module thermometer_to_binary (
    input [14:0] ith,
    output reg [3:0] binary
);

always @(*) begin
    case (ith)
        //16'b000000000000000: binary = 4'b0000; 	// ~0.0000
        16'b000000000000001: binary = 4'b0001; 	// ~0.1188
        16'b000000000000011: binary = 4'b0010; 	// ~0.2376
        16'b000000000000111: binary = 4'b0011; 	// ~0.3564
        16'b000000000001111: binary = 4'b0100; 	// ~0.4752
        16'b000000000011111: binary = 4'b0101; 	// ~0.5940
        16'b000000000111111: binary = 4'b0110; 	// ~0.7128
        16'b000000001111111: binary = 4'b0111; 	// ~0.8316
        16'b000000011111111: binary = 4'b1000; 	// ~0.9504
        16'b000000111111111: binary = 4'b1001; 	// ~1.0692
        16'b000001111111111: binary = 4'b1010; 	// ~1.1880
        16'b000011111111111: binary = 4'b1011; 	// ~1.3068
        16'b000111111111111: binary = 4'b1100; 	// ~1.4256
        16'b001111111111111: binary = 4'b1101; 	// ~1.5444
        16'b011111111111111: binary = 4'b1110; 	// ~1.6632
        16'b111111111111111: binary = 4'b1111;	// ~1.7820

        default: binary = 4'b0000; // Don't care
    endcase
end

endmodule
