magic
tech sky130A
magscale 1 2
timestamp 1706464016
<< viali >>
rect 901 82 935 116
rect 996 -737 1030 -703
rect 1682 -1125 1716 -1091
<< metal1 >>
rect 484 117 584 152
rect 892 117 946 122
rect 484 116 1052 117
rect 484 83 901 116
rect 484 52 584 83
rect 892 82 901 83
rect 935 83 1052 116
rect 935 82 946 83
rect 892 70 946 82
rect 499 -101 533 52
rect 608 -79 642 -78
rect 608 -101 666 -79
rect 499 -135 666 -101
rect 608 -156 666 -135
rect 632 -157 666 -156
rect 849 -111 883 -81
rect 849 -145 963 -111
rect 1018 -118 1052 83
rect 1780 -79 1814 -78
rect 1750 -97 1814 -79
rect 1750 -131 1893 -97
rect 1750 -138 1814 -131
rect 1750 -139 1784 -138
rect 849 -157 883 -145
rect 929 -197 963 -145
rect 929 -231 1543 -197
rect 747 -290 753 -238
rect 805 -290 811 -238
rect 1081 -311 1118 -231
rect 679 -443 815 -409
rect 597 -535 667 -501
rect 597 -878 631 -535
rect 633 -579 667 -535
rect 781 -639 815 -443
rect 1084 -632 1118 -311
rect 1859 -396 1893 -131
rect 1836 -402 1936 -396
rect 1596 -442 1936 -402
rect 1596 -544 1638 -442
rect 1836 -496 1936 -442
rect 1236 -584 1638 -544
rect 1598 -586 1638 -584
rect 1723 -596 1757 -593
rect 1710 -630 1757 -596
rect 687 -673 815 -639
rect 1346 -643 1380 -642
rect 687 -707 721 -673
rect 1225 -677 1551 -643
rect 983 -684 1047 -683
rect 982 -703 1047 -684
rect 982 -707 996 -703
rect 687 -737 996 -707
rect 1030 -712 1047 -703
rect 1318 -712 1381 -677
rect 1030 -737 1381 -712
rect 687 -741 1381 -737
rect 990 -743 1381 -741
rect 1001 -746 1381 -743
rect 1013 -749 1381 -746
rect 1723 -749 1757 -630
rect 1599 -783 1757 -749
rect 597 -912 1145 -878
rect 1599 -882 1633 -783
rect 1111 -943 1145 -912
rect 1568 -929 1633 -882
rect 1568 -942 1632 -929
rect 632 -1022 732 -966
rect 862 -1000 914 -994
rect 632 -1052 862 -1022
rect 1173 -1022 1533 -989
rect 914 -1023 1533 -1022
rect 914 -1052 1279 -1023
rect 632 -1056 1279 -1052
rect 632 -1066 732 -1056
rect 862 -1058 914 -1056
rect 1662 -1091 1762 -1056
rect 1662 -1125 1682 -1091
rect 1716 -1125 1762 -1091
rect 1662 -1156 1762 -1125
<< via1 >>
rect 753 -290 805 -238
rect 862 -1052 914 -1000
<< metal2 >>
rect 753 -238 805 -232
rect 753 -294 805 -290
rect 753 -296 904 -294
rect 762 -302 904 -296
rect 762 -336 905 -302
rect 871 -1000 905 -336
rect 856 -1052 862 -1000
rect 914 -1052 920 -1000
use sky130_fd_pr__pfet_01v8_LDQF7K  XM0
timestamp 1706462747
transform 1 0 707 0 1 -541
box -225 -269 225 269
use sky130_fd_pr__nfet_01v8_HZA4VB  XM1
timestamp 1706462747
transform 1 0 1356 0 1 -912
box -396 -252 396 252
use sky130_fd_pr__pfet_01v8_GEY2B5  XM2
timestamp 1706462747
transform 1 0 757 0 1 -118
box -275 -270 275 270
use sky130_fd_pr__pfet_01v8_KQKFM4  XM3
timestamp 1706462747
transform 1 0 1408 0 1 -109
box -526 -261 526 261
use sky130_fd_pr__nfet_01v8_5NW376  XM4
timestamp 1706462747
transform 0 -1 1421 1 0 -613
box -211 -461 211 461
<< labels >>
flabel metal1 1836 -496 1936 -396 0 FreeSans 256 0 0 0 V15
port 1 nsew
flabel metal1 484 52 584 152 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 1662 -1156 1762 -1056 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 632 -1066 732 -966 0 FreeSans 256 0 0 0 Vin
port 2 nsew
<< end >>
