magic
tech sky130A
magscale 1 2
timestamp 1704877912
<< error_p >>
rect -35 167 35 173
rect -35 133 -23 167
rect -35 127 35 133
rect -35 -133 35 -127
rect -35 -167 -23 -133
rect -35 -173 35 -167
<< pwell >>
rect -235 -305 235 305
<< nmos >>
rect -39 -95 39 95
<< ndiff >>
rect -97 83 -39 95
rect -97 -83 -85 83
rect -51 -83 -39 83
rect -97 -95 -39 -83
rect 39 83 97 95
rect 39 -83 51 83
rect 85 -83 97 83
rect 39 -95 97 -83
<< ndiffc >>
rect -85 -83 -51 83
rect 51 -83 85 83
<< psubdiff >>
rect -199 235 -103 269
rect 103 235 199 269
rect -199 173 -165 235
rect 165 173 199 235
rect -199 -235 -165 -173
rect 165 -235 199 -173
rect -199 -269 -103 -235
rect 103 -269 199 -235
<< psubdiffcont >>
rect -103 235 103 269
rect -199 -173 -165 173
rect 165 -173 199 173
rect -103 -269 103 -235
<< poly >>
rect -39 167 39 183
rect -39 133 -23 167
rect 23 133 39 167
rect -39 95 39 133
rect -39 -133 39 -95
rect -39 -167 -23 -133
rect 23 -167 39 -133
rect -39 -183 39 -167
<< polycont >>
rect -23 133 23 167
rect -23 -167 23 -133
<< locali >>
rect -199 235 -103 269
rect 103 235 199 269
rect -199 173 -165 235
rect 165 173 199 235
rect -39 133 -23 167
rect 23 133 39 167
rect -85 83 -51 99
rect -85 -99 -51 -83
rect 51 83 85 99
rect 51 -99 85 -83
rect -39 -167 -23 -133
rect 23 -167 39 -133
rect -199 -235 -165 -173
rect 165 -235 199 -173
rect -199 -269 -103 -235
rect 103 -269 199 -235
<< viali >>
rect -23 133 23 167
rect -85 -83 -51 83
rect 51 -83 85 83
rect -23 -167 23 -133
<< metal1 >>
rect -35 167 35 173
rect -35 133 -23 167
rect 23 133 35 167
rect -35 127 35 133
rect -91 83 -45 95
rect -91 -83 -85 83
rect -51 -83 -45 83
rect -91 -95 -45 -83
rect 45 83 91 95
rect 45 -83 51 83
rect 85 -83 91 83
rect 45 -95 91 -83
rect -35 -133 35 -127
rect -35 -167 -23 -133
rect 23 -167 35 -133
rect -35 -173 35 -167
<< properties >>
string FIXED_BBOX -182 -252 182 252
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.95 l 0.39 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
