magic
tech sky130A
magscale 1 2
timestamp 1705440136
<< checkpaint >>
rect -1260 -2460 1460 1460
<< locali >>
rect 834 500 976 554
rect 436 -20 582 44
<< metal1 >>
rect 1018 779 1218 780
rect 710 745 1218 779
rect 710 561 745 745
rect 774 600 834 658
rect 1018 580 1218 745
rect 710 497 777 561
rect 831 497 899 557
rect 710 496 744 497
rect 398 445 598 476
rect 398 411 829 445
rect 398 276 598 411
rect 865 404 899 497
rect 0 0 200 200
rect 0 -400 200 -200
rect 399 -221 433 276
rect 865 241 1068 404
rect 517 207 1068 241
rect 517 41 551 207
rect 868 204 1068 207
rect 517 7 583 41
rect 1270 40 1470 110
rect 518 -23 583 7
rect 1258 -18 1470 40
rect 660 -221 694 -78
rect 1270 -90 1470 -18
rect 399 -255 694 -221
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_FP437E  XM0
timestamp 1704962149
transform 1 0 921 0 1 11
box -521 -261 521 261
use sky130_fd_pr__nfet_01v8_L7T3GD  XM1
timestamp 1704336338
transform 1 0 805 0 1 528
box -211 -252 211 252
<< labels >>
flabel metal1 1270 -90 1470 110 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 1018 580 1218 780 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 398 276 598 476 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 868 204 1068 404 0 FreeSans 256 0 0 0 Vpamp
port 2 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vin
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vpamp
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
<< end >>
