magic
tech sky130A
magscale 1 2
timestamp 1696192038
<< pwell >>
rect -211 -310 211 310
<< nmos >>
rect -15 -100 15 100
<< ndiff >>
rect -73 88 -15 100
rect -73 -88 -61 88
rect -27 -88 -15 88
rect -73 -100 -15 -88
rect 15 88 73 100
rect 15 -88 27 88
rect 61 -88 73 88
rect 15 -100 73 -88
<< ndiffc >>
rect -61 -88 -27 88
rect 27 -88 61 88
<< psubdiff >>
rect -175 240 -79 274
rect 79 240 175 274
rect -175 178 -141 240
rect 141 178 175 240
rect -175 -240 -141 -178
rect 141 -240 175 -178
rect -175 -274 -79 -240
rect 79 -274 175 -240
<< psubdiffcont >>
rect -79 240 79 274
rect -175 -178 -141 178
rect 141 -178 175 178
rect -79 -274 79 -240
<< poly >>
rect -34 178 34 188
rect -34 144 -18 178
rect 16 144 34 178
rect -34 122 34 144
rect -15 100 15 122
rect -15 -122 15 -100
rect -34 -144 34 -122
rect -34 -178 -18 -144
rect 16 -178 34 -144
rect -34 -188 34 -178
<< polycont >>
rect -18 144 16 178
rect -18 -178 16 -144
<< locali >>
rect -175 240 -79 274
rect 79 240 175 274
rect -175 178 -141 240
rect -34 178 34 188
rect -34 144 -18 178
rect 16 144 34 178
rect -34 138 34 144
rect 141 178 175 240
rect -61 88 -27 104
rect -61 -104 -27 -88
rect 27 88 61 104
rect 27 -104 61 -88
rect -175 -240 -141 -178
rect -34 -144 34 -138
rect -34 -178 -18 -144
rect 16 -178 34 -144
rect -34 -188 34 -178
rect 141 -240 175 -178
rect -175 -274 -79 -240
rect 79 -274 175 -240
<< viali >>
rect -18 144 16 178
rect -61 -88 -27 88
rect 27 -88 61 88
rect -18 -178 16 -144
<< metal1 >>
rect -34 178 34 188
rect -34 144 -18 178
rect 16 144 34 178
rect -34 138 34 144
rect -67 88 -21 100
rect -67 -88 -61 88
rect -27 -88 -21 88
rect -67 -100 -21 -88
rect 21 88 67 100
rect 21 -88 27 88
rect 61 -88 67 88
rect 21 -100 67 -88
rect -34 -144 34 -138
rect -34 -178 -18 -144
rect 16 -178 34 -144
rect -34 -188 34 -178
<< properties >>
string FIXED_BBOX -158 -257 158 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
