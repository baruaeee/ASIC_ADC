magic
tech sky130A
magscale 1 2
timestamp 1706229878
<< nwell >>
rect -245 -261 245 261
<< pmos >>
rect -49 -42 49 42
<< pdiff >>
rect -107 30 -49 42
rect -107 -30 -95 30
rect -61 -30 -49 30
rect -107 -42 -49 -30
rect 49 30 107 42
rect 49 -30 61 30
rect 95 -30 107 30
rect 49 -42 107 -30
<< pdiffc >>
rect -95 -30 -61 30
rect 61 -30 95 30
<< nsubdiff >>
rect -175 191 -113 225
rect 113 191 175 225
<< nsubdiffcont >>
rect -113 191 113 225
<< poly >>
rect -49 123 49 139
rect -49 89 -33 123
rect 33 89 49 123
rect -49 42 49 89
rect -49 -89 49 -42
rect -49 -123 -33 -89
rect 33 -123 49 -89
rect -49 -139 49 -123
<< polycont >>
rect -33 89 33 123
rect -33 -123 33 -89
<< locali >>
rect -175 191 -113 225
rect 113 191 175 225
rect -49 89 -33 123
rect 33 89 49 123
rect -95 30 -61 46
rect -95 -46 -61 -30
rect 61 30 95 46
rect 61 -46 95 -30
rect -49 -123 -33 -89
rect 33 -123 49 -89
<< viali >>
rect -33 89 33 123
rect -95 -30 -61 30
rect 61 -30 95 30
rect -33 -123 33 -89
<< metal1 >>
rect -45 123 45 129
rect -45 89 -33 123
rect 33 89 45 123
rect -45 83 45 89
rect -101 30 -55 42
rect -101 -30 -95 30
rect -61 -30 -55 30
rect -101 -42 -55 -30
rect 55 30 101 42
rect 55 -30 61 30
rect 95 -30 101 30
rect 55 -42 101 -30
rect -45 -89 45 -83
rect -45 -123 -33 -89
rect 33 -123 45 -89
rect -45 -129 45 -123
<< properties >>
string FIXED_BBOX -192 -208 192 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.494 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
