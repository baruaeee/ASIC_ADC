magic
tech sky130A
magscale 1 2
timestamp 1706197322
<< error_p >>
rect -29 272 29 278
rect -29 238 -17 272
rect -29 232 29 238
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect -29 -278 29 -272
<< pwell >>
rect -211 -410 211 410
<< nmos >>
rect -15 -200 15 200
<< ndiff >>
rect -73 188 -15 200
rect -73 -188 -61 188
rect -27 -188 -15 188
rect -73 -200 -15 -188
rect 15 188 73 200
rect 15 -188 27 188
rect 61 -188 73 188
rect 15 -200 73 -188
<< ndiffc >>
rect -61 -188 -27 188
rect 27 -188 61 188
<< psubdiff >>
rect -141 340 -79 374
rect 79 340 175 374
rect 141 278 175 340
rect 141 -340 175 -278
rect -141 -374 -79 -340
rect 79 -374 175 -340
<< psubdiffcont >>
rect -79 340 79 374
rect 141 -278 175 278
rect -79 -374 79 -340
<< poly >>
rect -33 272 33 288
rect -33 238 -17 272
rect 17 238 33 272
rect -33 222 33 238
rect -15 200 15 222
rect -15 -222 15 -200
rect -33 -238 33 -222
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
<< polycont >>
rect -17 238 17 272
rect -17 -272 17 -238
<< locali >>
rect -141 340 -79 374
rect 79 340 175 374
rect 141 278 175 340
rect -33 238 -17 272
rect 17 238 33 272
rect -61 188 -27 204
rect -61 -204 -27 -188
rect 27 188 61 204
rect 27 -204 61 -188
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect 141 -340 175 -278
rect -141 -374 -79 -340
rect 79 -374 175 -340
<< viali >>
rect -17 238 17 272
rect -61 -188 -27 188
rect 27 -188 61 188
rect -17 -272 17 -238
<< metal1 >>
rect -29 272 29 278
rect -29 238 -17 272
rect 17 238 29 272
rect -29 232 29 238
rect -67 188 -21 200
rect -67 -188 -61 188
rect -27 -188 -21 188
rect -67 -200 -21 -188
rect 21 188 67 200
rect 21 -188 27 188
rect 61 -188 67 188
rect 21 -200 67 -188
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
<< properties >>
string FIXED_BBOX -158 -357 158 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
