magic
tech sky130A
magscale 1 2
timestamp 1706462747
<< nwell >>
rect -275 -270 275 270
<< pmos >>
rect -79 -51 79 51
<< pdiff >>
rect -137 39 -79 51
rect -137 -39 -125 39
rect -91 -39 -79 39
rect -137 -51 -79 -39
rect 79 39 137 51
rect 79 -39 91 39
rect 125 -39 137 39
rect 79 -51 137 -39
<< pdiffc >>
rect -125 -39 -91 39
rect 91 -39 125 39
<< nsubdiff >>
rect -205 200 -143 234
rect 143 200 205 234
<< nsubdiffcont >>
rect -143 200 143 234
<< poly >>
rect -79 132 79 148
rect -79 98 -63 132
rect 63 98 79 132
rect -79 51 79 98
rect -79 -98 79 -51
rect -79 -132 -63 -98
rect 63 -132 79 -98
rect -79 -148 79 -132
<< polycont >>
rect -63 98 63 132
rect -63 -132 63 -98
<< locali >>
rect -205 200 -143 234
rect 143 200 205 234
rect -79 98 -63 132
rect 63 98 79 132
rect -125 39 -91 55
rect -125 -55 -91 -39
rect 91 39 125 55
rect 91 -55 125 -39
rect -79 -132 -63 -98
rect 63 -132 79 -98
<< viali >>
rect -63 98 63 132
rect -125 -39 -91 39
rect 91 -39 125 39
rect -63 -132 63 -98
<< metal1 >>
rect -75 132 75 138
rect -75 98 -63 132
rect 63 98 75 132
rect -75 92 75 98
rect -131 39 -85 51
rect -131 -39 -125 39
rect -91 -39 -85 39
rect -131 -51 -85 -39
rect 85 39 131 51
rect 85 -39 91 39
rect 125 -39 131 39
rect 85 -51 131 -39
rect -75 -98 75 -92
rect -75 -132 -63 -98
rect 63 -132 75 -98
rect -75 -138 75 -132
<< properties >>
string FIXED_BBOX -222 -217 222 217
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.51 l 0.79 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
