magic
tech sky130A
magscale 1 2
timestamp 1706236419
<< error_p >>
rect -29 229 29 235
rect -29 195 -17 229
rect -29 189 29 195
rect -29 -195 29 -189
rect -29 -229 -17 -195
rect -29 -235 29 -229
<< pwell >>
rect -211 -367 211 367
<< nmos >>
rect -15 -157 15 157
<< ndiff >>
rect -73 145 -15 157
rect -73 -145 -61 145
rect -27 -145 -15 145
rect -73 -157 -15 -145
rect 15 145 73 157
rect 15 -145 27 145
rect 61 -145 73 145
rect 15 -157 73 -145
<< ndiffc >>
rect -61 -145 -27 145
rect 27 -145 61 145
<< psubdiff >>
rect -175 235 -141 297
rect -175 -297 -141 -235
<< psubdiffcont >>
rect -175 -235 -141 235
<< poly >>
rect -33 229 33 245
rect -33 195 -17 229
rect 17 195 33 229
rect -33 179 33 195
rect -15 157 15 179
rect -15 -179 15 -157
rect -33 -195 33 -179
rect -33 -229 -17 -195
rect 17 -229 33 -195
rect -33 -245 33 -229
<< polycont >>
rect -17 195 17 229
rect -17 -229 17 -195
<< locali >>
rect -175 235 -141 297
rect -33 195 -17 229
rect 17 195 33 229
rect -61 145 -27 161
rect -61 -161 -27 -145
rect 27 145 61 161
rect 27 -161 61 -145
rect -33 -229 -17 -195
rect 17 -229 33 -195
rect -175 -297 -141 -235
<< viali >>
rect -17 195 17 229
rect -61 -145 -27 145
rect 27 -145 61 145
rect -17 -229 17 -195
<< metal1 >>
rect -29 229 29 235
rect -29 195 -17 229
rect 17 195 29 229
rect -29 189 29 195
rect -67 145 -21 157
rect -67 -145 -61 145
rect -27 -145 -21 145
rect -67 -157 -21 -145
rect 21 145 67 157
rect 21 -145 27 145
rect 61 -145 67 145
rect 21 -157 67 -145
rect -29 -195 29 -189
rect -29 -229 -17 -195
rect 17 -229 29 -195
rect -29 -235 29 -229
<< properties >>
string FIXED_BBOX -158 -314 158 314
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.57 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
