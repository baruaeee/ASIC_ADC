magic
tech sky130A
magscale 1 2
timestamp 1702941823
<< checkpaint >>
rect -575 2329 2367 2339
rect -1313 2170 2367 2329
rect -1313 2117 2736 2170
rect -1313 2046 3105 2117
rect -1313 -713 3474 2046
rect -944 -766 3474 -713
rect -575 -819 3474 -766
rect -206 -872 3474 -819
rect 163 -925 3474 -872
rect 532 -978 3474 -925
<< error_s >>
rect 129 931 187 937
rect 129 897 141 931
rect 129 891 187 897
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_M479BZ  XM1
timestamp 0
transform 1 0 158 0 1 808
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 0
transform 1 0 896 0 1 760
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_L7T3GD  XM3
timestamp 0
transform 1 0 527 0 1 746
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_M479BZ  XM7
timestamp 0
transform 1 0 1265 0 1 649
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_M479BZ  XM9
timestamp 0
transform 1 0 1634 0 1 596
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_L7T3GD  XM10
timestamp 0
transform 1 0 2003 0 1 534
box -211 -252 211 252
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
