magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 1452 29 1458
rect -29 1418 -17 1452
rect -29 1412 29 1418
rect -29 -1418 29 -1412
rect -29 -1452 -17 -1418
rect -29 -1458 29 -1452
<< pwell >>
rect -211 -1590 211 1590
<< nmos >>
rect -15 -1380 15 1380
<< ndiff >>
rect -73 1368 -15 1380
rect -73 -1368 -61 1368
rect -27 -1368 -15 1368
rect -73 -1380 -15 -1368
rect 15 1368 73 1380
rect 15 -1368 27 1368
rect 61 -1368 73 1368
rect 15 -1380 73 -1368
<< ndiffc >>
rect -61 -1368 -27 1368
rect 27 -1368 61 1368
<< psubdiff >>
rect -175 1520 -79 1554
rect 79 1520 175 1554
rect -175 1458 -141 1520
rect 141 1458 175 1520
rect -175 -1520 -141 -1458
rect 141 -1520 175 -1458
rect -175 -1554 -79 -1520
rect 79 -1554 175 -1520
<< psubdiffcont >>
rect -79 1520 79 1554
rect -175 -1458 -141 1458
rect 141 -1458 175 1458
rect -79 -1554 79 -1520
<< poly >>
rect -33 1452 33 1468
rect -33 1418 -17 1452
rect 17 1418 33 1452
rect -33 1402 33 1418
rect -15 1380 15 1402
rect -15 -1402 15 -1380
rect -33 -1418 33 -1402
rect -33 -1452 -17 -1418
rect 17 -1452 33 -1418
rect -33 -1468 33 -1452
<< polycont >>
rect -17 1418 17 1452
rect -17 -1452 17 -1418
<< locali >>
rect -175 1520 -79 1554
rect 79 1520 175 1554
rect -175 1458 -141 1520
rect 141 1458 175 1520
rect -33 1418 -17 1452
rect 17 1418 33 1452
rect -61 1368 -27 1384
rect -61 -1384 -27 -1368
rect 27 1368 61 1384
rect 27 -1384 61 -1368
rect -33 -1452 -17 -1418
rect 17 -1452 33 -1418
rect -175 -1520 -141 -1458
rect 141 -1520 175 -1458
rect -175 -1554 -79 -1520
rect 79 -1554 175 -1520
<< viali >>
rect -17 1418 17 1452
rect -61 -1368 -27 1368
rect 27 -1368 61 1368
rect -17 -1452 17 -1418
<< metal1 >>
rect -29 1452 29 1458
rect -29 1418 -17 1452
rect 17 1418 29 1452
rect -29 1412 29 1418
rect -67 1368 -21 1380
rect -67 -1368 -61 1368
rect -27 -1368 -21 1368
rect -67 -1380 -21 -1368
rect 21 1368 67 1380
rect 21 -1368 27 1368
rect 61 -1368 67 1368
rect 21 -1380 67 -1368
rect -29 -1418 29 -1412
rect -29 -1452 -17 -1418
rect 17 -1452 29 -1418
rect -29 -1458 29 -1452
<< properties >>
string FIXED_BBOX -158 -1537 158 1537
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 13.8 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
