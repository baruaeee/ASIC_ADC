magic
tech sky130A
magscale 1 2
timestamp 1706400305
<< pwell >>
rect -351 210 351 252
rect -351 148 267 210
rect 333 148 351 210
rect -351 -252 351 148
<< nmos >>
rect -155 -42 155 42
<< ndiff >>
rect -213 30 -155 42
rect -213 -30 -201 30
rect -167 -30 -155 30
rect -213 -42 -155 -30
rect 155 30 213 42
rect 155 -30 167 30
rect 201 -30 213 30
rect 155 -42 213 -30
<< ndiffc >>
rect -201 -30 -167 30
rect 167 -30 201 30
<< psubdiff >>
rect 281 64 315 92
rect 281 -238 315 -176
<< psubdiffcont >>
rect 281 -176 315 64
<< poly >>
rect -155 114 155 130
rect -155 80 -139 114
rect 139 80 155 114
rect -155 42 155 80
rect -155 -80 155 -42
rect -155 -114 -139 -80
rect 139 -114 155 -80
rect -155 -130 155 -114
<< polycont >>
rect -139 80 139 114
rect -139 -114 139 -80
<< locali >>
rect -155 80 -139 114
rect 139 80 155 114
rect 281 64 315 92
rect -201 30 -167 46
rect -201 -46 -167 -30
rect 167 30 201 46
rect 167 -46 201 -30
rect -155 -114 -139 -80
rect 139 -114 155 -80
rect 281 -238 315 -176
<< viali >>
rect -139 80 139 114
rect -201 -30 -167 30
rect 167 -30 201 30
rect -139 -114 139 -80
<< metal1 >>
rect -151 114 151 120
rect -151 80 -139 114
rect 139 80 151 114
rect -151 74 151 80
rect -207 30 -161 42
rect -207 -30 -201 30
rect -167 -30 -161 30
rect -207 -42 -161 -30
rect 161 30 207 42
rect 161 -30 167 30
rect 201 -30 207 30
rect 161 -42 207 -30
rect -151 -80 151 -74
rect -151 -114 -139 -80
rect 139 -114 151 -80
rect -151 -120 151 -114
<< properties >>
string FIXED_BBOX -298 -199 298 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 1.55 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
