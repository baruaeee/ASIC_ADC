magic
tech sky130A
timestamp 1703732895
<< pwell >>
rect -208 -126 208 126
<< nmos >>
rect -110 -21 110 21
<< ndiff >>
rect -139 15 -110 21
rect -139 -15 -133 15
rect -116 -15 -110 15
rect -139 -21 -110 -15
rect 110 15 139 21
rect 110 -15 116 15
rect 133 -15 139 15
rect 110 -21 139 -15
<< ndiffc >>
rect -133 -15 -116 15
rect 116 -15 133 15
<< psubdiff >>
rect -190 91 -142 108
rect 142 91 190 108
rect -190 60 -173 91
rect 173 60 190 91
rect -190 -91 -173 -60
rect 173 -91 190 -60
rect -190 -108 -142 -91
rect 142 -108 190 -91
<< psubdiffcont >>
rect -142 91 142 108
rect -190 -60 -173 60
rect 173 -60 190 60
rect -142 -108 142 -91
<< poly >>
rect -110 57 110 65
rect -110 40 -102 57
rect 102 40 110 57
rect -110 21 110 40
rect -110 -40 110 -21
rect -110 -57 -102 -40
rect 102 -57 110 -40
rect -110 -65 110 -57
<< polycont >>
rect -102 40 102 57
rect -102 -57 102 -40
<< locali >>
rect -190 91 -142 108
rect 142 91 190 108
rect -190 60 -173 91
rect 173 60 190 91
rect -110 40 -102 57
rect 102 40 110 57
rect -133 15 -116 23
rect -133 -23 -116 -15
rect 116 15 133 23
rect 116 -23 133 -15
rect -110 -57 -102 -40
rect 102 -57 110 -40
rect -190 -91 -173 -60
rect 173 -91 190 -60
rect -190 -108 -142 -91
rect 142 -108 190 -91
<< viali >>
rect -102 40 102 57
rect -133 -15 -116 15
rect 116 -15 133 15
rect -102 -57 102 -40
<< metal1 >>
rect -108 57 108 60
rect -108 40 -102 57
rect 102 40 108 57
rect -108 37 108 40
rect -136 15 -113 21
rect -136 -15 -133 15
rect -116 -15 -113 15
rect -136 -21 -113 -15
rect 113 15 136 21
rect 113 -15 116 15
rect 133 -15 136 15
rect 113 -21 136 -15
rect -108 -40 108 -37
rect -108 -57 -102 -40
rect 102 -57 108 -40
rect -108 -60 108 -57
<< properties >>
string FIXED_BBOX -181 -99 181 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 2.2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
