magic
tech sky130A
magscale 1 2
timestamp 1702941819
<< checkpaint >>
rect 1426 -766 6738 2258
rect 10220 -1084 15532 1940
<< error_s >>
rect 2668 999 2703 1016
rect 2669 998 2703 999
rect 2669 962 2739 998
rect 5425 962 5478 963
rect 2686 928 2757 962
rect 5407 928 5478 962
rect 2686 583 2756 928
rect 5408 927 5478 928
rect 5425 893 5496 927
rect 5776 893 5811 910
rect 2686 547 2739 583
rect 5425 530 5495 893
rect 5777 892 5811 893
rect 5777 856 5847 892
rect 7033 856 7086 857
rect 5607 825 5665 831
rect 5607 791 5619 825
rect 5794 822 5865 856
rect 7015 822 7086 856
rect 5607 785 5665 791
rect 5607 613 5665 619
rect 5607 579 5619 613
rect 5607 573 5665 579
rect 5425 494 5478 530
rect 5794 477 5864 822
rect 7016 821 7086 822
rect 7033 787 7104 821
rect 8354 787 8389 804
rect 5794 441 5847 477
rect 7033 424 7103 787
rect 8355 786 8389 787
rect 8355 750 8425 786
rect 8741 750 8794 751
rect 8372 716 8443 750
rect 8723 716 8794 750
rect 7033 388 7086 424
rect 8372 371 8442 716
rect 8724 715 8794 716
rect 8741 681 8812 715
rect 8554 648 8612 654
rect 8554 614 8566 648
rect 8554 608 8612 614
rect 8554 454 8612 460
rect 8554 420 8566 454
rect 8554 414 8612 420
rect 8372 335 8425 371
rect 8741 318 8811 681
rect 8741 282 8794 318
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_MQKFYN  XM1
timestamp 0
transform 1 0 1343 0 1 808
box -1396 -261 1396 261
use sky130_fd_pr__nfet_01v8_RYBV7U  XM2
timestamp 0
transform 1 0 4082 0 1 746
box -1396 -252 1396 252
use sky130_fd_pr__pfet_01v8_VZ9GCW  XM3
timestamp 0
transform 1 0 7729 0 1 596
box -696 -261 696 261
use sky130_fd_pr__nfet_01v8_L7T3GD  XM4
timestamp 0
transform 1 0 8583 0 1 534
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_MQKFYN  XM5
timestamp 0
transform 1 0 10137 0 1 490
box -1396 -261 1396 261
use sky130_fd_pr__nfet_01v8_RYBV7U  XM6
timestamp 0
transform 1 0 12876 0 1 428
box -1396 -252 1396 252
use sky130_fd_pr__pfet_01v8_M479BZ  XM7
timestamp 0
transform 1 0 5636 0 1 702
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_LHZPBA  XM10
timestamp 0
transform 1 0 6440 0 1 640
box -646 -252 646 252
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
