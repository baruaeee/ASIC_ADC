magic
tech sky130A
magscale 1 2
timestamp 1704387395
<< nwell >>
rect -243 -261 243 261
<< pmos >>
rect -47 -42 47 42
<< pdiff >>
rect -105 30 -47 42
rect -105 -30 -93 30
rect -59 -30 -47 30
rect -105 -42 -47 -30
rect 47 30 105 42
rect 47 -30 59 30
rect 93 -30 105 30
rect 47 -42 105 -30
<< pdiffc >>
rect -93 -30 -59 30
rect 59 -30 93 30
<< nsubdiff >>
rect -207 191 -111 225
rect 111 191 207 225
rect -207 129 -173 191
rect 173 129 207 191
rect -207 -191 -173 -129
rect 173 -191 207 -129
rect -207 -225 -111 -191
rect 111 -225 207 -191
<< nsubdiffcont >>
rect -111 191 111 225
rect -207 -129 -173 129
rect 173 -129 207 129
rect -111 -225 111 -191
<< poly >>
rect -47 123 47 139
rect -47 89 -31 123
rect 31 89 47 123
rect -47 42 47 89
rect -47 -89 47 -42
rect -47 -123 -31 -89
rect 31 -123 47 -89
rect -47 -139 47 -123
<< polycont >>
rect -31 89 31 123
rect -31 -123 31 -89
<< locali >>
rect -207 191 -111 225
rect 111 191 207 225
rect -207 129 -173 191
rect 173 129 207 191
rect -47 89 -31 123
rect 31 89 47 123
rect -93 30 -59 46
rect -93 -46 -59 -30
rect 59 30 93 46
rect 59 -46 93 -30
rect -47 -123 -31 -89
rect 31 -123 47 -89
rect -207 -191 -173 -129
rect 173 -191 207 -129
rect -207 -225 -111 -191
rect 111 -225 207 -191
<< viali >>
rect -31 89 31 123
rect -93 -30 -59 30
rect 59 -30 93 30
rect -31 -123 31 -89
<< metal1 >>
rect -43 123 43 129
rect -43 89 -31 123
rect 31 89 43 123
rect -43 83 43 89
rect -99 30 -53 42
rect -99 -30 -93 30
rect -59 -30 -53 30
rect -99 -42 -53 -30
rect 53 30 99 42
rect 53 -30 59 30
rect 93 -30 99 30
rect 53 -42 99 -30
rect -43 -89 43 -83
rect -43 -123 -31 -89
rect 31 -123 43 -89
rect -43 -129 43 -123
<< properties >>
string FIXED_BBOX -190 -208 190 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.47 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
