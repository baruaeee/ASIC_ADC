* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : pre_therm                                    *
* Netlisted  : Wed Dec 11 23:34:13 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_C_CDNS_733956442880                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_C_CDNS_733956442880 1
** N=1 EP=1 FDC=0
.ends M1M2_C_CDNS_733956442880

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: PYL1CON_C_CDNS_733956442881                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt PYL1CON_C_CDNS_733956442881 1 2
** N=2 EP=2 FDC=0
.ends PYL1CON_C_CDNS_733956442881

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_733956442882                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_733956442882 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_733956442882

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_733956442884                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_733956442884 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_733956442884

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733956442880                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733956442880 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6.5e-07 W=4.45e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733956442880

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733956442881                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733956442881 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=6.3e-07 W=7.9e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733956442881

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv01f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv01f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733956442881 $T=575 1630 0 0 $X=390 $Y=1445
X1 3 L1M1_C_CDNS_733956442882 $T=575 1630 0 0 $X=410 $Y=1485
X2 4 L1M1_C_CDNS_733956442884 $T=1085 695 0 0 $X=970 $Y=530
X3 2 4 3 nfet_01v8_CDNS_733956442880 $T=295 475 0 0 $X=-110 $Y=325
X4 1 4 3 pfet_01v8_CDNS_733956442881 $T=295 2820 0 0 $X=-150 $Y=2640
.ends inv01f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_733956442885                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_733956442885 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_733956442885

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733956442882                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733956442882 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 pfet_01v8 L=1.05e-06 W=5.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733956442882

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733956442883                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733956442883 1 2 3 4
** N=10 EP=4 FDC=1
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=1.02e-06 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733956442883

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: preampF                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt preampF 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733956442881 $T=415 2135 0 0 $X=230 $Y=1950
X1 3 L1M1_C_CDNS_733956442882 $T=415 2135 0 0 $X=250 $Y=1990
X2 4 L1M1_C_CDNS_733956442884 $T=1100 3570 0 90 $X=935 $Y=3455
X3 1 L1M1_C_CDNS_733956442885 $T=130 995 0 0 $X=15 $Y=470
X4 4 L1M1_C_CDNS_733956442885 $T=570 995 0 0 $X=455 $Y=470
X5 4 2 3 1 pfet_01v8_CDNS_733956442882 $T=825 3430 0 270 $X=645 $Y=1935
X6 4 1 3 2 nfet_01v8_CDNS_733956442883 $T=430 485 1 180 $X=-125 $Y=335
.ends preampF

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pre_therm                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pre_therm
** N=5 EP=0 FDC=4
X0 1 M1M2_C_CDNS_733956442880 $T=390 2575 0 90 $X=230 $Y=2445
X1 2 M1M2_C_CDNS_733956442880 $T=2730 685 0 0 $X=2600 $Y=525
X2 3 4 5 2 inv01f $T=1630 0 0 0 $X=1450 $Y=-265
X3 3 4 1 5 preampF $T=0 0 0 0 $X=-180 $Y=-265
.ends pre_therm
