* NGSPICE file created from th01.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_9DPZTU w_n291_n261# a_n153_n42# a_n95_n139# a_95_n42#
+ VSUBS
X0 a_95_n42# a_n95_n139# a_n153_n42# w_n291_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.95
C0 w_n291_n261# a_n153_n42# 0.0499f
C1 a_n95_n139# a_n153_n42# 0.014f
C2 a_n95_n139# w_n291_n261# 0.419f
C3 a_n153_n42# a_95_n42# 0.0249f
C4 w_n291_n261# a_95_n42# 0.0499f
C5 a_n95_n139# a_95_n42# 0.014f
C6 a_95_n42# VSUBS 0.0313f
C7 a_n153_n42# VSUBS 0.0313f
C8 a_n95_n139# VSUBS 0.289f
C9 w_n291_n261# VSUBS 1.36f
.ends

.subckt sky130_fd_pr__nfet_01v8_586EUA a_n97_n95# a_n199_n269# a_n39_n183# a_39_n95#
X0 a_39_n95# a_n39_n183# a_n97_n95# a_n199_n269# sky130_fd_pr__nfet_01v8 ad=0.275 pd=2.48 as=0.275 ps=2.48 w=0.95 l=0.39
C0 a_n39_n183# a_39_n95# 0.0127f
C1 a_n97_n95# a_39_n95# 0.1f
C2 a_n97_n95# a_n39_n183# 0.0127f
C3 a_39_n95# a_n199_n269# 0.135f
C4 a_n97_n95# a_n199_n269# 0.135f
C5 a_n39_n183# a_n199_n269# 0.381f
.ends

.subckt sky130_fd_pr__nfet_01v8_PJBF84 a_n248_n222# a_n146_n48# a_88_n48# a_n88_n136#
X0 a_88_n48# a_n88_n136# a_n146_n48# a_n248_n222# sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.54 as=0.139 ps=1.54 w=0.48 l=0.88
C0 a_n88_n136# a_88_n48# 0.0146f
C1 a_n146_n48# a_88_n48# 0.03f
C2 a_n146_n48# a_n88_n136# 0.0146f
C3 a_88_n48# a_n248_n222# 0.088f
C4 a_n146_n48# a_n248_n222# 0.088f
C5 a_n88_n136# a_n248_n222# 0.649f
.ends

.subckt sky130_fd_pr__pfet_01v8_RVEGTV a_n69_n175# a_n127_n78# w_n265_n297# a_69_n78#
+ VSUBS
X0 a_69_n78# a_n69_n175# a_n127_n78# w_n265_n297# sky130_fd_pr__pfet_01v8 ad=0.226 pd=2.14 as=0.226 ps=2.14 w=0.78 l=0.69
C0 w_n265_n297# a_n127_n78# 0.0718f
C1 a_n69_n175# a_n127_n78# 0.0173f
C2 a_n69_n175# w_n265_n297# 0.338f
C3 a_n127_n78# a_69_n78# 0.0574f
C4 w_n265_n297# a_69_n78# 0.0718f
C5 a_n69_n175# a_69_n78# 0.0173f
C6 a_69_n78# VSUBS 0.0474f
C7 a_n127_n78# VSUBS 0.0474f
C8 a_n69_n175# VSUBS 0.227f
C9 w_n265_n297# VSUBS 1.41f
.ends

.subckt th01 Vp Vin Vout Vn
XXM2 Vp Vp Vin m1_732_n84# Vn sky130_fd_pr__pfet_01v8_9DPZTU
XXM3 Vn Vn Vin m1_732_n84# sky130_fd_pr__nfet_01v8_586EUA
XXM4 Vn Vn Vout m1_732_n84# sky130_fd_pr__nfet_01v8_PJBF84
XXM5 m1_732_n84# Vp Vp Vout Vn sky130_fd_pr__pfet_01v8_RVEGTV
C0 Vn Vp 0.167f
C1 Vn Vin 0.0827f
C2 Vn m1_732_n84# 0.18f
C3 Vout Vp 0.0895f
C4 Vout Vin 1.54e-19
C5 Vout m1_732_n84# 0.174f
C6 Vin Vp 0.228f
C7 Vn Vout 0.0643f
C8 m1_732_n84# Vp 0.305f
C9 m1_732_n84# Vin 0.174f
C10 Vin 0 0.683f
C11 Vp 0 2.57f
C12 Vout 0 0.247f
C13 m1_732_n84# 0 0.96f
C14 Vn 0 0.0948f
.ends

