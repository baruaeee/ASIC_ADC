magic
tech sky130A
magscale 1 2
timestamp 1706323418
<< pwell >>
rect 21812 -6304 21857 -6259
rect 26818 -6386 26842 -6384
rect 26818 -6456 26844 -6386
rect 26820 -6458 26844 -6456
<< psubdiff >>
rect 21642 -275 21676 -214
rect 21642 -309 21717 -275
rect 21645 -310 21717 -309
rect 21281 -4702 21349 -4668
<< nsubdiff >>
rect 20956 -4273 20990 -4211
<< locali >>
rect 27163 194 27211 228
rect 21642 -251 21676 -214
rect 21509 -2633 21543 -1601
rect 20956 -4249 20990 -4211
rect 21315 -4702 21335 -4668
<< viali >>
rect 27211 194 27245 228
rect 21642 -285 21676 -251
rect 20956 -4283 20990 -4249
rect 21281 -4702 21315 -4668
<< metal1 >>
rect 21123 1137 26569 1171
rect 21123 1119 23763 1137
rect 23533 1105 23763 1119
rect 23533 1097 23703 1105
rect 23669 1075 23703 1097
rect 22896 828 22948 834
rect 22896 770 22948 776
rect 23836 726 23842 778
rect 23894 726 23900 778
rect 25680 614 25732 620
rect 27037 619 27345 653
rect 25680 552 25732 558
rect 27311 473 27345 619
rect 27311 439 27503 473
rect 22806 89 22843 409
rect 27205 228 27251 240
rect 27205 194 27211 228
rect 27245 194 27251 228
rect 27205 182 27251 194
rect 22506 52 22843 89
rect 22806 -33 22843 52
rect 22806 -43 23096 -33
rect 25737 -43 25771 159
rect 22806 -70 24587 -43
rect 23059 -77 24587 -70
rect 24683 -77 25771 -43
rect 27211 98 27245 182
rect 27469 163 27503 439
rect 27469 129 28903 163
rect 21630 -246 21688 -245
rect 21630 -251 21694 -246
rect 23059 -250 23096 -77
rect 24446 -235 24480 -77
rect 27211 -89 27428 98
rect 27211 -123 27429 -89
rect 21630 -291 21642 -251
rect 21676 -252 21694 -251
rect 21642 -310 21694 -304
rect 21111 -484 21363 -457
rect 21111 -491 21374 -484
rect 21111 -1985 21145 -491
rect 21340 -492 21374 -491
rect 21199 -624 21205 -572
rect 21257 -624 21263 -572
rect 21912 -595 22173 -561
rect 21213 -1613 21247 -624
rect 21912 -645 21946 -595
rect 22139 -805 22173 -595
rect 27395 -768 27429 -123
rect 22139 -839 22499 -805
rect 27177 -815 27429 -768
rect 27177 -849 27515 -815
rect 27177 -864 27429 -849
rect 27395 -865 27429 -864
rect 27481 -1523 27515 -849
rect 27481 -1557 28807 -1523
rect 21213 -1647 21935 -1613
rect 22203 -1915 22503 -1881
rect 27481 -1887 27515 -1557
rect 22203 -1985 22237 -1915
rect 27253 -1921 27515 -1887
rect 20865 -2019 21369 -1985
rect 21483 -2019 22237 -1985
rect 20556 -2608 20756 -2574
rect 20556 -2660 20618 -2608
rect 20670 -2660 20756 -2608
rect 20556 -2774 20756 -2660
rect 20865 -3287 20899 -2019
rect 27562 -2054 27614 -2048
rect 27562 -2112 27614 -2106
rect 28636 -2182 28688 -2176
rect 28636 -2240 28688 -2234
rect 27215 -2467 27481 -2433
rect 27447 -2678 27481 -2467
rect 28243 -2678 28373 -2673
rect 27447 -2712 27733 -2678
rect 28179 -2696 28373 -2678
rect 28416 -2687 28468 -2681
rect 28179 -2712 28416 -2696
rect 28339 -2730 28416 -2712
rect 28416 -2745 28468 -2739
rect 28773 -2801 28807 -1557
rect 28869 -2756 28903 129
rect 28003 -2807 28807 -2801
rect 27475 -2835 28807 -2807
rect 28842 -2808 28848 -2756
rect 28900 -2808 28906 -2756
rect 27475 -2841 28013 -2835
rect 27475 -2979 27509 -2841
rect 27979 -2957 28013 -2841
rect 27253 -3013 27509 -2979
rect 27560 -3262 27612 -3256
rect 27560 -3320 27612 -3314
rect 28418 -3266 28470 -3260
rect 28418 -3324 28470 -3318
rect 27237 -3551 27455 -3517
rect 20790 -3654 20842 -3648
rect 20790 -3712 20842 -3706
rect 27421 -3751 27455 -3551
rect 28618 -3722 28670 -3716
rect 27421 -3785 27881 -3751
rect 28159 -3769 28618 -3726
rect 28618 -3780 28670 -3774
rect 27541 -3919 28245 -3885
rect 28773 -3893 28807 -2835
rect 28869 -3716 28903 -2808
rect 28856 -3722 28908 -3716
rect 28856 -3780 28908 -3774
rect 27541 -4075 27575 -3919
rect 28367 -3927 28807 -3893
rect 27251 -4109 27575 -4075
rect 20944 -4249 21002 -4243
rect 20944 -4283 20956 -4249
rect 20990 -4283 21002 -4249
rect 20944 -4289 21002 -4283
rect 20956 -4362 20990 -4289
rect 28344 -4320 28396 -4314
rect 20941 -4414 20947 -4362
rect 20999 -4414 21005 -4362
rect 27564 -4388 27570 -4336
rect 27622 -4388 27628 -4336
rect 28344 -4378 28396 -4372
rect 21457 -4588 21739 -4569
rect 21457 -4622 22034 -4588
rect 21127 -4704 21133 -4652
rect 21185 -4668 21191 -4652
rect 21275 -4668 21321 -4656
rect 21185 -4702 21281 -4668
rect 21315 -4702 21321 -4668
rect 21185 -4704 21191 -4702
rect 21275 -4714 21321 -4702
rect 20572 -5008 20578 -4956
rect 20630 -5008 20636 -4956
rect 20941 -4966 20947 -4962
rect 20587 -5339 20621 -5008
rect 20940 -5014 20947 -4966
rect 20999 -5014 21005 -4962
rect 20940 -5050 21002 -5014
rect 21088 -5050 21911 -5030
rect 21088 -5056 21932 -5050
rect 21088 -5064 21880 -5056
rect 21877 -5093 21880 -5064
rect 21880 -5114 21932 -5108
rect 20587 -5373 20669 -5339
rect 22000 -6082 22034 -4622
rect 27257 -4651 27367 -4617
rect 27333 -4895 27367 -4651
rect 28037 -4829 28071 -4777
rect 28001 -4853 28035 -4841
rect 28037 -4853 28079 -4829
rect 28001 -4861 28127 -4853
rect 28001 -4867 28134 -4861
rect 28001 -4895 28082 -4867
rect 27333 -4919 28082 -4895
rect 27333 -4925 28134 -4919
rect 27333 -4929 28105 -4925
rect 22496 -5021 22548 -5015
rect 22548 -5064 22669 -5030
rect 22496 -5079 22548 -5073
rect 22635 -5073 22669 -5064
rect 23853 -5073 25199 -5039
rect 22635 -5107 23887 -5073
rect 23853 -5181 23887 -5107
rect 25165 -5227 25199 -5073
rect 28771 -5123 28805 -3927
rect 28869 -4818 28903 -3780
rect 28838 -4870 28844 -4818
rect 28896 -4870 28903 -4818
rect 27567 -5181 27965 -5147
rect 28167 -5157 28805 -5123
rect 27567 -5205 27601 -5181
rect 25825 -5239 27601 -5205
rect 28869 -5221 28903 -4870
rect 25825 -5276 25872 -5239
rect 28725 -5255 28903 -5221
rect 24862 -5363 24914 -5357
rect 23512 -5429 23518 -5377
rect 23570 -5429 23576 -5377
rect 25825 -5369 25859 -5276
rect 28498 -5392 28504 -5340
rect 28556 -5392 28562 -5340
rect 24862 -5421 24914 -5415
rect 27648 -5598 27700 -5592
rect 27326 -5706 27332 -5654
rect 27384 -5706 27390 -5654
rect 27648 -5656 27700 -5650
rect 26124 -5832 26176 -5826
rect 26124 -5890 26176 -5884
rect 22000 -6134 22060 -6082
rect 22000 -6195 22034 -6134
rect 23814 -6160 23866 -6154
rect 20634 -6254 20640 -6202
rect 20692 -6254 20698 -6202
rect 21812 -6218 21866 -6211
rect 23814 -6218 23866 -6212
rect 21811 -6268 21817 -6218
rect 21770 -6270 21817 -6268
rect 21869 -6268 21875 -6218
rect 25096 -6256 25148 -6250
rect 21869 -6270 21970 -6268
rect 21770 -6295 21970 -6270
rect 21480 -6340 21970 -6295
rect 23057 -6316 23063 -6264
rect 23115 -6316 23121 -6264
rect 21770 -6420 21970 -6340
rect 21770 -6455 22981 -6420
rect 24313 -6447 24347 -6309
rect 25096 -6314 25148 -6308
rect 26394 -6280 26446 -6274
rect 26394 -6338 26446 -6332
rect 26818 -6386 26842 -6384
rect 26818 -6447 26844 -6386
rect 28215 -6447 28249 -6131
rect 28725 -6447 28759 -5255
rect 21770 -6468 21970 -6455
rect 23587 -6481 28759 -6447
<< via1 >>
rect 22896 776 22948 828
rect 23842 726 23894 778
rect 25680 558 25732 614
rect 21642 -285 21676 -252
rect 21676 -285 21694 -252
rect 21642 -304 21694 -285
rect 21205 -624 21257 -572
rect 20618 -2660 20670 -2608
rect 27562 -2106 27614 -2054
rect 28636 -2234 28688 -2182
rect 28416 -2739 28468 -2687
rect 28848 -2808 28900 -2756
rect 27560 -3314 27612 -3262
rect 28418 -3318 28470 -3266
rect 20790 -3706 20842 -3654
rect 28618 -3774 28670 -3722
rect 28856 -3774 28908 -3722
rect 20947 -4414 20999 -4362
rect 27570 -4388 27622 -4336
rect 28344 -4372 28396 -4320
rect 21133 -4704 21185 -4652
rect 20578 -5008 20630 -4956
rect 20947 -5014 20999 -4962
rect 21880 -5108 21932 -5056
rect 28082 -4919 28134 -4867
rect 22496 -5073 22548 -5021
rect 28844 -4870 28896 -4818
rect 23518 -5429 23570 -5377
rect 24862 -5415 24914 -5363
rect 28504 -5392 28556 -5340
rect 27648 -5650 27700 -5598
rect 27332 -5706 27384 -5654
rect 26124 -5884 26176 -5832
rect 20640 -6254 20692 -6202
rect 23814 -6212 23866 -6160
rect 21817 -6270 21869 -6218
rect 23063 -6316 23115 -6264
rect 25096 -6308 25148 -6256
rect 26394 -6332 26446 -6280
<< metal2 >>
rect 20991 1251 27157 1285
rect 20991 -783 21025 1251
rect 22792 820 22848 827
rect 22890 820 22896 828
rect 22792 818 22896 820
rect 22848 783 22896 818
rect 22890 776 22896 783
rect 22948 776 22954 828
rect 23851 784 23885 1251
rect 23842 778 23894 784
rect 22792 753 22848 762
rect 23842 720 23894 726
rect 25447 513 25481 1251
rect 27123 763 27157 1251
rect 25576 558 25680 614
rect 25732 558 25738 614
rect 25343 479 25481 513
rect 21464 16 21504 42
rect 21371 -40 21380 16
rect 21436 -32 21504 16
rect 21436 -40 21445 -32
rect 21636 -261 21642 -252
rect 21214 -295 21642 -261
rect 21214 -566 21248 -295
rect 21636 -304 21642 -295
rect 21694 -304 21700 -252
rect 21205 -572 21257 -566
rect 21205 -630 21257 -624
rect 20991 -817 21335 -783
rect 20991 -1691 21025 -817
rect 20627 -1725 21025 -1691
rect 20627 -2602 20661 -1725
rect 20991 -2090 21025 -1725
rect 27556 -2062 27562 -2054
rect 20991 -2108 21054 -2090
rect 27364 -2098 27562 -2062
rect 20991 -2133 21025 -2108
rect 20618 -2608 20670 -2602
rect 20618 -2666 20670 -2660
rect 20627 -2836 20661 -2666
rect 20610 -2892 20619 -2836
rect 20675 -2892 20684 -2836
rect 20769 -3004 20778 -2948
rect 20834 -3004 20843 -2948
rect 20588 -3175 20621 -3174
rect 20789 -3175 20823 -3004
rect 20588 -3209 20823 -3175
rect 20588 -3230 20621 -3209
rect 20587 -3663 20621 -3230
rect 20784 -3663 20790 -3654
rect 20587 -3697 20790 -3663
rect 20784 -3706 20790 -3697
rect 20842 -3706 20848 -3654
rect 20947 -4362 20999 -4356
rect 20947 -4420 20999 -4414
rect 20567 -4874 20576 -4818
rect 20632 -4874 20641 -4818
rect 20587 -4950 20621 -4874
rect 20578 -4956 20630 -4950
rect 20956 -4956 20990 -4420
rect 27364 -4474 27400 -2098
rect 27556 -2106 27562 -2098
rect 27614 -2106 27620 -2054
rect 28630 -2234 28636 -2182
rect 28688 -2184 28694 -2182
rect 28688 -2234 28758 -2184
rect 28676 -2260 28758 -2234
rect 28532 -2685 28588 -2676
rect 28410 -2739 28416 -2687
rect 28468 -2689 28474 -2687
rect 28468 -2737 28532 -2689
rect 28468 -2739 28474 -2737
rect 28532 -2750 28588 -2741
rect 28710 -2810 28758 -2260
rect 28846 -2685 28902 -2676
rect 28846 -2750 28902 -2741
rect 28498 -2858 28758 -2810
rect 28848 -2756 28900 -2750
rect 28848 -2814 28900 -2808
rect 28498 -3234 28546 -2858
rect 27554 -3268 27560 -3262
rect 27463 -3309 27560 -3268
rect 21133 -4652 21185 -4646
rect 21133 -4710 21185 -4704
rect 21142 -4794 21176 -4710
rect 27463 -4723 27504 -3309
rect 27554 -3314 27560 -3309
rect 27612 -3314 27618 -3262
rect 28458 -3266 28546 -3234
rect 28412 -3318 28418 -3266
rect 28470 -3318 28546 -3266
rect 28460 -3342 28546 -3318
rect 27570 -4336 27622 -4330
rect 28338 -4372 28344 -4320
rect 28396 -4322 28402 -4320
rect 28498 -4322 28546 -3342
rect 28612 -3774 28618 -3722
rect 28670 -3724 28676 -3722
rect 28850 -3724 28856 -3722
rect 28670 -3772 28856 -3724
rect 28670 -3774 28676 -3772
rect 28850 -3774 28856 -3772
rect 28908 -3774 28914 -3722
rect 28396 -4370 28676 -4322
rect 28396 -4372 28402 -4370
rect 27570 -4394 27622 -4388
rect 21122 -4850 21131 -4794
rect 21187 -4850 21196 -4794
rect 23848 -4919 23889 -4771
rect 24481 -4821 24667 -4781
rect 24964 -4784 25468 -4744
rect 26700 -4764 27504 -4723
rect 24481 -4831 24872 -4821
rect 24617 -4834 24872 -4831
rect 25056 -4834 25323 -4821
rect 24617 -4871 25323 -4834
rect 24836 -4880 25072 -4871
rect 20578 -5014 20630 -5008
rect 20947 -4962 20999 -4956
rect 22794 -4979 23561 -4944
rect 23848 -4960 24908 -4919
rect 20947 -5020 20999 -5014
rect 22490 -5030 22496 -5021
rect 21879 -5056 22496 -5030
rect 21874 -5108 21880 -5056
rect 21932 -5064 22496 -5056
rect 21932 -5108 21938 -5064
rect 22490 -5073 22496 -5064
rect 22548 -5073 22554 -5021
rect 23526 -5371 23561 -4979
rect 24867 -5363 24908 -4960
rect 25273 -4977 25323 -4871
rect 25428 -4874 25468 -4784
rect 25757 -4823 25951 -4781
rect 26179 -4815 26489 -4777
rect 25909 -4863 25951 -4823
rect 26451 -4829 26489 -4815
rect 27577 -4829 27615 -4394
rect 25428 -4914 25812 -4874
rect 25909 -4905 26353 -4863
rect 26451 -4867 27615 -4829
rect 28408 -4865 28464 -4856
rect 25772 -4958 25812 -4914
rect 26311 -4915 26353 -4905
rect 26311 -4957 27559 -4915
rect 28076 -4919 28082 -4867
rect 28134 -4869 28140 -4867
rect 28134 -4917 28408 -4869
rect 28134 -4919 28140 -4917
rect 28408 -4930 28464 -4921
rect 25273 -5027 25701 -4977
rect 25772 -4998 26206 -4958
rect 25651 -5033 25701 -5027
rect 26166 -5014 26206 -4998
rect 27517 -4999 27559 -4957
rect 25651 -5083 26083 -5033
rect 26166 -5054 27378 -5014
rect 27517 -5041 28551 -4999
rect 26033 -5109 26083 -5083
rect 26033 -5159 26175 -5109
rect 23518 -5377 23570 -5371
rect 24856 -5415 24862 -5363
rect 24914 -5415 24920 -5363
rect 23518 -5435 23570 -5429
rect 26125 -5832 26175 -5159
rect 27338 -5648 27378 -5054
rect 28509 -5334 28551 -5041
rect 28504 -5340 28556 -5334
rect 28504 -5398 28556 -5392
rect 27642 -5600 27648 -5598
rect 27534 -5648 27648 -5600
rect 27332 -5654 27384 -5648
rect 27332 -5712 27384 -5706
rect 23072 -5872 23689 -5838
rect 21805 -6182 21814 -6126
rect 21870 -6182 21879 -6126
rect 20640 -6202 20692 -6196
rect 21818 -6212 21868 -6182
rect 20640 -6260 20692 -6254
rect 21817 -6218 21869 -6212
rect 20642 -6510 20690 -6260
rect 23072 -6258 23106 -5872
rect 23655 -6169 23689 -5872
rect 26118 -5884 26124 -5832
rect 26176 -5884 26182 -5832
rect 23808 -6169 23814 -6160
rect 23655 -6203 23814 -6169
rect 23808 -6212 23814 -6203
rect 23866 -6212 23872 -6160
rect 27534 -6240 27582 -5648
rect 27642 -5650 27648 -5648
rect 27700 -5650 27706 -5598
rect 28628 -6240 28676 -4370
rect 28844 -4818 28896 -4812
rect 28842 -4865 28844 -4856
rect 28896 -4865 28898 -4856
rect 28842 -4930 28898 -4921
rect 25090 -6258 25096 -6256
rect 21817 -6276 21869 -6270
rect 23063 -6264 23115 -6258
rect 23063 -6322 23115 -6316
rect 24976 -6306 25096 -6258
rect 24976 -6510 25024 -6306
rect 25090 -6308 25096 -6306
rect 25148 -6308 25154 -6256
rect 26388 -6282 26394 -6280
rect 26354 -6332 26394 -6282
rect 26446 -6332 26452 -6280
rect 27534 -6288 28676 -6240
rect 26354 -6510 26402 -6332
rect 27534 -6510 27582 -6288
rect 20642 -6558 27582 -6510
<< via2 >>
rect 22792 762 22848 818
rect 21380 -40 21436 16
rect 20619 -2892 20675 -2836
rect 20778 -3004 20834 -2948
rect 20576 -4874 20632 -4818
rect 28532 -2741 28588 -2685
rect 28846 -2741 28902 -2685
rect 21131 -4850 21187 -4794
rect 28408 -4921 28464 -4865
rect 21814 -6182 21870 -6126
rect 28842 -4870 28844 -4865
rect 28844 -4870 28896 -4865
rect 28896 -4870 28898 -4865
rect 28842 -4921 28898 -4870
<< metal3 >>
rect 22787 821 22853 823
rect 22732 818 22853 821
rect 22732 762 22792 818
rect 22848 762 22853 818
rect 22732 757 22853 762
rect 21375 16 21441 21
rect 21375 -40 21380 16
rect 21436 -40 21441 16
rect 21375 -45 21441 -40
rect 21377 -183 21439 -45
rect 22732 -51 22794 757
rect 22403 -113 22794 -51
rect 20863 -245 21567 -183
rect 20863 -1795 20925 -245
rect 21505 -331 21567 -245
rect 22403 -331 22465 -113
rect 21505 -393 22465 -331
rect 20775 -1857 20925 -1795
rect 20614 -2836 20680 -2831
rect 20614 -2892 20619 -2836
rect 20675 -2892 20680 -2836
rect 20614 -2897 20680 -2892
rect 20616 -3103 20678 -2897
rect 20775 -2943 20837 -1857
rect 28527 -2682 28593 -2680
rect 28841 -2682 28907 -2680
rect 28527 -2685 28907 -2682
rect 28527 -2741 28532 -2685
rect 28588 -2741 28846 -2685
rect 28902 -2741 28907 -2685
rect 28527 -2744 28907 -2741
rect 28527 -2746 28593 -2744
rect 28841 -2746 28907 -2744
rect 20773 -2948 20839 -2943
rect 20773 -3004 20778 -2948
rect 20834 -3004 20839 -2948
rect 20773 -3009 20839 -3004
rect 20573 -3165 20678 -3103
rect 20573 -4813 20635 -3165
rect 21128 -4789 21190 -4729
rect 21126 -4794 21192 -4789
rect 20571 -4818 20637 -4813
rect 20571 -4874 20576 -4818
rect 20632 -4874 20637 -4818
rect 21126 -4828 21131 -4794
rect 21187 -4828 21192 -4794
rect 20571 -4879 20637 -4874
rect 21121 -4892 21127 -4828
rect 21191 -4892 21197 -4828
rect 28403 -4862 28469 -4860
rect 28837 -4862 28903 -4860
rect 28403 -4865 28903 -4862
rect 28403 -4921 28408 -4865
rect 28464 -4921 28842 -4865
rect 28898 -4921 28903 -4865
rect 28403 -4924 28903 -4921
rect 28403 -4926 28469 -4924
rect 28837 -4926 28903 -4924
rect 21810 -6114 21874 -6108
rect 21809 -6178 21810 -6121
rect 21874 -6178 21875 -6121
rect 21809 -6182 21814 -6178
rect 21870 -6182 21875 -6178
rect 21809 -6187 21875 -6182
rect 21811 -6289 21873 -6187
<< via3 >>
rect 21127 -4850 21131 -4828
rect 21131 -4850 21187 -4828
rect 21187 -4850 21191 -4828
rect 21127 -4892 21191 -4850
rect 21810 -6126 21874 -6114
rect 21810 -6178 21814 -6126
rect 21814 -6178 21870 -6126
rect 21870 -6178 21874 -6126
<< metal4 >>
rect 21126 -4828 21192 -4827
rect 21126 -4892 21127 -4828
rect 21191 -4853 21192 -4828
rect 21283 -4833 21811 -4771
rect 21283 -4853 21345 -4833
rect 21191 -4892 21345 -4853
rect 21126 -4893 21345 -4892
rect 21128 -4959 21345 -4893
rect 21749 -5653 21811 -4833
rect 21749 -5715 21873 -5653
rect 21811 -6113 21873 -5715
rect 21809 -6114 21875 -6113
rect 21809 -6178 21810 -6114
rect 21874 -6178 21875 -6114
rect 21809 -6179 21875 -6178
use th12  th12_0
timestamp 1706270854
transform 1 0 20666 0 1 -2146
box 278 -1078 1572 236
use preamp  x0
timestamp 1706271137
transform -1 0 24300 0 1 -210
box 394 136 1494 1340
use th01  x1
timestamp 1706270854
transform 1 0 21652 0 1 -5044
box 316 -1456 1968 6
use th02  x2
timestamp 1706270854
transform 1 0 23352 0 1 -5442
box 378 -1044 1518 426
use th03  x3
timestamp 1706270854
transform 1 0 24566 0 1 -5385
box 516 -1083 1680 238
use th04  x4
timestamp 1706270854
transform 1 0 26058 0 1 -5340
box 374 -1126 1336 148
use th05  x5
timestamp 1706270876
transform -1 0 29178 0 1 -1669
box 474 -1043 1620 148
use th06  x6
timestamp 1706231216
transform -1 0 28658 0 1 -2810
box 200 -976 1084 2
use th07  x7
timestamp 1706236611
transform -1 0 28708 0 1 -3916
box 314 -1014 1088 32
use th08  x8
timestamp 1706233216
transform 1 0 27292 0 1 -5110
box 356 -1052 1272 -2
use th09  x9
timestamp 1706236419
transform -1 0 25784 0 1 676
box 368 -754 1692 526
use th10  x10
timestamp 1706270854
transform 1 0 21036 0 1 -876
box 270 -794 1168 452
use th11  x11
timestamp 1706241174
transform 1 0 20160 0 1 -5462
box 466 -880 1630 468
use th13  x13
timestamp 1706270854
transform -1 0 27716 0 1 562
box 438 -680 2042 646
use th14  x14
timestamp 1706271011
transform 1 0 20086 0 1 -3934
box 502 -804 2110 674
use th15  x15
timestamp 1706283436
transform 1 0 20536 0 1 462
box 470 -808 2076 675
<< labels >>
flabel metal1 21770 -6468 21970 -6268 0 FreeSans 256 0 0 0 Vn
port 17 nsew
flabel metal1 27228 -102 27428 98 0 FreeSans 256 0 0 0 Vp
port 1 nsew
flabel metal1 20556 -2774 20756 -2574 0 FreeSans 256 0 0 0 Vin
port 0 nsew
<< end >>
