* NGSPICE file created from adc1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X a_208_47# a_75_199#
+ a_544_297# a_315_47# a_201_297#
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPWR VGND 0.0735f
C1 a_75_199# a_544_297# 0.0176f
C2 a_201_297# B1 0.00594f
C3 C1 VPB 0.0394f
C4 a_315_47# VGND 0.00427f
C5 a_75_199# VPB 0.0486f
C6 VGND A3 0.0161f
C7 VGND a_208_47# 0.00302f
C8 X B1 7.79e-20
C9 VGND A2 0.0119f
C10 VPWR A1 0.0151f
C11 VGND a_201_297# 0.00403f
C12 a_315_47# A1 0.00313f
C13 B1 a_544_297# 1.13e-19
C14 VPB B1 0.0292f
C15 a_75_199# C1 0.0628f
C16 A2 A1 0.0689f
C17 X VGND 0.0609f
C18 a_201_297# A1 0.011f
C19 a_315_47# VPWR 0.00154f
C20 VGND a_544_297# 0.00256f
C21 VPWR A3 0.0181f
C22 VGND VPB 0.00772f
C23 VPWR a_208_47# 8.35e-19
C24 VPWR A2 0.0174f
C25 X A1 1.2e-19
C26 C1 B1 0.066f
C27 a_75_199# B1 0.102f
C28 VPWR a_201_297# 0.211f
C29 a_315_47# A2 0.00335f
C30 A3 a_208_47# 3.65e-19
C31 VPB A1 0.0306f
C32 A3 A2 0.0747f
C33 A3 a_201_297# 0.00642f
C34 A2 a_208_47# 0.00102f
C35 X VPWR 0.0676f
C36 C1 VGND 0.0181f
C37 a_75_199# VGND 0.362f
C38 a_201_297# A2 0.0112f
C39 VPWR a_544_297# 0.0105f
C40 X A3 0.00317f
C41 VPWR VPB 0.0749f
C42 X a_208_47# 1.91e-19
C43 X A2 3.01e-19
C44 C1 A1 3.21e-19
C45 VPB A3 0.0268f
C46 a_75_199# A1 0.0696f
C47 X a_201_297# 0.0131f
C48 VGND B1 0.0171f
C49 a_201_297# a_544_297# 0.00702f
C50 VPB A2 0.0376f
C51 VPB a_201_297# 0.00186f
C52 C1 VPWR 0.0146f
C53 a_75_199# VPWR 0.109f
C54 X a_544_297# 2.35e-19
C55 A1 B1 0.0716f
C56 a_315_47# a_75_199# 0.0202f
C57 X VPB 0.0107f
C58 a_75_199# A3 0.163f
C59 a_75_199# a_208_47# 0.0159f
C60 a_75_199# A2 0.0621f
C61 C1 a_201_297# 0.00243f
C62 a_75_199# a_201_297# 0.16f
C63 VPWR B1 0.0125f
C64 VGND A1 0.0113f
C65 C1 X 5.14e-20
C66 a_75_199# X 0.0959f
C67 VGND VNB 0.437f
C68 VPWR VNB 0.365f
C69 X VNB 0.0906f
C70 C1 VNB 0.148f
C71 B1 VNB 0.0947f
C72 A1 VNB 0.101f
C73 A2 VNB 0.11f
C74 A3 VNB 0.0908f
C75 VPB VNB 0.782f
C76 a_201_297# VNB 0.00345f
C77 a_75_199# VNB 0.205f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_181_47# a_109_47# a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_181_47# VGND 0.00261f
C1 a_27_47# a_181_47# 0.00401f
C2 B VPWR 0.128f
C3 C X 0.0149f
C4 A VPWR 0.0185f
C5 VPWR VGND 0.0475f
C6 VPWR a_27_47# 0.145f
C7 A a_109_47# 6.45e-19
C8 a_109_47# VGND 0.00123f
C9 a_27_47# a_109_47# 0.00517f
C10 VPB VPWR 0.0795f
C11 A B 0.0869f
C12 VPWR X 0.0766f
C13 B VGND 0.00714f
C14 B a_27_47# 0.0625f
C15 A VGND 0.0154f
C16 A a_27_47# 0.157f
C17 a_181_47# C 0.00151f
C18 a_27_47# VGND 0.134f
C19 VPB B 0.0836f
C20 A VPB 0.0426f
C21 B X 0.00111f
C22 VPWR C 0.00464f
C23 VPB VGND 0.00604f
C24 VPB a_27_47# 0.0501f
C25 X VGND 0.0708f
C26 a_27_47# X 0.087f
C27 VPWR a_181_47# 3.97e-19
C28 B C 0.0746f
C29 VPB X 0.0121f
C30 C VGND 0.0703f
C31 a_27_47# C 0.186f
C32 VPWR a_109_47# 3.29e-19
C33 VPB C 0.0347f
C34 VGND VNB 0.3f
C35 X VNB 0.0923f
C36 C VNB 0.12f
C37 A VNB 0.174f
C38 VPWR VNB 0.274f
C39 B VNB 0.102f
C40 VPB VNB 0.516f
C41 a_27_47# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
C0 VGND VPWR 0.353f
C1 VPB VPWR 0.0625f
C2 VPB VGND 0.0797f
C3 VPWR VNB 0.47f
C4 VGND VNB 0.427f
C5 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VGND VPWR 0.546f
C1 VPB VPWR 0.0787f
C2 VPB VGND 0.116f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_384_47# a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
C0 B1 A1 0.0817f
C1 VPB A2 0.0373f
C2 a_81_21# B1 0.148f
C3 A2 VPWR 0.0201f
C4 VGND A2 0.0495f
C5 a_384_47# VPWR 4.08e-19
C6 a_299_297# A2 0.0468f
C7 VPB VPWR 0.068f
C8 VPB X 0.0108f
C9 A2 A1 0.0921f
C10 a_384_47# VGND 0.00366f
C11 VPB VGND 0.00713f
C12 X VPWR 0.0847f
C13 a_299_297# a_384_47# 1.48e-19
C14 VPB a_299_297# 0.0111f
C15 a_384_47# A1 0.00884f
C16 VGND VPWR 0.0579f
C17 VGND X 0.0512f
C18 VPB A1 0.0264f
C19 a_299_297# VPWR 0.202f
C20 a_81_21# A2 7.47e-19
C21 A1 VPWR 0.0209f
C22 a_299_297# VGND 0.00772f
C23 VGND A1 0.0786f
C24 a_81_21# a_384_47# 0.00138f
C25 VPB a_81_21# 0.0593f
C26 a_299_297# A1 0.0585f
C27 VPB B1 0.0387f
C28 a_81_21# VPWR 0.146f
C29 a_81_21# X 0.112f
C30 B1 VPWR 0.0196f
C31 X B1 3.04e-20
C32 a_81_21# VGND 0.173f
C33 VGND B1 0.0181f
C34 a_81_21# a_299_297# 0.0821f
C35 a_81_21# A1 0.0568f
C36 a_299_297# B1 0.00863f
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_pr__nfet_01v8_D7Y3TR a_n63_n101# a_n33_n75# a_n249_n145# a_63_n75#
+ a_n125_n75#
X0 a_63_n75# a_n63_n101# a_n33_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.233 pd=2.12 as=0.124 ps=1.08 w=0.75 l=0.15
X1 a_n33_n75# a_n63_n101# a_n125_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.08 as=0.233 ps=2.12 w=0.75 l=0.15
C0 a_n125_n75# a_n33_n75# 0.113f
C1 a_n63_n101# a_63_n75# 0.0104f
C2 a_63_n75# a_n33_n75# 0.113f
C3 a_n63_n101# a_n33_n75# 0.0186f
C4 a_n63_n101# a_n125_n75# 0.00451f
C5 a_63_n75# a_n249_n145# 0.0963f
C6 a_n33_n75# a_n249_n145# 0.0361f
C7 a_n125_n75# a_n249_n145# 0.105f
C8 a_n63_n101# a_n249_n145# 0.294f
.ends

.subckt sky130_fd_pr__pfet_01v8_2ZD99F w_n349_n261# a_n153_n139# a_n211_n42# a_153_n42#
+ VSUBS
X0 a_153_n42# a_n153_n139# a_n211_n42# w_n349_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.53
C0 a_n153_n139# a_n211_n42# 0.0177f
C1 w_n349_n261# a_153_n42# 0.0179f
C2 a_153_n42# a_n211_n42# 0.0169f
C3 w_n349_n261# a_n211_n42# 0.034f
C4 a_153_n42# a_n153_n139# 0.0177f
C5 w_n349_n261# a_n153_n139# 0.388f
C6 a_153_n42# VSUBS 0.0558f
C7 a_n211_n42# VSUBS 0.0456f
C8 a_n153_n139# VSUBS 0.556f
C9 w_n349_n261# VSUBS 1.16f
.ends

.subckt sky130_fd_pr__nfet_01v8_2BW22M a_154_n42# a_n154_n130# a_n314_n182# a_n212_n42#
X0 a_154_n42# a_n154_n130# a_n212_n42# a_n314_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.54
C0 a_n212_n42# a_154_n42# 0.0169f
C1 a_n154_n130# a_154_n42# 0.0178f
C2 a_n154_n130# a_n212_n42# 0.0178f
C3 a_154_n42# a_n314_n182# 0.0737f
C4 a_n212_n42# a_n314_n182# 0.0816f
C5 a_n154_n130# a_n314_n182# 0.924f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJP3BL a_15_n150# w_n211_n369# a_n73_n150# a_n33_n247#
+ VSUBS
X0 a_15_n150# a_n33_n247# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.15
C0 a_n33_n247# a_n73_n150# 0.0267f
C1 w_n211_n369# a_15_n150# 0.0292f
C2 a_15_n150# a_n73_n150# 0.242f
C3 w_n211_n369# a_n73_n150# 0.0292f
C4 a_15_n150# a_n33_n247# 0.0267f
C5 w_n211_n369# a_n33_n247# 0.19f
C6 a_15_n150# VSUBS 0.126f
C7 a_n73_n150# VSUBS 0.126f
C8 a_n33_n247# VSUBS 0.146f
C9 w_n211_n369# VSUBS 1.02f
.ends

.subckt sky130_fd_pr__nfet_01v8_LH5FDA a_n150_n130# a_276_n182# a_n208_n42# a_150_n42#
X0 a_150_n42# a_n150_n130# a_n208_n42# a_276_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.5
C0 a_n208_n42# a_150_n42# 0.0172f
C1 a_n150_n130# a_150_n42# 0.0176f
C2 a_n150_n130# a_n208_n42# 0.0176f
C3 a_150_n42# a_276_n182# 0.0815f
C4 a_n208_n42# a_276_n182# 0.0736f
C5 a_n150_n130# a_276_n182# 0.904f
.ends

.subckt th02 Vin V02 m1_983_133# Vp m1_571_144# Vn
XXM0 Vin Vn Vn m1_983_133# m1_983_133# sky130_fd_pr__nfet_01v8_D7Y3TR
XXM1 Vp Vin m1_571_144# m1_983_133# Vn sky130_fd_pr__pfet_01v8_2ZD99F
XXM2 m1_571_144# Vp Vn Vp sky130_fd_pr__nfet_01v8_2BW22M
XXM3 V02 Vp Vp m1_983_133# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_983_133# Vn V02 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 m1_571_144# Vn 0.00115f
C1 Vp Vn 0.0235f
C2 m1_983_133# V02 0.155f
C3 Vp m1_571_144# 0.176f
C4 m1_983_133# Vn 0.216f
C5 m1_571_144# m1_983_133# 0.0183f
C6 Vp m1_983_133# 0.366f
C7 Vin V02 0.00845f
C8 Vin Vn 0.0263f
C9 m1_571_144# Vin 0.332f
C10 Vp Vin 0.25f
C11 V02 Vn 0.00239f
C12 Vin m1_983_133# 0.279f
C13 m1_571_144# V02 0.011f
C14 Vp V02 0.118f
C15 Vn 0 0.263f
C16 V02 0 0.334f
C17 m1_983_133# 0 1.44f
C18 Vp 0 3.16f
C19 m1_571_144# 0 0.252f
C20 Vin 0 0.949f
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 VPWR Y 0.209f
C1 VPWR VPB 0.0521f
C2 A VGND 0.0638f
C3 A Y 0.0894f
C4 VGND Y 0.155f
C5 A VPB 0.0742f
C6 VGND VPB 0.00649f
C7 A VPWR 0.0631f
C8 VGND VPWR 0.0423f
C9 Y VPB 0.0061f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X a_29_53# a_183_297# a_111_297#
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 a_29_53# VPB 0.0491f
C1 C A 0.0343f
C2 B C 0.0802f
C3 a_29_53# a_111_297# 0.005f
C4 VGND C 0.0161f
C5 VPB A 0.0377f
C6 X VPB 0.0109f
C7 B VPB 0.0962f
C8 VGND VPB 0.00724f
C9 a_111_297# A 0.00223f
C10 a_183_297# VPWR 8.13e-19
C11 a_29_53# A 0.242f
C12 a_29_53# X 0.0991f
C13 a_29_53# B 0.121f
C14 VGND a_111_297# 3.96e-19
C15 a_29_53# VGND 0.217f
C16 X A 0.00127f
C17 B A 0.0787f
C18 B X 6.52e-19
C19 VGND A 0.0187f
C20 VPWR C 0.00457f
C21 VGND X 0.036f
C22 B VGND 0.0152f
C23 VPWR VPB 0.0649f
C24 VPWR a_111_297# 5.94e-19
C25 a_29_53# a_183_297# 0.00868f
C26 a_29_53# VPWR 0.0833f
C27 VPB C 0.0396f
C28 a_183_297# A 0.00239f
C29 VPWR A 0.00936f
C30 VPWR X 0.0885f
C31 B VPWR 0.147f
C32 a_183_297# VGND 5.75e-19
C33 VPWR VGND 0.0459f
C34 a_29_53# C 0.0857f
C35 VGND VNB 0.306f
C36 X VNB 0.0882f
C37 A VNB 0.117f
C38 C VNB 0.16f
C39 B VNB 0.117f
C40 VPWR VNB 0.253f
C41 VPB VNB 0.516f
C42 a_29_53# VNB 0.18f
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
C0 VPB VPWR 0.0858f
C1 VGND VPWR 0.903f
C2 VGND VPB 0.161f
C3 VPWR VNB 0.867f
C4 VGND VNB 0.761f
C5 VPB VNB 0.605f
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPB VGND 0.00456f
C1 VPB B 0.0367f
C2 VGND A 0.0486f
C3 B A 0.0584f
C4 VGND VPWR 0.0314f
C5 B VPWR 0.0148f
C6 Y a_109_297# 0.0113f
C7 VPB Y 0.0139f
C8 A Y 0.0471f
C9 B VGND 0.0451f
C10 VPWR Y 0.0995f
C11 VPB A 0.0415f
C12 VPWR a_109_297# 0.00638f
C13 VPB VPWR 0.0449f
C14 VPWR A 0.0528f
C15 VGND Y 0.154f
C16 B Y 0.0877f
C17 VGND a_109_297# 0.00128f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X a_193_297# a_465_47#
+ a_205_47# a_109_297# a_27_47#
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
C0 a_205_47# a_27_47# 0.00762f
C1 C1 A1 1.77e-20
C2 B2 VPB 0.0256f
C3 B2 X 6.77e-20
C4 B2 B1 0.0784f
C5 VPB A1 0.0343f
C6 a_109_297# VPWR 0.15f
C7 X A1 2.77e-19
C8 a_465_47# X 1.56e-19
C9 B2 a_27_47# 0.0959f
C10 C1 VPWR 0.0139f
C11 B1 A1 0.0609f
C12 VGND a_193_297# 0.00438f
C13 VGND A2 0.0168f
C14 a_205_47# VGND 0.00156f
C15 a_193_297# A2 0.00683f
C16 a_27_47# A1 0.0984f
C17 VPB VPWR 0.0799f
C18 a_27_47# a_465_47# 0.013f
C19 X VPWR 0.0897f
C20 C1 a_109_297# 0.00739f
C21 B1 VPWR 0.00982f
C22 a_27_47# VPWR 0.099f
C23 a_109_297# VPB 0.00421f
C24 VGND B2 0.0174f
C25 a_109_297# X 3.99e-19
C26 B2 a_193_297# 0.00126f
C27 C1 VPB 0.0367f
C28 C1 X 5.03e-20
C29 a_109_297# B1 0.00736f
C30 C1 B1 6.46e-19
C31 VGND A1 0.0126f
C32 VGND a_465_47# 0.00257f
C33 a_193_297# A1 0.0109f
C34 a_27_47# a_109_297# 0.0961f
C35 X VPB 0.0113f
C36 A1 A2 0.0692f
C37 C1 a_27_47# 0.0792f
C38 B1 VPB 0.0321f
C39 B1 X 9.58e-20
C40 VGND VPWR 0.0722f
C41 a_193_297# VPWR 0.169f
C42 a_27_47# VPB 0.0512f
C43 a_27_47# X 0.0921f
C44 VPWR A2 0.0209f
C45 a_205_47# VPWR 1.62e-19
C46 a_27_47# B1 0.112f
C47 VGND a_109_297# 0.00284f
C48 a_193_297# a_109_297# 0.0927f
C49 VGND C1 0.0196f
C50 a_465_47# A1 7.06e-19
C51 B2 VPWR 0.00842f
C52 C1 A2 9.03e-21
C53 VGND VPB 0.00844f
C54 a_193_297# VPB 0.00774f
C55 VGND X 0.061f
C56 a_193_297# X 0.00367f
C57 VPWR A1 0.0161f
C58 VPB A2 0.027f
C59 VGND B1 0.0133f
C60 a_465_47# VPWR 5.05e-19
C61 X A2 0.00157f
C62 a_193_297# B1 0.00869f
C63 B2 a_109_297# 0.0133f
C64 C1 B2 0.0726f
C65 VGND a_27_47# 0.395f
C66 a_193_297# a_27_47# 0.144f
C67 a_109_297# A1 1.05e-19
C68 a_27_47# A2 0.153f
C69 VGND VNB 0.437f
C70 X VNB 0.0919f
C71 VPWR VNB 0.364f
C72 A2 VNB 0.0896f
C73 A1 VNB 0.106f
C74 B1 VNB 0.108f
C75 B2 VNB 0.0887f
C76 C1 VNB 0.139f
C77 VPB VNB 0.782f
C78 a_193_297# VNB 0.0011f
C79 a_109_297# VNB 7.11e-19
C80 a_27_47# VNB 0.216f
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X a_256_47# a_584_47#
+ a_93_21# a_250_297# a_346_47#
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
C0 B2 A2 1.46e-19
C1 A1 X 6.03e-20
C2 A3 a_256_47# 4.42e-19
C3 a_93_21# VGND 0.251f
C4 a_346_47# VPWR 0.00109f
C5 B2 VPWR 0.0108f
C6 A3 X 2.45e-19
C7 a_93_21# a_250_297# 0.188f
C8 VGND a_256_47# 0.00394f
C9 X VGND 0.06f
C10 a_93_21# A2 0.0747f
C11 a_93_21# VPWR 0.0907f
C12 VPB B1 0.0276f
C13 X a_250_297# 5.42e-19
C14 B2 VPB 0.0355f
C15 A2 a_256_47# 0.00256f
C16 B1 a_346_47# 5.39e-20
C17 B2 B1 0.0823f
C18 VGND a_584_47# 0.00683f
C19 A2 X 1.19e-19
C20 a_256_47# VPWR 9.47e-19
C21 X VPWR 0.0849f
C22 a_250_297# a_584_47# 2.43e-19
C23 A1 VGND 0.0133f
C24 VPB a_93_21# 0.0485f
C25 a_93_21# B1 0.0774f
C26 A3 VGND 0.00974f
C27 a_584_47# VPWR 9.47e-19
C28 a_93_21# a_346_47# 0.0119f
C29 A1 a_250_297# 0.0129f
C30 B2 a_93_21# 0.0147f
C31 A3 a_250_297# 0.00602f
C32 VPB X 0.0108f
C33 B1 a_256_47# 2.07e-20
C34 B1 X 3.83e-20
C35 A2 A1 0.0971f
C36 A3 A2 0.0788f
C37 A1 VPWR 0.016f
C38 a_250_297# VGND 0.0072f
C39 A3 VPWR 0.0158f
C40 A2 VGND 0.0114f
C41 B1 a_584_47# 0.00143f
C42 VGND VPWR 0.076f
C43 a_93_21# a_256_47# 0.0114f
C44 A2 a_250_297# 0.0129f
C45 a_93_21# X 0.0841f
C46 a_250_297# VPWR 0.313f
C47 VPB A1 0.0296f
C48 B1 A1 0.0965f
C49 VPB A3 0.0291f
C50 A3 B1 7.88e-22
C51 A1 a_346_47# 0.00465f
C52 A2 VPWR 0.0133f
C53 B2 A1 3.14e-19
C54 a_93_21# a_584_47# 0.00278f
C55 B2 A3 9.12e-20
C56 VPB VGND 0.00788f
C57 B1 VGND 0.0344f
C58 VGND a_346_47# 0.00514f
C59 B2 VGND 0.0469f
C60 VPB a_250_297# 0.00616f
C61 B1 a_250_297# 0.0125f
C62 a_93_21# A1 0.0641f
C63 A3 a_93_21# 0.124f
C64 B2 a_250_297# 0.0344f
C65 VPB A2 0.0287f
C66 B1 A2 1.44e-20
C67 VPB VPWR 0.0756f
C68 A2 a_346_47# 0.00252f
C69 B1 VPWR 0.01f
C70 VGND VNB 0.465f
C71 VPWR VNB 0.365f
C72 X VNB 0.0937f
C73 B2 VNB 0.14f
C74 B1 VNB 0.101f
C75 A1 VNB 0.0951f
C76 A2 VNB 0.0921f
C77 A3 VNB 0.0929f
C78 VPB VNB 0.782f
C79 a_250_297# VNB 0.0278f
C80 a_93_21# VNB 0.151f
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X a_277_297# a_205_297# a_27_297#
+ a_109_297#
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 a_277_297# a_27_297# 0.00876f
C1 D VPWR 0.00503f
C2 B A 0.0639f
C3 X VPB 0.0109f
C4 D C 0.0954f
C5 VPWR A 0.00769f
C6 a_109_297# VGND 7.58e-19
C7 D a_27_297# 0.054f
C8 B VGND 0.0159f
C9 C A 0.028f
C10 D VPB 0.0405f
C11 a_27_297# A 0.163f
C12 VPWR VGND 0.0546f
C13 A VPB 0.033f
C14 a_277_297# X 6.43e-20
C15 C VGND 0.0191f
C16 a_27_297# VGND 0.235f
C17 a_109_297# VPWR 9.23e-19
C18 B VPWR 0.193f
C19 VGND VPB 0.00796f
C20 a_109_297# C 0.00356f
C21 B C 0.0917f
C22 a_27_297# a_109_297# 0.00695f
C23 A X 0.00133f
C24 B a_27_297# 0.159f
C25 a_277_297# A 2.28e-19
C26 C VPWR 0.00723f
C27 B VPB 0.106f
C28 a_205_297# VGND 3.36e-19
C29 a_27_297# VPWR 0.084f
C30 VGND X 0.0354f
C31 VPWR VPB 0.075f
C32 a_277_297# VGND 4.65e-19
C33 D A 2.13e-19
C34 a_27_297# C 0.158f
C35 C VPB 0.0338f
C36 a_27_297# VPB 0.0517f
C37 D VGND 0.0517f
C38 B X 6.42e-19
C39 a_277_297# B 2.29e-19
C40 a_205_297# VPWR 5.16e-19
C41 VGND A 0.016f
C42 VPWR X 0.0878f
C43 a_277_297# VPWR 7.48e-19
C44 a_205_297# C 0.00261f
C45 B D 0.00287f
C46 a_277_297# C 5.54e-19
C47 a_205_297# a_27_297# 0.00412f
C48 a_27_297# X 0.0991f
C49 VGND VNB 0.367f
C50 X VNB 0.0883f
C51 A VNB 0.109f
C52 C VNB 0.105f
C53 D VNB 0.175f
C54 B VNB 0.115f
C55 VPWR VNB 0.29f
C56 VPB VNB 0.605f
C57 a_27_297# VNB 0.163f
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
C0 VPB VGND 0.35f
C1 VGND VPWR 1.57f
C2 VPB VPWR 0.137f
C3 VPWR VNB 1.67f
C4 VGND VNB 1.47f
C5 VPB VNB 1.14f
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X a_369_47# a_469_47#
+ a_297_47# a_193_413# a_27_47#
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPWR B 0.0186f
C1 C X 0.00479f
C2 a_369_47# VGND 0.00505f
C3 VPWR VGND 0.0727f
C4 a_27_47# a_193_413# 0.125f
C5 C a_469_47# 0.00202f
C6 a_27_47# B 0.0794f
C7 a_193_413# a_297_47# 0.00137f
C8 a_27_47# VGND 0.103f
C9 VPB D 0.0763f
C10 X a_193_413# 0.108f
C11 VPWR VPB 0.0818f
C12 B a_297_47# 0.00353f
C13 VPWR D 0.0186f
C14 a_297_47# VGND 0.00183f
C15 VPWR a_369_47# 6.65e-19
C16 X VGND 0.0588f
C17 a_193_413# a_469_47# 0.00109f
C18 VPB a_27_47# 0.092f
C19 a_469_47# VGND 0.00551f
C20 C a_193_413# 0.0389f
C21 VPWR a_27_47# 0.106f
C22 A_N a_193_413# 0.00151f
C23 VPB X 0.0108f
C24 D X 0.0168f
C25 B C 0.164f
C26 VPWR a_297_47# 2.82e-19
C27 C VGND 0.0395f
C28 VPWR X 0.0586f
C29 A_N VGND 0.0205f
C30 D a_469_47# 0.00183f
C31 VPWR a_469_47# 7.77e-19
C32 B a_193_413# 0.144f
C33 a_193_413# VGND 0.0915f
C34 VPB C 0.0742f
C35 D C 0.183f
C36 VPB A_N 0.0832f
C37 B VGND 0.037f
C38 C a_369_47# 0.00448f
C39 VPWR C 0.0182f
C40 VPWR A_N 0.02f
C41 VPB a_193_413# 0.0644f
C42 X a_469_47# 0.001f
C43 D a_193_413# 0.155f
C44 a_193_413# a_369_47# 0.00181f
C45 A_N a_27_47# 0.237f
C46 VPWR a_193_413# 0.281f
C47 VPB B 0.089f
C48 VPB VGND 0.0123f
C49 D VGND 0.0372f
C50 B a_369_47# 0.00129f
C51 VGND VNB 0.456f
C52 X VNB 0.0934f
C53 VPWR VNB 0.368f
C54 D VNB 0.123f
C55 C VNB 0.108f
C56 B VNB 0.12f
C57 A_N VNB 0.198f
C58 VPB VNB 0.782f
C59 a_193_413# VNB 0.136f
C60 a_27_47# VNB 0.224f
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X a_109_93# a_368_53# a_209_311#
+ a_296_53#
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
C0 VPWR X 0.0732f
C1 B A_N 2.03e-19
C2 VGND VPB 0.00909f
C3 B C 0.0671f
C4 A_N X 1.44e-19
C5 B a_109_93# 0.0802f
C6 C X 0.0176f
C7 B VPB 0.0914f
C8 a_296_53# VGND 6.07e-19
C9 X VPB 0.0119f
C10 VPWR a_209_311# 0.155f
C11 a_368_53# VGND 0.0031f
C12 a_209_311# A_N 0.00515f
C13 VPWR A_N 0.0513f
C14 B VGND 0.00796f
C15 a_209_311# C 0.19f
C16 VPWR C 0.005f
C17 a_109_93# a_209_311# 0.168f
C18 X VGND 0.0647f
C19 VPWR a_109_93# 0.0984f
C20 a_209_311# VPB 0.0515f
C21 C A_N 7.6e-19
C22 VPWR VPB 0.104f
C23 a_109_93# A_N 0.117f
C24 A_N VPB 0.111f
C25 B X 0.00119f
C26 a_109_93# C 3.91e-20
C27 C VPB 0.0339f
C28 a_296_53# a_209_311# 0.0049f
C29 VPWR a_296_53# 1.15e-19
C30 a_109_93# VPB 0.0652f
C31 a_209_311# VGND 0.131f
C32 a_368_53# a_209_311# 0.0026f
C33 VPWR VGND 0.0657f
C34 a_368_53# VPWR 4.26e-19
C35 A_N VGND 0.045f
C36 B a_209_311# 0.0609f
C37 C VGND 0.0678f
C38 VPWR B 0.131f
C39 a_368_53# C 0.00415f
C40 a_296_53# a_109_93# 1.84e-19
C41 a_209_311# X 0.0877f
C42 a_109_93# VGND 0.0784f
C43 VGND VNB 0.44f
C44 X VNB 0.0925f
C45 C VNB 0.114f
C46 B VNB 0.101f
C47 VPWR VNB 0.342f
C48 A_N VNB 0.197f
C49 VPB VNB 0.693f
C50 a_209_311# VNB 0.143f
C51 a_109_93# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
C0 a_27_47# X 0.328f
C1 X VPB 0.0122f
C2 VGND A 0.0431f
C3 X VPWR 0.317f
C4 VGND a_27_47# 0.148f
C5 a_27_47# A 0.195f
C6 VGND VPB 0.00583f
C7 VPB A 0.0321f
C8 VGND VPWR 0.057f
C9 VPWR A 0.022f
C10 a_27_47# VPB 0.139f
C11 a_27_47# VPWR 0.219f
C12 VGND X 0.216f
C13 VPWR VPB 0.0632f
C14 X A 0.014f
C15 VGND VNB 0.358f
C16 X VNB 0.067f
C17 VPWR VNB 0.308f
C18 A VNB 0.148f
C19 VPB VNB 0.605f
C20 a_27_47# VNB 0.543f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
C0 a_59_75# A 0.0809f
C1 a_59_75# a_145_75# 0.00658f
C2 a_59_75# VGND 0.116f
C3 X VPWR 0.111f
C4 B VPB 0.0629f
C5 A VPWR 0.0362f
C6 a_145_75# VPWR 6.31e-19
C7 VGND VPWR 0.0461f
C8 B a_59_75# 0.143f
C9 X A 1.68e-19
C10 a_59_75# VPB 0.0563f
C11 X a_145_75# 5.76e-19
C12 X VGND 0.0993f
C13 B VPWR 0.0117f
C14 VGND A 0.0147f
C15 VPWR VPB 0.0729f
C16 VGND a_145_75# 0.00468f
C17 B X 0.00276f
C18 X VPB 0.0127f
C19 a_59_75# VPWR 0.15f
C20 B A 0.0971f
C21 A VPB 0.0806f
C22 X a_59_75# 0.109f
C23 B VGND 0.0115f
C24 VGND VPB 0.008f
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y a_297_297# a_191_297#
+ a_109_297#
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
C0 A C 0.00268f
C1 B VPWR 0.0887f
C2 VGND D 0.0456f
C3 B VPB 0.0304f
C4 A Y 0.0175f
C5 C VPWR 0.0509f
C6 VPB C 0.0299f
C7 Y VPWR 0.0561f
C8 VPB Y 0.0127f
C9 a_297_297# VGND 8.1e-19
C10 a_109_297# VPWR 0.00576f
C11 VPWR D 0.0128f
C12 B a_191_297# 0.00223f
C13 VPB D 0.0376f
C14 a_191_297# C 0.0195f
C15 A a_297_297# 3.16e-19
C16 B C 0.173f
C17 A VGND 0.0526f
C18 a_191_297# Y 0.00142f
C19 B Y 0.0403f
C20 a_297_297# VPWR 0.00317f
C21 VPWR VGND 0.0492f
C22 VPB VGND 0.0048f
C23 Y C 0.125f
C24 a_109_297# C 0.0062f
C25 C D 0.0523f
C26 A VPWR 0.0483f
C27 a_109_297# Y 0.0122f
C28 A VPB 0.041f
C29 Y D 0.108f
C30 B a_297_297# 0.0132f
C31 a_191_297# VGND 9.29e-19
C32 VPB VPWR 0.0524f
C33 B VGND 0.0191f
C34 C VGND 0.0184f
C35 a_297_297# Y 1.24e-19
C36 Y VGND 0.151f
C37 B A 0.11f
C38 a_109_297# VGND 0.00181f
C39 a_191_297# VPWR 0.0049f
C40 VGND VNB 0.322f
C41 VPWR VNB 0.276f
C42 Y VNB 0.0645f
C43 A VNB 0.174f
C44 B VNB 0.0968f
C45 C VNB 0.0911f
C46 D VNB 0.159f
C47 VPB VNB 0.516f
.ends

.subckt sky130_fd_pr__nfet_01v8_2V6S9N a_n216_n42# a_158_n42# a_n158_n130# a_n284_n216#
X0 a_158_n42# a_n158_n130# a_n216_n42# a_n284_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.58
C0 a_n158_n130# a_n216_n42# 0.018f
C1 a_n216_n42# a_158_n42# 0.0165f
C2 a_n158_n130# a_158_n42# 0.018f
C3 a_158_n42# a_n284_n216# 0.0746f
C4 a_n216_n42# a_n284_n216# 0.0746f
C5 a_n158_n130# a_n284_n216# 0.981f
.ends

.subckt sky130_fd_pr__pfet_01v8_XYZSMQ a_n33_n255# a_15_n158# w_n211_n377# a_n73_n158#
+ VSUBS
X0 a_15_n158# a_n33_n255# a_n73_n158# w_n211_n377# sky130_fd_pr__pfet_01v8 ad=0.458 pd=3.74 as=0.458 ps=3.74 w=1.58 l=0.15
C0 w_n211_n377# a_n33_n255# 0.191f
C1 w_n211_n377# a_15_n158# 0.0299f
C2 a_n33_n255# a_n73_n158# 0.0271f
C3 a_15_n158# a_n73_n158# 0.254f
C4 a_15_n158# a_n33_n255# 0.0271f
C5 w_n211_n377# a_n73_n158# 0.0299f
C6 a_15_n158# VSUBS 0.132f
C7 a_n73_n158# VSUBS 0.132f
C8 a_n33_n255# VSUBS 0.146f
C9 w_n211_n377# VSUBS 1.04f
.ends

.subckt sky130_fd_pr__pfet_01v8_AZD9DW w_n353_n261# a_n157_n139# a_n215_n42# a_157_n42#
+ VSUBS
X0 a_157_n42# a_n157_n139# a_n215_n42# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.57
C0 w_n353_n261# a_n157_n139# 0.396f
C1 w_n353_n261# a_157_n42# 0.0323f
C2 a_n157_n139# a_n215_n42# 0.0179f
C3 a_157_n42# a_n215_n42# 0.0166f
C4 a_157_n42# a_n157_n139# 0.0179f
C5 w_n353_n261# a_n215_n42# 0.0179f
C6 a_157_n42# VSUBS 0.0468f
C7 a_n215_n42# VSUBS 0.0559f
C8 a_n157_n139# VSUBS 0.569f
C9 w_n353_n261# VSUBS 1.17f
.ends

.subckt sky130_fd_pr__nfet_01v8_T8HSQ7 a_n175_n297# a_15_n157# a_n33_n245# a_n73_n157#
X0 a_15_n157# a_n33_n245# a_n73_n157# a_n175_n297# sky130_fd_pr__nfet_01v8 ad=0.455 pd=3.72 as=0.455 ps=3.72 w=1.57 l=0.15
C0 a_n33_n245# a_n73_n157# 0.0289f
C1 a_n73_n157# a_15_n157# 0.253f
C2 a_n33_n245# a_15_n157# 0.0289f
C3 a_15_n157# a_n175_n297# 0.161f
C4 a_n73_n157# a_n175_n297# 0.188f
C5 a_n33_n245# a_n175_n297# 0.322f
.ends

.subckt th09 V09 Vin Vn m1_485_n505# Vp m1_962_372#
XXM0 m1_485_n505# Vn Vin Vn sky130_fd_pr__nfet_01v8_2V6S9N
XXM1 Vin m1_485_n505# Vp Vp Vn sky130_fd_pr__pfet_01v8_XYZSMQ
XXM2 Vp m1_485_n505# Vp m1_962_372# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM3 Vp m1_485_n505# V09 m1_962_372# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM4 Vn V09 m1_485_n505# Vn sky130_fd_pr__nfet_01v8_T8HSQ7
C0 Vn Vin 0.0386f
C1 Vn V09 0.00364f
C2 V09 Vin 2.77e-19
C3 Vn m1_962_372# 6.71e-21
C4 m1_485_n505# Vn 0.0846f
C5 Vin m1_962_372# 0.00821f
C6 m1_485_n505# Vin 0.372f
C7 Vn Vp 0.0176f
C8 Vin Vp 0.187f
C9 V09 m1_962_372# 0.00205f
C10 m1_485_n505# V09 0.104f
C11 V09 Vp 0.0743f
C12 m1_485_n505# m1_962_372# 0.0822f
C13 Vp m1_962_372# 0.0579f
C14 m1_485_n505# Vp 0.372f
C15 Vin 0 1.1f
C16 m1_485_n505# 0 1.18f
C17 V09 0 0.27f
C18 Vn 0 0.344f
C19 m1_962_372# 0 0.118f
C20 Vp 0 3.27f
.ends

.subckt sky130_fd_pr__pfet_01v8_HPNF99 a_n33_n147# a_23_n50# a_n81_n50# w_n219_n269#
+ VSUBS
X0 a_23_n50# a_n33_n147# a_n81_n50# w_n219_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.23
C0 a_n81_n50# a_23_n50# 0.07f
C1 a_23_n50# w_n219_n269# 0.0185f
C2 a_n81_n50# w_n219_n269# 0.0419f
C3 a_23_n50# a_n33_n147# 0.00814f
C4 a_n81_n50# a_n33_n147# 0.00814f
C5 w_n219_n269# a_n33_n147# 0.173f
C6 a_23_n50# VSUBS 0.0578f
C7 a_n81_n50# VSUBS 0.0428f
C8 a_n33_n147# VSUBS 0.157f
C9 w_n219_n269# VSUBS 0.779f
.ends

.subckt sky130_fd_pr__nfet_01v8_JZU22M a_n213_n42# a_155_n42# a_n155_n130# a_281_n238#
X0 a_155_n42# a_n155_n130# a_n213_n42# a_281_n238# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.55
C0 a_155_n42# a_n155_n130# 0.0178f
C1 a_155_n42# a_n213_n42# 0.0168f
C2 a_n155_n130# a_n213_n42# 0.0178f
C3 a_155_n42# a_281_n238# 0.0816f
C4 a_n213_n42# a_281_n238# 0.0737f
C5 a_n155_n130# a_281_n238# 0.928f
.ends

.subckt sky130_fd_pr__pfet_01v8_TM5S5A a_n80_n147# a_n138_n50# a_80_n50# w_n276_n269#
+ VSUBS
X0 a_80_n50# a_n80_n147# a_n138_n50# w_n276_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.8
C0 a_n138_n50# a_80_n50# 0.0335f
C1 a_80_n50# w_n276_n269# 0.0231f
C2 a_n138_n50# w_n276_n269# 0.0231f
C3 a_80_n50# a_n80_n147# 0.0141f
C4 a_n138_n50# a_n80_n147# 0.0141f
C5 w_n276_n269# a_n80_n147# 0.297f
C6 a_80_n50# VSUBS 0.0565f
C7 a_n138_n50# VSUBS 0.0565f
C8 a_n80_n147# VSUBS 0.296f
C9 w_n276_n269# VSUBS 1.01f
.ends

.subckt sky130_fd_pr__pfet_01v8_AM8GZ5 w_n526_n261# a_n330_n139# a_330_n42# a_n388_n42#
+ VSUBS
X0 a_330_n42# a_n330_n139# a_n388_n42# w_n526_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.3
C0 a_n388_n42# a_330_n42# 0.00853f
C1 a_330_n42# w_n526_n261# 0.0408f
C2 a_n388_n42# w_n526_n261# 0.0179f
C3 a_330_n42# a_n330_n139# 0.0223f
C4 a_n388_n42# a_n330_n139# 0.0223f
C5 w_n526_n261# a_n330_n139# 0.719f
C6 a_330_n42# VSUBS 0.0435f
C7 a_n388_n42# VSUBS 0.0585f
C8 a_n330_n139# VSUBS 1.13f
C9 w_n526_n261# VSUBS 1.76f
.ends

.subckt sky130_fd_pr__nfet_01v8_H7HSAV a_n73_n250# a_15_n250# a_n33_n338# a_n141_n424#
X0 a_15_n250# a_n33_n338# a_n73_n250# a_n141_n424# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.15
C0 a_15_n250# a_n33_n338# 0.0337f
C1 a_15_n250# a_n73_n250# 0.401f
C2 a_n33_n338# a_n73_n250# 0.0337f
C3 a_15_n250# a_n141_n424# 0.24f
C4 a_n73_n250# a_n141_n424# 0.24f
C5 a_n33_n338# a_n141_n424# 0.327f
.ends

.subckt th14 V14 Vin Vn m1_641_n318# Vp m1_891_419#
XXM0 Vn Vn m1_641_n318# Vp Vn sky130_fd_pr__pfet_01v8_HPNF99
XXM1 m1_641_n318# m1_891_419# Vin Vn sky130_fd_pr__nfet_01v8_JZU22M
XXM2 Vin Vp m1_891_419# Vp Vn sky130_fd_pr__pfet_01v8_TM5S5A
XXM3 Vp m1_891_419# V14 Vp Vn sky130_fd_pr__pfet_01v8_AM8GZ5
XXM4 Vn V14 m1_891_419# Vn sky130_fd_pr__nfet_01v8_H7HSAV
C0 V14 Vp 0.082f
C1 m1_641_n318# m1_891_419# 0.00289f
C2 Vin Vp 0.201f
C3 V14 Vin 0.00516f
C4 m1_641_n318# Vp 0.0629f
C5 m1_891_419# Vp 0.227f
C6 V14 m1_891_419# 0.249f
C7 m1_641_n318# Vin 0.229f
C8 Vin m1_891_419# 0.132f
C9 m1_891_419# Vn 1.7f
C10 V14 Vn 0.273f
C11 Vp Vn 3.39f
C12 Vin Vn 1.76f
C13 m1_641_n318# Vn 0.313f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X a_75_212#
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 VPWR a_75_212# 0.134f
C1 VPWR A 0.0217f
C2 A a_75_212# 0.178f
C3 VPWR VPB 0.0355f
C4 a_75_212# VPB 0.0571f
C5 VPWR X 0.0896f
C6 a_75_212# X 0.107f
C7 VPWR VGND 0.0289f
C8 VGND a_75_212# 0.105f
C9 A VPB 0.0525f
C10 A X 8.48e-19
C11 VPB X 0.0128f
C12 VGND A 0.0184f
C13 VGND VPB 0.00507f
C14 VGND X 0.0545f
C15 VGND VNB 0.207f
C16 VPWR VNB 0.176f
C17 X VNB 0.0942f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_75_212# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 X a_27_47# 0.107f
C1 X A 8.48e-19
C2 A a_27_47# 0.181f
C3 X VPB 0.0128f
C4 a_27_47# VPB 0.0592f
C5 X VPWR 0.0897f
C6 a_27_47# VPWR 0.135f
C7 X VGND 0.0546f
C8 VGND a_27_47# 0.105f
C9 A VPB 0.0524f
C10 A VPWR 0.0215f
C11 VPB VPWR 0.0355f
C12 VGND A 0.0184f
C13 VGND VPB 0.00505f
C14 VGND VPWR 0.029f
C15 VGND VNB 0.207f
C16 X VNB 0.0941f
C17 VPWR VNB 0.175f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_27_47# VNB 0.208f
.ends

.subckt sky130_fd_pr__pfet_01v8_P28Q2U a_n33_n232# a_15_n135# w_n211_n354# a_n73_n135#
+ VSUBS
X0 a_15_n135# a_n33_n232# a_n73_n135# w_n211_n354# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.28 as=0.391 ps=3.28 w=1.35 l=0.15
C0 w_n211_n354# a_n73_n135# 0.0279f
C1 w_n211_n354# a_n33_n232# 0.19f
C2 w_n211_n354# a_15_n135# 0.0279f
C3 a_n73_n135# a_n33_n232# 0.0258f
C4 a_n73_n135# a_15_n135# 0.218f
C5 a_n33_n232# a_15_n135# 0.0258f
C6 a_15_n135# VSUBS 0.115f
C7 a_n73_n135# VSUBS 0.115f
C8 a_n33_n232# VSUBS 0.146f
C9 w_n211_n354# VSUBS 0.983f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZMY3VB a_n348_n42# a_n290_n130# a_n450_n182# a_290_n42#
X0 a_290_n42# a_n290_n130# a_n348_n42# a_n450_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.9
C0 a_n290_n130# a_290_n42# 0.0217f
C1 a_n290_n130# a_n348_n42# 0.0217f
C2 a_290_n42# a_n348_n42# 0.00961f
C3 a_290_n42# a_n450_n182# 0.076f
C4 a_n348_n42# a_n450_n182# 0.0839f
C5 a_n290_n130# a_n450_n182# 1.6f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 w_n211_n319# a_n73_n100# 0.0248f
C1 w_n211_n319# a_n33_n197# 0.189f
C2 w_n211_n319# a_15_n100# 0.0248f
C3 a_n73_n100# a_n33_n197# 0.0236f
C4 a_n73_n100# a_15_n100# 0.162f
C5 a_n33_n197# a_15_n100# 0.0236f
C6 a_15_n100# VSUBS 0.0885f
C7 a_n73_n100# VSUBS 0.0885f
C8 a_n33_n197# VSUBS 0.145f
C9 w_n211_n319# VSUBS 0.894f
.ends

.subckt sky130_fd_pr__pfet_01v8_WV9GCW a_n158_n42# w_n296_n261# a_n100_n139# a_100_n42#
+ VSUBS
X0 a_100_n42# a_n100_n139# a_n158_n42# w_n296_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1
C0 w_n296_n261# a_n158_n42# 0.0224f
C1 w_n296_n261# a_n100_n139# 0.346f
C2 w_n296_n261# a_100_n42# 0.0224f
C3 a_n158_n42# a_n100_n139# 0.0144f
C4 a_n158_n42# a_100_n42# 0.024f
C5 a_n100_n139# a_100_n42# 0.0144f
C6 a_100_n42# VSUBS 0.0504f
C7 a_n158_n42# VSUBS 0.0504f
C8 a_n100_n139# VSUBS 0.353f
C9 w_n296_n261# VSUBS 1.06f
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n141_240# a_n33_n188# a_15_n100#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n141_240# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n33_n188# a_15_n100# 0.0254f
C1 a_n33_n188# a_n73_n100# 0.0254f
C2 a_15_n100# a_n73_n100# 0.162f
C3 a_15_n100# a_n141_240# 0.113f
C4 a_n73_n100# a_n141_240# 0.113f
C5 a_n33_n188# a_n141_240# 0.322f
.ends

.subckt th12 V12 Vin m1_394_n856# m1_529_n42# Vp Vn
XXM0 Vn Vn Vp m1_394_n856# Vn sky130_fd_pr__pfet_01v8_P28Q2U
XXM1 m1_529_n42# Vin Vn m1_394_n856# sky130_fd_pr__nfet_01v8_ZMY3VB
XXM2 m1_529_n42# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM3 Vp Vp m1_529_n42# V12 Vn sky130_fd_pr__pfet_01v8_WV9GCW
XXM4 V12 Vn m1_529_n42# Vn sky130_fd_pr__nfet_01v8_648S5X
C0 m1_394_n856# Vp 0.04f
C1 m1_529_n42# Vp 0.322f
C2 m1_394_n856# Vn 0.0338f
C3 m1_529_n42# Vn 0.254f
C4 V12 Vp 0.0454f
C5 V12 Vn 0.0234f
C6 Vin Vp 0.238f
C7 Vin Vn 0.135f
C8 m1_394_n856# m1_529_n42# 0.0134f
C9 m1_394_n856# V12 4.74e-19
C10 V12 m1_529_n42# 0.0929f
C11 Vp Vn 0.132f
C12 Vin m1_394_n856# 0.321f
C13 Vin m1_529_n42# 0.0965f
C14 Vin V12 0.00205f
C15 Vn 0 0.29f
C16 Vp 0 2.88f
C17 m1_529_n42# 0 0.861f
C18 V12 0 0.359f
C19 Vin 0 1.9f
C20 m1_394_n856# 0 0.215f
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X a_664_47# a_841_47#
+ a_381_47# a_62_47# a_558_47#
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPB a_841_47# 0.0108f
C1 VPB a_381_47# 0.0447f
C2 VPB X 0.126f
C3 VPB a_62_47# 0.0515f
C4 VPB A 0.105f
C5 X a_381_47# 0.318f
C6 VPB VPWR 0.103f
C7 A a_381_47# 5.42e-19
C8 a_62_47# X 0.156f
C9 VPWR a_841_47# 0.0614f
C10 VPB VGND 0.008f
C11 X A 0.0142f
C12 VGND a_841_47# 0.0585f
C13 a_664_47# VPB 0.043f
C14 a_664_47# a_841_47# 0.134f
C15 a_62_47# A 0.244f
C16 VPWR a_381_47# 0.134f
C17 VPB a_558_47# 0.115f
C18 VGND a_381_47# 0.125f
C19 a_558_47# a_841_47# 0.00368f
C20 X VPWR 0.108f
C21 X VGND 0.106f
C22 a_664_47# X 6.67e-19
C23 a_62_47# VPWR 0.149f
C24 VPWR A 0.0174f
C25 a_62_47# VGND 0.144f
C26 a_558_47# a_381_47# 0.16f
C27 VGND A 0.0176f
C28 a_558_47# X 0.0144f
C29 VPWR VGND 0.0902f
C30 a_664_47# VPWR 0.131f
C31 a_664_47# VGND 0.125f
C32 a_558_47# VPWR 0.084f
C33 a_558_47# VGND 0.0816f
C34 a_664_47# a_558_47# 0.314f
C35 VGND VNB 0.537f
C36 VPWR VNB 0.439f
C37 X VNB 0.163f
C38 A VNB 0.198f
C39 VPB VNB 0.959f
C40 a_841_47# VNB 0.0929f
C41 a_664_47# VNB 0.13f
C42 a_558_47# VNB 0.164f
C43 a_381_47# VNB 0.11f
C44 a_62_47# VNB 0.169f
.ends

.subckt sky130_fd_pr__nfet_01v8_4L9AWD a_n206_n182# a_n46_n130# a_n104_n42# a_46_n42#
X0 a_46_n42# a_n46_n130# a_n104_n42# a_n206_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.46
C0 a_46_n42# a_n46_n130# 0.00852f
C1 a_46_n42# a_n104_n42# 0.0412f
C2 a_n46_n130# a_n104_n42# 0.00852f
C3 a_46_n42# a_n206_n182# 0.0705f
C4 a_n104_n42# a_n206_n182# 0.0784f
C5 a_n46_n130# a_n206_n182# 0.388f
.ends

.subckt sky130_fd_pr__pfet_01v8_EZD9Q7 w_n224_n261# a_28_n42# a_n33_n139# a_n86_n42#
+ VSUBS
X0 a_28_n42# a_n33_n139# a_n86_n42# w_n224_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.28
C0 a_28_n42# w_n224_n261# 0.0224f
C1 a_28_n42# a_n33_n139# 0.00625f
C2 a_n86_n42# w_n224_n261# 0.0224f
C3 a_n86_n42# a_n33_n139# 0.00625f
C4 w_n224_n261# a_n33_n139# 0.183f
C5 a_n86_n42# a_28_n42# 0.0541f
C6 a_28_n42# VSUBS 0.0479f
C7 a_n86_n42# VSUBS 0.0479f
C8 a_n33_n139# VSUBS 0.155f
C9 w_n224_n261# VSUBS 0.799f
.ends

.subckt sky130_fd_pr__pfet_01v8_M479BZ a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_15_n42# w_n211_n261# 0.0389f
C1 a_15_n42# a_n33_n139# 0.0192f
C2 a_n73_n42# w_n211_n261# 0.016f
C3 a_n73_n42# a_n33_n139# 0.0192f
C4 w_n211_n261# a_n33_n139# 0.182f
C5 a_n73_n42# a_15_n42# 0.0699f
C6 a_15_n42# VSUBS 0.0328f
C7 a_n73_n42# VSUBS 0.0478f
C8 a_n33_n139# VSUBS 0.145f
C9 w_n211_n261# VSUBS 0.785f
.ends

.subckt sky130_fd_pr__nfet_01v8_4BNSKG a_n144_n216# a_18_n42# a_n33_n130# a_n76_n42#
X0 a_18_n42# a_n33_n130# a_n76_n42# a_n144_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.18
C0 a_18_n42# a_n33_n130# 0.0154f
C1 a_18_n42# a_n76_n42# 0.0655f
C2 a_n33_n130# a_n76_n42# 0.0154f
C3 a_18_n42# a_n144_n216# 0.0668f
C4 a_n76_n42# a_n144_n216# 0.0668f
C5 a_n33_n130# a_n144_n216# 0.319f
.ends

.subckt th10 V10 Vin m1_502_n495# m1_536_174# Vn Vp
XXM0 m1_502_n495# Vn Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vn Vin m1_536_174# m1_502_n495# sky130_fd_pr__nfet_01v8_4L9AWD
XXM2 Vp m1_536_174# Vin Vp Vn sky130_fd_pr__pfet_01v8_EZD9Q7
XXM3 Vp Vp m1_536_174# V10 Vn sky130_fd_pr__pfet_01v8_M479BZ
XXM4 Vn V10 m1_536_174# Vn sky130_fd_pr__nfet_01v8_4BNSKG
C0 Vin V10 0.0187f
C1 m1_502_n495# V10 0.042f
C2 Vp m1_536_174# 0.172f
C3 Vin m1_502_n495# 0.0207f
C4 Vp Vn 0.102f
C5 Vn m1_536_174# 0.233f
C6 Vp V10 0.0702f
C7 m1_536_174# V10 0.177f
C8 Vin Vp 0.175f
C9 m1_502_n495# Vp 0.0256f
C10 Vin m1_536_174# 0.0971f
C11 m1_502_n495# m1_536_174# 0.00612f
C12 Vn V10 0.0577f
C13 Vin Vn 0.114f
C14 m1_502_n495# Vn 0.0348f
C15 Vin 0 0.664f
C16 V10 0 0.249f
C17 Vn 0 0.463f
C18 m1_536_174# 0 0.825f
C19 Vp 0 2.17f
C20 m1_502_n495# 0 0.146f
.ends

.subckt sky130_fd_pr__nfet_01v8_X33H33 a_n73_n110# a_n175_n250# a_n33_n198# a_15_n110#
X0 a_15_n110# a_n33_n198# a_n73_n110# a_n175_n250# sky130_fd_pr__nfet_01v8 ad=0.319 pd=2.78 as=0.319 ps=2.78 w=1.1 l=0.15
C0 a_n33_n198# a_15_n110# 0.0261f
C1 a_15_n110# a_n73_n110# 0.178f
C2 a_n33_n198# a_n73_n110# 0.0261f
C3 a_15_n110# a_n175_n250# 0.121f
C4 a_n73_n110# a_n175_n250# 0.141f
C5 a_n33_n198# a_n175_n250# 0.32f
.ends

.subckt sky130_fd_pr__pfet_01v8_AMA9E4 a_n194_n44# a_n136_n141# w_n332_n263# a_136_n44#
+ VSUBS
X0 a_136_n44# a_n136_n141# a_n194_n44# w_n332_n263# sky130_fd_pr__pfet_01v8 ad=0.128 pd=1.46 as=0.128 ps=1.46 w=0.44 l=1.36
C0 a_136_n44# a_n194_n44# 0.0196f
C1 w_n332_n263# a_n194_n44# 0.0226f
C2 a_136_n44# w_n332_n263# 0.0226f
C3 a_n194_n44# a_n136_n141# 0.0174f
C4 a_136_n44# a_n136_n141# 0.0174f
C5 w_n332_n263# a_n136_n141# 0.434f
C6 a_136_n44# VSUBS 0.0532f
C7 a_n194_n44# VSUBS 0.0532f
C8 a_n136_n141# VSUBS 0.457f
C9 w_n332_n263# VSUBS 1.2f
.ends

.subckt sky130_fd_pr__pfet_01v8_8DZSNJ a_n74_n100# a_16_n100# w_n212_n319# a_n33_n197#
+ VSUBS
X0 a_16_n100# a_n33_n197# a_n74_n100# w_n212_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.16
C0 a_16_n100# a_n74_n100# 0.159f
C1 w_n212_n319# a_n74_n100# 0.0252f
C2 a_16_n100# w_n212_n319# 0.0252f
C3 a_n74_n100# a_n33_n197# 0.0223f
C4 a_16_n100# a_n33_n197# 0.0223f
C5 w_n212_n319# a_n33_n197# 0.189f
C6 a_16_n100# VSUBS 0.089f
C7 a_n74_n100# VSUBS 0.089f
C8 a_n33_n197# VSUBS 0.146f
C9 w_n212_n319# VSUBS 0.899f
.ends

.subckt th03 V03 Vin Vp m1_890_n844# m1_638_n591# Vn
XXM0 Vn Vn Vin m1_890_n844# sky130_fd_pr__nfet_01v8_X33H33
XXM1 m1_638_n591# Vin Vp m1_890_n844# Vn sky130_fd_pr__pfet_01v8_AMA9E4
XXM2 Vp Vn Vp m1_638_n591# sky130_fd_pr__nfet_01v8_LH5FDA
XXM3 Vp V03 Vp m1_890_n844# Vn sky130_fd_pr__pfet_01v8_8DZSNJ
XXM4 m1_890_n844# Vn Vn V03 sky130_fd_pr__nfet_01v8_LH5FDA
C0 Vin Vn 0.105f
C1 Vp m1_638_n591# 0.169f
C2 Vp V03 0.0492f
C3 Vin m1_638_n591# 0.0439f
C4 Vin V03 0.0036f
C5 Vp Vin 0.313f
C6 Vn m1_890_n844# 0.183f
C7 m1_890_n844# m1_638_n591# 0.0187f
C8 m1_890_n844# V03 0.129f
C9 Vn m1_638_n591# 0.0097f
C10 Vp m1_890_n844# 0.459f
C11 Vn V03 0.0337f
C12 Vin m1_890_n844# 0.188f
C13 Vp Vn 0.023f
C14 Vp 0 3.07f
C15 V03 0 0.308f
C16 Vn 0 0.446f
C17 m1_890_n844# 0 1.05f
C18 m1_638_n591# 0 0.224f
C19 Vin 0 0.924f
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y a_129_47# a_47_47# a_285_47#
+ a_377_297#
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 A Y 0.00181f
C1 VPWR VPB 0.0718f
C2 VPWR a_129_47# 9.47e-19
C3 VPWR B 0.0408f
C4 a_377_297# VPWR 0.00559f
C5 a_47_47# Y 0.143f
C6 a_47_47# A 0.0307f
C7 a_285_47# VPWR 0.00255f
C8 VPB Y 0.00878f
C9 B Y 0.00334f
C10 A VPB 0.0822f
C11 a_377_297# Y 0.00188f
C12 A B 0.236f
C13 VPWR VGND 0.0665f
C14 a_285_47# Y 0.0439f
C15 a_47_47# VPB 0.0444f
C16 a_47_47# a_129_47# 0.00369f
C17 a_285_47# A 0.0353f
C18 a_47_47# B 0.356f
C19 a_377_297# a_47_47# 0.00899f
C20 VGND Y 0.0381f
C21 a_285_47# a_47_47# 0.0175f
C22 B VPB 0.0643f
C23 B a_129_47# 0.00236f
C24 A VGND 0.0635f
C25 a_377_297# B 0.00254f
C26 a_285_47# VPB 5.53e-19
C27 a_285_47# B 0.067f
C28 a_47_47# VGND 0.104f
C29 VPWR Y 0.107f
C30 VGND VPB 0.00568f
C31 a_129_47# VGND 0.00547f
C32 VPWR A 0.0349f
C33 B VGND 0.0389f
C34 a_377_297# VGND 0.00125f
C35 VPWR a_47_47# 0.273f
C36 a_285_47# VGND 0.211f
C37 VGND VNB 0.4f
C38 Y VNB 0.0783f
C39 VPWR VNB 0.352f
C40 A VNB 0.217f
C41 B VNB 0.212f
C42 VPB VNB 0.693f
C43 a_285_47# VNB 0.0174f
C44 a_47_47# VNB 0.199f
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X a_472_297# a_80_21#
+ a_300_47# a_217_297#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
C0 C1 X 7.15e-20
C1 a_300_47# X 5.31e-19
C2 VGND X 0.0654f
C3 A1 a_217_297# 0.0124f
C4 a_80_21# VPWR 0.119f
C5 A2 VPB 0.0384f
C6 B1 a_217_297# 0.00651f
C7 A1 B1 0.0834f
C8 a_80_21# A2 0.128f
C9 VPWR X 0.0884f
C10 C1 a_217_297# 0.00262f
C11 VGND a_217_297# 0.00342f
C12 A1 a_300_47# 5.95e-19
C13 VGND A1 0.0147f
C14 A2 X 6.82e-19
C15 C1 B1 0.0846f
C16 VGND B1 0.0175f
C17 VPWR a_217_297# 0.197f
C18 A1 VPWR 0.0149f
C19 VGND C1 0.0176f
C20 VGND a_300_47# 0.00536f
C21 a_80_21# a_472_297# 0.0164f
C22 A2 a_217_297# 0.0135f
C23 B1 VPWR 0.0129f
C24 A1 A2 0.0881f
C25 a_472_297# X 2.6e-19
C26 C1 VPWR 0.0137f
C27 VPWR a_300_47# 8.53e-19
C28 VGND VPWR 0.0665f
C29 VGND A2 0.0191f
C30 a_80_21# VPB 0.0661f
C31 a_472_297# a_217_297# 0.00517f
C32 VPB X 0.0118f
C33 A2 VPWR 0.0161f
C34 B1 a_472_297# 1.87e-19
C35 a_80_21# X 0.118f
C36 VGND a_472_297# 0.00188f
C37 a_217_297# VPB 0.00494f
C38 A1 VPB 0.0266f
C39 a_80_21# a_217_297# 0.127f
C40 a_472_297# VPWR 0.00703f
C41 B1 VPB 0.0267f
C42 a_80_21# A1 0.111f
C43 a_217_297# X 0.00271f
C44 C1 VPB 0.0379f
C45 a_80_21# B1 0.0964f
C46 VGND VPB 0.00775f
C47 A1 X 3.62e-19
C48 a_80_21# C1 0.079f
C49 a_80_21# a_300_47# 0.00997f
C50 a_80_21# VGND 0.293f
C51 B1 X 1.18e-19
C52 VPWR VPB 0.0754f
C53 VGND VNB 0.385f
C54 VPWR VNB 0.325f
C55 X VNB 0.0899f
C56 C1 VNB 0.144f
C57 B1 VNB 0.0899f
C58 A1 VNB 0.0905f
C59 A2 VNB 0.108f
C60 VPB VNB 0.693f
C61 a_217_297# VNB 0.00117f
C62 a_80_21# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
C0 C VPB 0.0609f
C1 a_27_47# B 0.13f
C2 VPB VGND 0.00852f
C3 C a_27_47# 0.0516f
C4 a_27_47# VGND 0.132f
C5 a_303_47# D 0.00119f
C6 X D 0.00746f
C7 VPB D 0.0782f
C8 VPWR B 0.0231f
C9 C VPWR 0.021f
C10 a_27_47# D 0.107f
C11 VPWR VGND 0.0662f
C12 a_109_47# a_27_47# 0.00578f
C13 A VPB 0.0907f
C14 VPB X 0.0111f
C15 a_27_47# a_197_47# 0.00167f
C16 a_303_47# a_27_47# 0.00119f
C17 A a_27_47# 0.153f
C18 a_27_47# X 0.0754f
C19 C B 0.161f
C20 VGND B 0.0453f
C21 VPWR D 0.0207f
C22 a_109_47# VPWR 4.66e-19
C23 C VGND 0.0408f
C24 a_27_47# VPB 0.082f
C25 a_197_47# VPWR 5.24e-19
C26 a_303_47# VPWR 4.83e-19
C27 A VPWR 0.044f
C28 VPWR X 0.0945f
C29 a_109_47# B 0.00153f
C30 C D 0.18f
C31 VGND D 0.0898f
C32 a_197_47# B 0.00623f
C33 VPWR VPB 0.077f
C34 C a_109_47# 1.72e-20
C35 a_109_47# VGND 0.00223f
C36 C a_197_47# 0.00123f
C37 A B 0.0839f
C38 a_27_47# VPWR 0.326f
C39 a_197_47# VGND 0.00387f
C40 C a_303_47# 0.00527f
C41 a_303_47# VGND 0.00381f
C42 A VGND 0.0151f
C43 VGND X 0.0903f
C44 VPB B 0.0643f
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt sky130_fd_pr__nfet_01v8_SHU4BF a_n73_n353# a_n141_493# a_15_n353# a_n33_n441#
X0 a_15_n353# a_n33_n441# a_n73_n353# a_n141_493# sky130_fd_pr__nfet_01v8 ad=1.02 pd=7.64 as=1.02 ps=7.64 w=3.53 l=0.15
C0 a_n73_n353# a_n33_n441# 0.0384f
C1 a_15_n353# a_n33_n441# 0.0384f
C2 a_n73_n353# a_15_n353# 0.564f
C3 a_15_n353# a_n141_493# 0.327f
C4 a_n73_n353# a_n141_493# 0.327f
C5 a_n33_n441# a_n141_493# 0.329f
.ends

.subckt sky130_fd_pr__pfet_01v8_HE9GT9 a_n408_n42# a_350_n42# w_n546_n261# a_n350_n139#
+ VSUBS
X0 a_350_n42# a_n350_n139# a_n408_n42# w_n546_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 a_350_n42# w_n546_n261# 0.0179f
C1 a_n350_n139# a_350_n42# 0.0226f
C2 a_n350_n139# w_n546_n261# 0.756f
C3 a_350_n42# a_n408_n42# 0.00807f
C4 a_n408_n42# w_n546_n261# 0.0408f
C5 a_n350_n139# a_n408_n42# 0.0226f
C6 a_350_n42# VSUBS 0.0587f
C7 a_n408_n42# VSUBS 0.0437f
C8 a_n350_n139# VSUBS 1.19f
C9 w_n546_n261# VSUBS 1.83f
.ends

.subckt sky130_fd_pr__nfet_01v8_LHD8GA a_n408_n42# a_350_n42# a_n350_n130# a_n510_n182#
X0 a_350_n42# a_n350_n130# a_n408_n42# a_n510_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 a_n408_n42# a_n350_n130# 0.0226f
C1 a_350_n42# a_n350_n130# 0.0226f
C2 a_n408_n42# a_350_n42# 0.00807f
C3 a_350_n42# a_n510_n182# 0.0766f
C4 a_n408_n42# a_n510_n182# 0.0845f
C5 a_n350_n130# a_n510_n182# 1.9f
.ends

.subckt th01 V01 Vn m1_991_n1219# m1_571_n501# Vp Vin
XXM0 Vn Vn m1_991_n1219# Vin sky130_fd_pr__nfet_01v8_SHU4BF
XXM1 m1_571_n501# m1_991_n1219# Vp Vin Vn sky130_fd_pr__pfet_01v8_HE9GT9
XXM2 Vp m1_571_n501# Vp Vn sky130_fd_pr__nfet_01v8_LHD8GA
XXM3 Vp Vp V01 m1_991_n1219# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_991_n1219# Vn V01 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 m1_991_n1219# Vn 0.0569f
C1 Vin V01 0.00412f
C2 m1_571_n501# Vin 0.274f
C3 Vp m1_991_n1219# 0.423f
C4 Vin Vn 0.0582f
C5 Vin Vp 0.354f
C6 Vin m1_991_n1219# 0.208f
C7 m1_571_n501# V01 2.16e-20
C8 V01 Vn 0.0149f
C9 m1_571_n501# Vn 2.57e-20
C10 Vp V01 0.0684f
C11 m1_571_n501# Vp 0.32f
C12 Vp Vn 0.0233f
C13 m1_991_n1219# V01 0.0901f
C14 m1_571_n501# m1_991_n1219# 0.0899f
C15 Vn 0 0.633f
C16 V01 0 0.373f
C17 m1_991_n1219# 0 1.24f
C18 Vp 0 4.41f
C19 m1_571_n501# 0 0.194f
C20 Vin 0 1.87f
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X a_489_413# a_226_47#
+ a_556_47# a_226_297# a_76_199#
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_76_199# a_226_47# 0.188f
C1 X a_76_199# 0.0995f
C2 VGND a_226_47# 0.149f
C3 X VGND 0.0627f
C4 VPWR a_226_297# 8.54e-19
C5 a_489_413# a_226_47# 0.00579f
C6 A2_N a_226_47# 0.141f
C7 X A2_N 2.55e-19
C8 a_226_297# a_76_199# 0.00354f
C9 A1_N VPB 0.0339f
C10 B2 VPB 0.0645f
C11 a_556_47# B2 0.00291f
C12 X a_226_47# 0.0108f
C13 a_226_297# VGND 5.63e-19
C14 B1 B2 0.182f
C15 VPWR A1_N 0.00672f
C16 VPWR B2 0.0161f
C17 B1 VPB 0.0803f
C18 A1_N a_76_199# 0.119f
C19 VPWR VPB 0.0951f
C20 a_226_297# a_226_47# 0.00128f
C21 a_76_199# B2 0.0626f
C22 VPWR a_556_47# 7.24e-19
C23 VGND A1_N 0.0261f
C24 VPWR B1 0.0188f
C25 a_76_199# VPB 0.0817f
C26 a_76_199# a_556_47# 0.0017f
C27 VGND B2 0.0335f
C28 A2_N A1_N 0.11f
C29 B1 a_76_199# 0.00185f
C30 a_489_413# B2 0.0541f
C31 VGND VPB 0.0128f
C32 VGND a_556_47# 0.00639f
C33 VPWR a_76_199# 0.2f
C34 a_489_413# VPB 0.015f
C35 A1_N a_226_47# 0.0209f
C36 VGND B1 0.0471f
C37 A2_N VPB 0.0327f
C38 X A1_N 0.00211f
C39 a_489_413# B1 0.0382f
C40 B2 a_226_47# 0.0975f
C41 VPWR VGND 0.0743f
C42 VPWR a_489_413# 0.143f
C43 a_226_47# VPB 0.111f
C44 X VPB 0.0113f
C45 VPWR A2_N 0.00449f
C46 VGND a_76_199# 0.108f
C47 a_489_413# a_76_199# 0.0473f
C48 a_226_297# A1_N 0.00184f
C49 A2_N a_76_199# 0.0125f
C50 VPWR a_226_47# 0.0187f
C51 VPWR X 0.0589f
C52 VGND a_489_413# 0.0058f
C53 A2_N VGND 0.0174f
C54 VGND VNB 0.462f
C55 A2_N VNB 0.103f
C56 A1_N VNB 0.111f
C57 VPWR VNB 0.369f
C58 X VNB 0.0975f
C59 B1 VNB 0.206f
C60 B2 VNB 0.106f
C61 VPB VNB 0.782f
C62 a_489_413# VNB 0.0254f
C63 a_226_47# VNB 0.162f
C64 a_76_199# VNB 0.141f
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X a_515_93# a_223_47#
+ a_615_93# a_343_93# a_429_93# a_27_47#
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
C0 VPWR A_N 0.0318f
C1 a_223_47# A_N 0.00833f
C2 VGND a_615_93# 0.0044f
C3 a_343_93# D 0.114f
C4 VPB a_27_47# 0.154f
C5 VGND B_N 0.0427f
C6 a_343_93# C 0.0397f
C7 a_615_93# VPWR 8.49e-19
C8 a_515_93# VGND 0.00408f
C9 a_343_93# VPB 0.0857f
C10 X B_N 4.64e-20
C11 VPWR B_N 0.0168f
C12 a_223_47# B_N 0.0431f
C13 a_223_47# a_515_93# 0.00482f
C14 a_515_93# VPWR 7.86e-19
C15 VPB A_N 0.0848f
C16 a_615_93# D 0.00564f
C17 X VGND 0.0609f
C18 a_223_47# VGND 0.199f
C19 VGND VPWR 0.0906f
C20 D B_N 6.67e-20
C21 a_615_93# C 0.00407f
C22 X VPWR 0.0582f
C23 a_223_47# VPWR 0.114f
C24 B_N C 9.56e-20
C25 a_343_93# a_429_93# 0.00484f
C26 VPB B_N 0.0646f
C27 VGND D 0.0414f
C28 a_515_93# C 0.00389f
C29 VGND C 0.025f
C30 X D 0.0193f
C31 a_223_47# D 4.03e-19
C32 D VPWR 0.0143f
C33 VPB VGND 0.0167f
C34 VPWR C 0.012f
C35 a_223_47# C 0.151f
C36 X VPB 0.0103f
C37 a_223_47# VPB 0.0799f
C38 VPB VPWR 0.106f
C39 a_343_93# a_27_47# 0.0406f
C40 D C 0.163f
C41 a_27_47# A_N 0.0906f
C42 VPB D 0.081f
C43 VGND a_429_93# 0.00122f
C44 VPB C 0.0686f
C45 a_429_93# VPWR 5.19e-19
C46 a_223_47# a_429_93# 0.00492f
C47 B_N a_27_47# 0.138f
C48 a_343_93# a_615_93# 0.00103f
C49 a_343_93# B_N 0.00112f
C50 VGND a_27_47# 0.0715f
C51 a_343_93# a_515_93# 0.00115f
C52 B_N A_N 0.117f
C53 a_343_93# VGND 0.0548f
C54 VPWR a_27_47# 0.0897f
C55 a_223_47# a_27_47# 0.267f
C56 a_343_93# X 0.126f
C57 a_343_93# VPWR 0.255f
C58 a_343_93# a_223_47# 0.269f
C59 VGND A_N 0.0146f
C60 VGND VNB 0.553f
C61 X VNB 0.0908f
C62 VPWR VNB 0.453f
C63 D VNB 0.124f
C64 C VNB 0.107f
C65 B_N VNB 0.134f
C66 A_N VNB 0.144f
C67 VPB VNB 0.959f
C68 a_343_93# VNB 0.172f
C69 a_223_47# VNB 0.141f
C70 a_27_47# VNB 0.259f
.ends

.subckt sky130_fd_pr__pfet_01v8_MWHFPY a_n73_n63# a_n33_n160# w_n211_n282# a_15_n63#
+ VSUBS
X0 a_15_n63# a_n33_n160# a_n73_n63# w_n211_n282# sky130_fd_pr__pfet_01v8 ad=0.183 pd=1.84 as=0.183 ps=1.84 w=0.63 l=0.15
C0 a_n73_n63# a_15_n63# 0.103f
C1 a_15_n63# a_n33_n160# 0.021f
C2 a_n73_n63# a_n33_n160# 0.021f
C3 a_15_n63# w_n211_n282# 0.0591f
C4 a_n73_n63# w_n211_n282# 0.0591f
C5 w_n211_n282# a_n33_n160# 0.237f
C6 a_15_n63# VSUBS 0.0348f
C7 a_n73_n63# VSUBS 0.0348f
C8 a_n33_n160# VSUBS 0.116f
C9 w_n211_n282# VSUBS 1.1f
.ends

.subckt sky130_fd_pr__nfet_01v8_DPSGWY a_350_n100# a_n408_n100# a_n350_n188# a_n510_n274#
X0 a_350_n100# a_n350_n188# a_n408_n100# a_n510_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3.5
C0 a_350_n100# a_n408_n100# 0.0188f
C1 a_350_n100# a_n350_n188# 0.0439f
C2 a_n350_n188# a_n408_n100# 0.0439f
C3 a_350_n100# a_n510_n274# 0.159f
C4 a_n408_n100# a_n510_n274# 0.159f
C5 a_n350_n188# a_n510_n274# 2.13f
.ends

.subckt preamp Vin Vpamp Vn Vp
XXM0 Vn Vin Vp Vpamp Vn sky130_fd_pr__pfet_01v8_MWHFPY
XXM1 Vpamp Vp Vin Vn sky130_fd_pr__nfet_01v8_DPSGWY
C0 Vn Vp 0.297f
C1 Vpamp Vin 0.0777f
C2 Vp Vin 0.324f
C3 Vn Vin 0.29f
C4 Vpamp Vp 0.0552f
C5 Vpamp Vn 0.047f
C6 Vn 0 0.193f
C7 Vpamp 0 0.444f
C8 Vp 0 1.53f
C9 Vin 0 2.21f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 B X 0.0149f
C1 VGND A 0.0325f
C2 a_35_297# A 0.0633f
C3 VPWR a_285_47# 8.6e-19
C4 A VPB 0.051f
C5 VGND VPWR 0.0643f
C6 a_35_297# VPWR 0.096f
C7 VPWR VPB 0.0689f
C8 VGND a_285_47# 0.00552f
C9 a_35_297# a_285_47# 0.00723f
C10 A X 0.00166f
C11 VPWR a_117_297# 0.00852f
C12 a_35_297# VGND 0.177f
C13 VGND VPB 0.00696f
C14 a_35_297# VPB 0.0699f
C15 B a_285_297# 0.0553f
C16 VPWR X 0.0537f
C17 a_285_47# X 0.00206f
C18 VGND a_117_297# 0.00177f
C19 a_35_297# a_117_297# 0.00641f
C20 VGND X 0.173f
C21 a_35_297# X 0.166f
C22 X VPB 0.0154f
C23 A a_285_297# 0.00749f
C24 a_117_297# X 2.25e-19
C25 VPWR a_285_297# 0.246f
C26 A B 0.221f
C27 VPWR B 0.0703f
C28 VGND a_285_297# 0.00394f
C29 a_35_297# a_285_297# 0.025f
C30 a_285_297# VPB 0.0133f
C31 a_285_47# B 3.98e-19
C32 VGND B 0.0304f
C33 a_35_297# B 0.203f
C34 B VPB 0.0697f
C35 a_285_297# X 0.0712f
C36 a_117_297# B 0.00777f
C37 VPWR A 0.0348f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt sky130_fd_pr__pfet_01v8_LDQF7K a_n33_n147# a_29_n50# a_n87_n50# w_n225_n269#
+ VSUBS
X0 a_29_n50# a_n33_n147# a_n87_n50# w_n225_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.29
C0 a_n87_n50# w_n225_n269# 0.0457f
C1 a_29_n50# a_n87_n50# 0.0628f
C2 a_n33_n147# w_n225_n269# 0.176f
C3 a_n33_n147# a_29_n50# 0.00691f
C4 a_29_n50# w_n225_n269# 0.0186f
C5 a_n33_n147# a_n87_n50# 0.00691f
C6 a_29_n50# VSUBS 0.0581f
C7 a_n87_n50# VSUBS 0.0403f
C8 a_n33_n147# VSUBS 0.158f
C9 w_n225_n269# VSUBS 0.854f
.ends

.subckt sky130_fd_pr__nfet_01v8_HZA4VB a_326_n230# a_n200_n130# a_200_n42# li_n360_158#
+ a_n258_n42#
X0 a_200_n42# a_n200_n130# a_n258_n42# a_326_n230# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_200_n42# a_n200_n130# 0.0196f
C1 a_n258_n42# a_n200_n130# 0.0196f
C2 a_n258_n42# a_200_n42# 0.0134f
C3 li_n360_158# a_326_n230# 0.0244f
C4 a_200_n42# a_326_n230# 0.0748f
C5 a_n258_n42# a_326_n230# 0.0746f
C6 a_n200_n130# a_326_n230# 1.15f
.ends

.subckt sky130_fd_pr__pfet_01v8_GEY2B5 w_n275_n270# a_n137_n51# a_79_n51# a_n79_n148#
+ VSUBS
X0 a_79_n51# a_n79_n148# a_n137_n51# w_n275_n270# sky130_fd_pr__pfet_01v8 ad=0.148 pd=1.6 as=0.148 ps=1.6 w=0.51 l=0.79
C0 a_n137_n51# w_n275_n270# 0.0232f
C1 a_79_n51# a_n137_n51# 0.0345f
C2 a_n79_n148# w_n275_n270# 0.294f
C3 a_n79_n148# a_79_n51# 0.0141f
C4 a_79_n51# w_n275_n270# 0.0232f
C5 a_n79_n148# a_n137_n51# 0.0141f
C6 a_79_n51# VSUBS 0.0573f
C7 a_n137_n51# VSUBS 0.0573f
C8 a_n79_n148# VSUBS 0.294f
C9 w_n275_n270# VSUBS 1.01f
.ends

.subckt sky130_fd_pr__pfet_01v8_KQKFM4 w_n526_n261# a_n330_n139# a_330_n42# a_n388_n42#
+ VSUBS
X0 a_330_n42# a_n330_n139# a_n388_n42# w_n526_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.3
C0 a_n388_n42# w_n526_n261# 0.0224f
C1 a_330_n42# a_n388_n42# 0.00853f
C2 a_n330_n139# w_n526_n261# 0.911f
C3 a_n330_n139# a_330_n42# 0.0223f
C4 a_330_n42# w_n526_n261# 0.0224f
C5 a_n330_n139# a_n388_n42# 0.0223f
C6 a_330_n42# VSUBS 0.0545f
C7 a_n388_n42# VSUBS 0.0545f
C8 a_n330_n139# VSUBS 1.02f
C9 w_n526_n261# VSUBS 1.89f
.ends

.subckt sky130_fd_pr__nfet_01v8_5NW376 a_n73_n251# a_n141_391# a_15_n251# a_n33_n339#
X0 a_15_n251# a_n33_n339# a_n73_n251# a_n141_391# sky130_fd_pr__nfet_01v8 ad=0.728 pd=5.6 as=0.728 ps=5.6 w=2.51 l=0.15
C0 a_15_n251# a_n33_n339# 0.0337f
C1 a_n73_n251# a_n33_n339# 0.0337f
C2 a_n73_n251# a_15_n251# 0.402f
C3 a_15_n251# a_n141_391# 0.241f
C4 a_n73_n251# a_n141_391# 0.241f
C5 a_n33_n339# a_n141_391# 0.327f
.ends

.subckt th15 V15 Vin m1_597_n912# m1_849_n157# Vp Vn
XXM0 Vn Vn m1_597_n912# Vp Vn sky130_fd_pr__pfet_01v8_LDQF7K
XXM1 Vn Vin m1_849_n157# Vn m1_597_n912# sky130_fd_pr__nfet_01v8_HZA4VB
XXM2 Vp Vp m1_849_n157# Vin Vn sky130_fd_pr__pfet_01v8_GEY2B5
XXM3 Vp m1_849_n157# V15 Vp Vn sky130_fd_pr__pfet_01v8_KQKFM4
XXM4 Vn Vn V15 m1_849_n157# sky130_fd_pr__nfet_01v8_5NW376
C0 Vn Vp 0.0678f
C1 m1_849_n157# V15 0.202f
C2 m1_597_n912# Vin 0.211f
C3 V15 Vp 0.0762f
C4 Vn V15 2.72e-19
C5 m1_597_n912# m1_849_n157# 0.00715f
C6 m1_597_n912# Vp 0.0557f
C7 m1_597_n912# Vn 0.175f
C8 m1_849_n157# Vin 0.0977f
C9 Vin Vp 0.166f
C10 Vn Vin 0.38f
C11 V15 Vin 0.00573f
C12 m1_849_n157# Vp 0.226f
C13 m1_849_n157# Vn 0.171f
C14 V15 0 0.332f
C15 Vn 0 0.276f
C16 m1_849_n157# 0 1.28f
C17 Vp 0 3.52f
C18 m1_597_n912# 0 0.19f
C19 Vin 0 1.58f
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X a_465_297# a_297_297#
+ a_215_297# a_392_297# a_109_53#
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 VGND a_109_53# 0.118f
C1 C a_465_297# 6.89e-19
C2 VPWR a_297_297# 8.59e-19
C3 a_297_297# a_109_53# 7.06e-21
C4 B a_215_297# 0.159f
C5 A VPB 0.0325f
C6 A VGND 0.0158f
C7 C B 0.0893f
C8 a_392_297# VGND 3.44e-19
C9 VPWR a_465_297# 7.08e-19
C10 C a_215_297# 0.161f
C11 VPB VGND 0.0115f
C12 B X 6.65e-19
C13 a_297_297# VGND 6.5e-19
C14 a_215_297# X 0.0991f
C15 B VPWR 0.255f
C16 B a_109_53# 0.0246f
C17 A a_465_297# 5.42e-19
C18 D_N a_215_297# 3.19e-19
C19 a_215_297# VPWR 0.0871f
C20 a_215_297# a_109_53# 0.0807f
C21 a_465_297# VGND 5.02e-19
C22 C VPWR 0.00753f
C23 C a_109_53# 0.0984f
C24 B A 0.0666f
C25 X VPWR 0.0885f
C26 a_215_297# A 0.157f
C27 B VPB 0.116f
C28 B VGND 0.0161f
C29 D_N VPWR 0.0412f
C30 a_215_297# a_392_297# 0.00419f
C31 C A 0.0281f
C32 a_215_297# VPB 0.0508f
C33 a_215_297# VGND 0.237f
C34 D_N a_109_53# 0.0889f
C35 VPWR a_109_53# 0.0418f
C36 C a_392_297# 0.00267f
C37 C VPB 0.0337f
C38 C VGND 0.0202f
C39 a_215_297# a_297_297# 0.00659f
C40 A X 0.00127f
C41 C a_297_297# 0.00375f
C42 X VPB 0.011f
C43 X VGND 0.0359f
C44 A VPWR 0.0073f
C45 A a_109_53# 1.19e-19
C46 D_N VPB 0.0461f
C47 D_N VGND 0.0531f
C48 a_392_297# VPWR 5.29e-19
C49 a_215_297# a_465_297# 0.00827f
C50 VPWR VPB 0.122f
C51 VPWR VGND 0.075f
C52 VPB a_109_53# 0.0547f
C53 VGND VNB 0.469f
C54 X VNB 0.0884f
C55 A VNB 0.108f
C56 C VNB 0.101f
C57 D_N VNB 0.185f
C58 B VNB 0.101f
C59 VPWR VNB 0.399f
C60 VPB VNB 0.782f
C61 a_109_53# VNB 0.159f
C62 a_215_297# VNB 0.142f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFRTVB a_n410_n216# a_n250_n130# a_n308_n42# a_250_n42#
X0 a_250_n42# a_n250_n130# a_n308_n42# a_n410_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.5
C0 a_n308_n42# a_n250_n130# 0.0209f
C1 a_n308_n42# a_250_n42# 0.011f
C2 a_n250_n130# a_250_n42# 0.0209f
C3 a_250_n42# a_n410_n216# 0.0852f
C4 a_n308_n42# a_n410_n216# 0.0853f
C5 a_n250_n130# a_n410_n216# 1.48f
.ends

.subckt sky130_fd_pr__pfet_01v8_XQZLDL a_15_n240# w_n211_n459# a_n73_n240# a_n33_n337#
+ VSUBS
X0 a_15_n240# a_n33_n337# a_n73_n240# w_n211_n459# sky130_fd_pr__pfet_01v8 ad=0.696 pd=5.38 as=0.696 ps=5.38 w=2.4 l=0.15
C0 a_n33_n337# a_15_n240# 0.0313f
C1 a_n33_n337# w_n211_n459# 0.206f
C2 w_n211_n459# a_15_n240# 0.163f
C3 a_n33_n337# a_n73_n240# 0.0313f
C4 a_n73_n240# a_15_n240# 0.385f
C5 w_n211_n459# a_n73_n240# 0.0371f
C6 a_15_n240# VSUBS 0.11f
C7 a_n73_n240# VSUBS 0.195f
C8 a_n33_n337# VSUBS 0.139f
C9 w_n211_n459# VSUBS 1.47f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GC6 a_200_n42# w_n396_n261# a_n200_n139# a_n258_n42#
+ VSUBS
X0 a_200_n42# a_n200_n139# a_n258_n42# w_n396_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_n200_n139# a_200_n42# 0.0196f
C1 a_n200_n139# w_n396_n261# 0.73f
C2 w_n396_n261# a_200_n42# 0.0498f
C3 a_n200_n139# a_n258_n42# 0.0196f
C4 a_n258_n42# a_200_n42# 0.0134f
C5 w_n396_n261# a_n258_n42# 0.0269f
C6 a_200_n42# VSUBS 0.0338f
C7 a_n258_n42# VSUBS 0.0488f
C8 a_n200_n139# VSUBS 0.563f
C9 w_n396_n261# VSUBS 1.69f
.ends

.subckt sky130_fd_pr__nfet_01v8_ATLS57 a_15_n200# a_n73_n200# a_n33_n288# a_n141_n374#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n141_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n73_n200# a_n33_n288# 0.0312f
C1 a_n73_n200# a_15_n200# 0.321f
C2 a_n33_n288# a_15_n200# 0.0312f
C3 a_15_n200# a_n141_n374# 0.233f
C4 a_n73_n200# a_n141_n374# 0.199f
C5 a_n33_n288# a_n141_n374# 0.341f
.ends

.subckt th13 V13 Vin m1_831_275# Vn m1_559_n458# Vp
XXM0 Vn m1_559_n458# Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vn Vin m1_559_n458# m1_831_275# sky130_fd_pr__nfet_01v8_ZFRTVB
XXM2 Vp Vp m1_831_275# Vin Vn sky130_fd_pr__pfet_01v8_XQZLDL
XXM3 V13 Vp m1_831_275# Vp Vn sky130_fd_pr__pfet_01v8_VZ9GC6
XXM4 V13 Vn m1_831_275# Vn sky130_fd_pr__nfet_01v8_ATLS57
C0 Vin m1_831_275# 0.197f
C1 Vin V13 0.0076f
C2 Vin Vp 0.176f
C3 Vin m1_559_n458# 0.181f
C4 Vin Vn 0.347f
C5 m1_831_275# V13 0.184f
C6 m1_831_275# Vp 0.215f
C7 m1_831_275# m1_559_n458# 0.0183f
C8 m1_831_275# Vn 0.232f
C9 V13 Vp 0.135f
C10 m1_559_n458# Vp 0.0628f
C11 V13 Vn 0.0706f
C12 Vn Vp 0.206f
C13 m1_559_n458# Vn 0.152f
C14 m1_831_275# 0 1.05f
C15 Vin 0 1.79f
C16 V13 0 0.365f
C17 Vn 0 0.117f
C18 Vp 0 3.98f
C19 m1_559_n458# 0 0.286f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGAKDL a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
+ VSUBS
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_15_n200# w_n211_n419# 0.0336f
C1 a_15_n200# a_n33_n297# 0.0293f
C2 w_n211_n419# a_n73_n200# 0.0336f
C3 a_n73_n200# a_n33_n297# 0.0293f
C4 w_n211_n419# a_n33_n297# 0.191f
C5 a_15_n200# a_n73_n200# 0.321f
C6 a_15_n200# VSUBS 0.164f
C7 a_n73_n200# VSUBS 0.164f
C8 a_n33_n297# VSUBS 0.147f
C9 w_n211_n419# VSUBS 1.14f
.ends

.subckt sky130_fd_pr__nfet_01v8_4X3CDA a_n306_n216# a_n180_n130# a_n238_n42# a_180_n42#
X0 a_180_n42# a_n180_n130# a_n238_n42# a_n306_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.8
C0 a_n180_n130# a_180_n42# 0.0189f
C1 a_180_n42# a_n238_n42# 0.0147f
C2 a_n180_n130# a_n238_n42# 0.0189f
C3 a_180_n42# a_n306_n216# 0.075f
C4 a_n238_n42# a_n306_n216# 0.075f
C5 a_n180_n130# a_n306_n216# 1.1f
.ends

.subckt sky130_fd_pr__pfet_01v8_MWB9BZ a_15_n43# w_n211_n262# a_n73_n43# a_n33_n140#
+ VSUBS
X0 a_15_n43# a_n33_n140# a_n73_n43# w_n211_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.15
C0 a_15_n43# w_n211_n262# 0.0198f
C1 a_15_n43# a_n33_n140# 0.0193f
C2 w_n211_n262# a_n73_n43# 0.0198f
C3 a_n73_n43# a_n33_n140# 0.0193f
C4 w_n211_n262# a_n33_n140# 0.187f
C5 a_15_n43# a_n73_n43# 0.0715f
C6 a_15_n43# VSUBS 0.0453f
C7 a_n73_n43# VSUBS 0.0453f
C8 a_n33_n140# VSUBS 0.143f
C9 w_n211_n262# VSUBS 0.752f
.ends

.subckt sky130_fd_pr__pfet_01v8_JM8GTH a_50_n42# w_n246_n261# a_n50_n139# a_n108_n42#
+ VSUBS
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 a_50_n42# w_n246_n261# 0.0224f
C1 a_50_n42# a_n50_n139# 0.00909f
C2 w_n246_n261# a_n108_n42# 0.0224f
C3 a_n108_n42# a_n50_n139# 0.00909f
C4 w_n246_n261# a_n50_n139# 0.223f
C5 a_50_n42# a_n108_n42# 0.0391f
C6 a_50_n42# VSUBS 0.0488f
C7 a_n108_n42# VSUBS 0.0488f
C8 a_n50_n139# VSUBS 0.209f
C9 w_n246_n261# VSUBS 0.88f
.ends

.subckt sky130_fd_pr__nfet_01v8_L9ESAD a_n175_n190# a_n73_n50# a_n33_n138# a_15_n50#
X0 a_15_n50# a_n33_n138# a_n73_n50# a_n175_n190# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_n33_n138# a_15_n50# 0.0216f
C1 a_15_n50# a_n73_n50# 0.0826f
C2 a_n33_n138# a_n73_n50# 0.0216f
C3 a_15_n50# a_n175_n190# 0.0704f
C4 a_n73_n50# a_n175_n190# 0.0797f
C5 a_n33_n138# a_n175_n190# 0.315f
.ends

.subckt th11 V11 Vin Vp m1_705_187# Vn m1_577_n654#
XXM0 Vn Vp Vn m1_577_n654# Vn sky130_fd_pr__pfet_01v8_XGAKDL
XXM1 Vn Vin m1_577_n654# m1_705_187# sky130_fd_pr__nfet_01v8_4X3CDA
XXM2 m1_705_187# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_MWB9BZ
XXM3 V11 Vp m1_705_187# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM4 Vn Vn m1_705_187# V11 sky130_fd_pr__nfet_01v8_L9ESAD
C0 m1_577_n654# Vin 0.213f
C1 Vin V11 2.69e-19
C2 m1_705_187# Vin 0.0649f
C3 Vin Vp 0.285f
C4 m1_577_n654# V11 5.55e-19
C5 m1_577_n654# m1_705_187# 0.0258f
C6 m1_577_n654# Vp 0.0405f
C7 Vin Vn 0.135f
C8 m1_705_187# V11 0.377f
C9 m1_577_n654# Vn 0.0457f
C10 V11 Vp 0.026f
C11 m1_705_187# Vp 0.286f
C12 V11 Vn 0.00287f
C13 m1_705_187# Vn 0.463f
C14 Vp Vn 0.0775f
C15 Vin 0 1.27f
C16 m1_705_187# 0 0.602f
C17 V11 0 0.346f
C18 Vn 0 0.355f
C19 Vp 0 2.61f
C20 m1_577_n654# 0 0.286f
.ends

.subckt adc1 VGND b[0] b[1] b[2] b[3] p[0] p[10] p[11] p[12] p[13] p[14] p[1] p[2]
+ p[7] p[8] p[9] Vin
X_49_ net7 _02_ _19_ _20_ _21_ VGND VGND p[7] p[7] net17 _49_/a_208_47# _49_/a_75_199#
+ _49_/a_544_297# _49_/a_315_47# _49_/a_201_297# sky130_fd_sc_hd__a311o_1
X_48_ net11 _02_ _07_ VGND VGND p[7] p[7] _21_ _48_/a_181_47# _48_/a_109_47# _48_/a_27_47#
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_4
X_47_ net5 _12_ _17_ VGND VGND p[7] p[7] _20_ _47_/a_384_47# _47_/a_81_21# _47_/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xth02_0 th15_0/Vin p[1] th02_0/m1_983_133# p[7] th02_0/m1_571_144# VGND th02
X_46_ _04_ VGND VGND p[7] p[7] _19_ sky130_fd_sc_hd__inv_2
X_29_ net11 net13 net12 VGND VGND p[7] p[7] _03_ _29_/a_29_53# _29_/a_183_297# _29_/a_111_297#
+ sky130_fd_sc_hd__or3_1
XFILLER_0_1_43 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_6
X_28_ _00_ _01_ VGND VGND p[7] p[7] _02_ _28_/a_109_297# sky130_fd_sc_hd__nor2_1
X_45_ _02_ _09_ _12_ _13_ _18_ VGND VGND p[7] p[7] net16 _45_/a_193_297# _45_/a_465_47#
+ _45_/a_205_47# _45_/a_109_297# _45_/a_27_47# sky130_fd_sc_hd__a221o_1
X_44_ net14 _14_ _15_ _17_ net2 VGND VGND p[7] p[7] _18_ _44_/a_256_47# _44_/a_584_47#
+ _44_/a_93_21# _44_/a_250_297# _44_/a_346_47# sky130_fd_sc_hd__a32o_1
X_27_ net14 net15 net3 net2 VGND VGND p[7] p[7] _01_ _27_/a_277_297# _27_/a_205_297#
+ _27_/a_27_297# _27_/a_109_297# sky130_fd_sc_hd__or4_1
XFILLER_0_7_32 VGND p[7] p[7] VGND sky130_ef_sc_hd__decap_12
X_43_ _00_ _06_ _10_ _16_ VGND VGND p[7] p[7] _17_ _43_/a_369_47# _43_/a_469_47# _43_/a_297_47#
+ _43_/a_193_413# _43_/a_27_47# sky130_fd_sc_hd__and4b_1
X_26_ net5 net4 net6 VGND VGND p[7] p[7] _00_ _26_/a_29_53# _26_/a_183_297# _26_/a_111_297#
+ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
XFILLER_0_7_44 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_4
X_42_ net3 net15 net14 VGND VGND p[7] p[7] _16_ _42_/a_109_93# _42_/a_368_53# _42_/a_209_311#
+ _42_/a_296_53# sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_3_Left_11 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND p[7] p[7] b[0] output16/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_41_ _06_ _10_ VGND VGND p[7] p[7] _15_ _41_/a_145_75# _41_/a_59_75# sky130_fd_sc_hd__and2_1
Xoutput17 net17 VGND VGND p[7] p[7] b[1] output17/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_40_ net15 net3 net2 _00_ VGND VGND p[7] p[7] _14_ _40_/a_297_297# _40_/a_191_297#
+ _40_/a_109_297# sky130_fd_sc_hd__nor4_1
Xoutput18 net18 VGND VGND p[7] p[7] b[2] output18/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
Xth09_0 p[8] Vin VGND th09_0/m1_485_n505# p[7] th09_0/m1_962_372# th09
XPHY_EDGE_ROW_0_Left_8 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_15 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND p[7] p[7] b[3] output19/a_27_47# sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_15 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_6
Xth14_0 p[13] th15_0/Vin VGND th14_0/m1_641_n318# p[7] th14_0/m1_891_419# th14
Xinput1 p[0] VGND VGND p[7] p[7] net1 input1/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput2 p[10] VGND VGND p[7] p[7] net2 input2/a_27_47# sky130_fd_sc_hd__buf_1
Xinput3 p[11] VGND VGND p[7] p[7] net3 input3/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
Xth12_0 p[11] Vin th12_0/m1_394_n856# th12_0/m1_529_n42# p[7] VGND th12
Xinput4 p[12] VGND VGND p[7] p[7] net4 input4/a_75_212# sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_10 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
XFILLER_0_2_42 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_6
Xinput5 p[13] VGND VGND p[7] p[7] net5 input5/a_664_47# input5/a_841_47# input5/a_381_47#
+ input5/a_62_47# input5/a_558_47# sky130_fd_sc_hd__dlymetal6s2s_1
Xinput6 p[14] VGND VGND p[7] p[7] net6 input6/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_1_Left_9 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Right_4 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
Xth10_0 p[9] Vin th10_0/m1_502_n495# th10_0/m1_536_174# VGND p[7] th10
Xinput7 p[1] VGND VGND p[7] p[7] net7 input7/a_27_47# sky130_fd_sc_hd__buf_1
Xinput10 p[7] VGND VGND p[7] p[7] net10 input10/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_14 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
Xth03_0 p[2] Vin p[7] th03_0/m1_890_n844# th03_0/m1_638_n591# VGND th03
XFILLER_0_5_45 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_4
Xinput8 p[2] VGND VGND p[7] p[7] net8 input8/a_27_47# sky130_fd_sc_hd__buf_1
Xinput11 p[7] VGND VGND p[7] p[7] net11 input11/a_27_47# sky130_fd_sc_hd__buf_1
X_39_ net5 net6 VGND VGND p[7] p[7] _13_ _39_/a_129_47# _39_/a_47_47# _39_/a_285_47#
+ _39_/a_377_297# sky130_fd_sc_hd__xnor2_1
Xinput9 p[7] VGND VGND p[7] p[7] net9 input9/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput12 p[7] VGND VGND p[7] p[7] net12 input12/a_27_47# sky130_fd_sc_hd__buf_1
X_55_ _14_ _15_ _20_ _22_ VGND VGND p[7] p[7] net19 _55_/a_472_297# _55_/a_80_21#
+ _55_/a_300_47# _55_/a_217_297# sky130_fd_sc_hd__a211o_1
X_38_ net4 _06_ _10_ _11_ VGND VGND p[7] p[7] _12_ _38_/a_109_47# _38_/a_197_47# _38_/a_303_47#
+ _38_/a_27_47# sky130_fd_sc_hd__and4_1
X_54_ _25_ VGND VGND p[7] p[7] net18 _54_/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput13 p[7] VGND VGND p[7] p[7] net13 input13/a_27_47# sky130_fd_sc_hd__buf_1
X_37_ net14 net15 net3 net2 VGND VGND p[7] p[7] _11_ _37_/a_109_47# _37_/a_197_47#
+ _37_/a_303_47# _37_/a_27_47# sky130_fd_sc_hd__and4_1
Xth01_0 p[0] VGND th01_0/m1_991_n1219# th01_0/m1_571_n501# p[7] th15_0/Vin th01
Xinput14 p[8] VGND VGND p[7] p[7] net14 input14/a_27_47# sky130_fd_sc_hd__buf_1
X_53_ _21_ _22_ _24_ VGND VGND p[7] p[7] _25_ _53_/a_29_53# _53_/a_183_297# _53_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_36_ net11 net10 net13 net12 VGND VGND p[7] p[7] _10_ _36_/a_109_47# _36_/a_197_47#
+ _36_/a_303_47# _36_/a_27_47# sky130_fd_sc_hd__and4_1
X_52_ _02_ _06_ _23_ _12_ net5 VGND VGND p[7] p[7] _24_ _52_/a_256_47# _52_/a_584_47#
+ _52_/a_93_21# _52_/a_250_297# _52_/a_346_47# sky130_fd_sc_hd__a32o_1
Xinput15 p[9] VGND VGND p[7] p[7] net15 input15/a_27_47# sky130_fd_sc_hd__buf_1
X_35_ _04_ _05_ _07_ _08_ VGND VGND p[7] p[7] _09_ _35_/a_489_413# _35_/a_226_47#
+ _35_/a_556_47# _35_/a_226_297# _35_/a_76_199# sky130_fd_sc_hd__a2bb2o_1
X_51_ _03_ VGND VGND p[7] p[7] _23_ sky130_fd_sc_hd__inv_2
X_34_ net11 net12 VGND VGND p[7] p[7] _08_ _34_/a_129_47# _34_/a_47_47# _34_/a_285_47#
+ _34_/a_377_297# sky130_fd_sc_hd__xnor2_1
X_33_ net13 _06_ net10 VGND VGND p[7] p[7] _07_ _33_/a_109_93# _33_/a_368_53# _33_/a_209_311#
+ _33_/a_296_53# sky130_fd_sc_hd__and3b_1
X_50_ net5 net6 _15_ _11_ VGND VGND p[7] p[7] _22_ _50_/a_515_93# _50_/a_223_47# _50_/a_615_93#
+ _50_/a_343_93# _50_/a_429_93# _50_/a_27_47# sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
Xpreamp_0 Vin th15_0/Vin VGND p[7] preamp
X_32_ net7 net1 net9 net8 VGND VGND p[7] p[7] _06_ _32_/a_109_47# _32_/a_197_47# _32_/a_303_47#
+ _32_/a_27_47# sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_5_Left_13 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
XFILLER_0_0_20 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_4
X_31_ net7 net8 VGND VGND p[7] p[7] _05_ _31_/a_117_297# _31_/a_285_297# _31_/a_285_47#
+ _31_/a_35_297# sky130_fd_sc_hd__xor2_1
Xth15_0 p[14] th15_0/Vin th15_0/m1_597_n912# th15_0/m1_849_n157# p[7] VGND th15
X_30_ net9 net10 _03_ net1 VGND VGND p[7] p[7] _04_ _30_/a_465_297# _30_/a_297_297#
+ _30_/a_215_297# _30_/a_392_297# _30_/a_109_53# sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
XFILLER_0_0_34 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_4
XFILLER_0_3_45 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_4
XFILLER_0_0_13 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_4
Xth13_0 p[12] Vin th13_0/m1_831_275# VGND th13_0/m1_559_n458# p[7] th13
XFILLER_0_3_13 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_4
XFILLER_0_6_25 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
XFILLER_0_6_36 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_6
XFILLER_0_3_37 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_4
Xth11_0 p[10] Vin p[7] th11_0/m1_705_187# VGND th11_0/m1_577_n654# th11
XPHY_EDGE_ROW_2_Right_2 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_12 VGND VGND p[7] p[7] sky130_fd_sc_hd__decap_3
C0 _27_/a_277_297# net15 1.93e-19
C1 _04_ _33_/a_109_93# 0.0299f
C2 _34_/a_47_47# _25_ 1.08e-19
C3 _10_ _30_/a_297_297# 1.25e-20
C4 _08_ _21_ 0.00139f
C5 p[7] _50_/a_615_93# -5.34e-19
C6 VGND th02_0/m1_571_144# 0.00939f
C7 p[2] th03_0/m1_890_n844# 0.0404f
C8 _27_/a_27_297# _01_ 8.04e-19
C9 _29_/a_183_297# _03_ 7.36e-19
C10 input9/a_75_212# net13 4.4e-19
C11 net10 _31_/a_285_297# 1.68e-19
C12 VGND _18_ 0.0166f
C13 _12_ _50_/a_27_47# 0.00354f
C14 VGND _26_/a_111_297# -2.75e-19
C15 _01_ _31_/a_285_47# 3.36e-19
C16 _08_ _35_/a_226_47# 0.00117f
C17 net3 p[10] 3.61e-19
C18 net4 _50_/a_429_93# 4.16e-19
C19 net6 _50_/a_343_93# 0.00214f
C20 Vin p[10] 0.0929f
C21 th14_0/m1_891_419# input5/a_558_47# 3.96e-20
C22 _44_/a_250_297# _16_ 3.25e-19
C23 net2 net10 2.05e-20
C24 _10_ _50_/a_223_47# 0.0295f
C25 _06_ _41_/a_59_75# 0.0457f
C26 _13_ _50_/a_343_93# 5.63e-20
C27 _52_/a_346_47# _06_ 0.0031f
C28 input8/a_27_47# input7/a_27_47# 3.2e-20
C29 VGND _26_/a_29_53# 0.0381f
C30 _17_ _37_/a_109_47# 8.86e-21
C31 p[7] _42_/a_296_53# -6.37e-20
C32 p[7] _16_ 0.126f
C33 _04_ _27_/a_27_297# 0.0526f
C34 _44_/a_584_47# net14 7.2e-19
C35 net11 _12_ 0.00799f
C36 VGND b[3] 0.148f
C37 net12 input13/a_27_47# 0.0163f
C38 _09_ _23_ 0.207f
C39 input5/a_841_47# net15 0.00585f
C40 net9 _30_/a_297_297# 7.53e-19
C41 p[7] th03_0/m1_890_n844# 0.0198f
C42 _47_/a_81_21# _18_ 7.96e-20
C43 _47_/a_384_47# _17_ 1.1e-20
C44 _07_ _24_ 5.67e-19
C45 _06_ _22_ 0.124f
C46 _11_ _39_/a_377_297# 2.57e-20
C47 p[0] net1 0.00473f
C48 p[7] _48_/a_27_47# 0.0162f
C49 _06_ _11_ 0.493f
C50 _06_ net7 0.00447f
C51 p[7] _31_/a_117_297# 5.04e-19
C52 net2 _44_/a_93_21# 0.0273f
C53 _22_ output18/a_27_47# 7.51e-19
C54 _02_ _39_/a_47_47# 0.0127f
C55 _44_/a_256_47# _44_/a_93_21# -6.6e-20
C56 net2 th11_0/m1_705_187# 1.39e-19
C57 net9 _50_/a_223_47# 2e-19
C58 _45_/a_27_47# _50_/a_27_47# 0.109f
C59 p[11] p[13] 0.0167f
C60 net7 p[2] 0.00157f
C61 _02_ net10 6.74e-19
C62 net6 net5 0.727f
C63 _41_/a_59_75# p[7] 0.0186f
C64 _13_ net5 0.0381f
C65 p[7] input2/a_27_47# 0.00832f
C66 _52_/a_346_47# p[7] -0.00109f
C67 net17 input5/a_558_47# 2.88e-21
C68 _42_/a_368_53# net3 3.82e-19
C69 p[2] _49_/a_208_47# 4.19e-20
C70 _41_/a_59_75# th15_0/m1_849_n157# 0.00112f
C71 th15_0/Vin _40_/a_297_297# 1.26e-19
C72 input5/a_664_47# _19_ 2.19e-21
C73 _45_/a_27_47# net11 3.64e-20
C74 input3/a_27_47# net3 0.03f
C75 _06_ net12 0.284f
C76 net14 _21_ 7.17e-21
C77 net1 _27_/a_27_297# 6.05e-21
C78 _52_/a_93_21# net6 2.33e-19
C79 _52_/a_250_297# net4 0.00136f
C80 _54_/a_75_212# _38_/a_27_47# 2.67e-19
C81 _52_/a_93_21# _13_ 1.31e-19
C82 input5/a_664_47# net5 0.0536f
C83 _03_ _27_/a_277_297# 2.1e-20
C84 VGND _33_/a_209_311# -0.00749f
C85 _30_/a_109_53# net10 5.6e-20
C86 th15_0/Vin input7/a_27_47# 2.79e-19
C87 _22_ p[7] 1.4f
C88 net11 _36_/a_303_47# 7.63e-20
C89 p[7] _11_ 0.352f
C90 net7 p[7] 0.786f
C91 _44_/a_584_47# b[3] 1.27e-19
C92 _38_/a_27_47# net16 0.114f
C93 net2 net15 0.324f
C94 p[13] net8 0.00375f
C95 _14_ p[14] 1.13e-19
C96 _23_ _39_/a_47_47# 5.24e-21
C97 _35_/a_76_199# _01_ 3.08e-21
C98 _11_ th15_0/m1_849_n157# 7.84e-20
C99 VGND _47_/a_81_21# -0.0112f
C100 net4 _24_ 8.65e-20
C101 net6 _15_ 0.17f
C102 _10_ _12_ 0.19f
C103 VGND th10_0/m1_502_n495# 0.0046f
C104 net4 _14_ 1.54e-20
C105 _15_ _13_ 3.69e-20
C106 p[7] _49_/a_208_47# -5.93e-19
C107 _38_/a_27_47# _21_ 3.87e-19
C108 _23_ net10 0.00216f
C109 _49_/a_544_297# net13 3.43e-19
C110 Vin th02_0/m1_983_133# 0.0615f
C111 input5/a_664_47# b[1] 0.00195f
C112 _18_ net16 8.17e-21
C113 p[9] net14 1.05e-19
C114 _04_ _35_/a_76_199# 0.0269f
C115 _42_/a_209_311# th14_0/m1_641_n318# 1.87e-19
C116 _19_ _42_/a_109_93# 1.14e-21
C117 net19 net14 0.148f
C118 p[0] p[10] 0.00247f
C119 VGND output17/a_27_47# 0.00246f
C120 p[7] th15_0/m1_597_n912# 2.46e-19
C121 _07_ _20_ 1.28e-21
C122 _15_ input5/a_664_47# 9.15e-22
C123 net12 p[7] 0.9f
C124 _42_/a_109_93# net5 0.00109f
C125 input7/a_27_47# input5/a_558_47# 1.22e-20
C126 _34_/a_285_47# _06_ 0.00598f
C127 _34_/a_377_297# _07_ 5.8e-19
C128 th15_0/m1_849_n157# th15_0/m1_597_n912# -5.55e-35
C129 _17_ _00_ 0.0851f
C130 VGND _44_/a_584_47# -0.00145f
C131 _45_/a_465_47# p[7] -5.05e-19
C132 _08_ _04_ 5.99e-19
C133 _02_ net15 0.0806f
C134 net9 _12_ 4.39e-22
C135 _15_ _50_/a_429_93# 6.82e-19
C136 _14_ _50_/a_343_93# 9.76e-19
C137 net4 _45_/a_193_297# 7.41e-19
C138 _12_ _53_/a_29_53# 3.46e-20
C139 net6 _45_/a_109_297# 7.82e-19
C140 _42_/a_109_93# b[1] 2.38e-19
C141 _10_ _45_/a_27_47# 0.0143f
C142 _06_ _48_/a_109_47# 9.47e-19
C143 _43_/a_297_47# _00_ 1.26e-19
C144 p[1] _19_ 3.92e-20
C145 VGND th13_0/m1_559_n458# 0.0449f
C146 _27_/a_27_297# p[10] 1.63e-19
C147 _10_ _36_/a_303_47# 4.09e-19
C148 input15/a_27_47# net15 0.00325f
C149 _18_ net19 4.89e-20
C150 _15_ _42_/a_109_93# 0.00367f
C151 VGND _54_/a_75_212# 0.053f
C152 _10_ input6/a_27_47# 4.57e-20
C153 _52_/a_250_297# net5 0.018f
C154 _31_/a_285_47# p[10] 2.16e-20
C155 _06_ input5/a_381_47# 1.6e-19
C156 _03_ _31_/a_285_297# 0.00677f
C157 net17 _31_/a_117_297# 0.00149f
C158 p[12] _39_/a_129_47# 2.4e-20
C159 _38_/a_27_47# output16/a_27_47# 9.02e-19
C160 VGND net16 0.144f
C161 _07_ _29_/a_29_53# 1.19e-20
C162 _32_/a_27_47# _43_/a_27_47# 2.01e-20
C163 p[9] b[3] 0.134f
C164 _34_/a_285_47# p[7] -0.00191f
C165 _39_/a_47_47# net3 1.66e-20
C166 _14_ _19_ 2.71e-21
C167 _12_ _05_ 2.52e-19
C168 _07_ net11 0.0206f
C169 net2 _03_ 1.89e-19
C170 net7 _49_/a_315_47# 0.00706f
C171 net19 b[3] 0.0546f
C172 VGND _21_ 0.295f
C173 net4 _20_ 3.01e-20
C174 _52_/a_93_21# _52_/a_250_297# -6.97e-22
C175 _24_ net5 5.83e-20
C176 _14_ net5 3.89e-19
C177 input2/a_27_47# net17 0.0398f
C178 p[1] b[1] 0.00395f
C179 VGND input11/a_27_47# 0.0274f
C180 p[7] _48_/a_109_47# 3.35e-21
C181 net14 _01_ 8.29e-19
C182 VGND _35_/a_226_47# -0.0111f
C183 _36_/a_109_47# net13 0.00126f
C184 p[7] th12_0/m1_529_n42# 0.0444f
C185 _52_/a_93_21# _24_ 0.0211f
C186 _24_ b[1] 2.68e-19
C187 _14_ b[1] 1.1e-19
C188 p[0] th02_0/m1_983_133# 0.0563f
C189 net9 p[13] 1.72e-19
C190 _35_/a_226_47# _33_/a_209_311# 1.31e-19
C191 VGND p[9] 0.443f
C192 _04_ net14 0.0863f
C193 net7 net17 0.2f
C194 input5/a_381_47# p[7] 8.33e-19
C195 _12_ input4/a_75_212# 2.09e-20
C196 p[7] _29_/a_183_297# -8.13e-19
C197 _44_/a_93_21# net3 0.0102f
C198 Vin _44_/a_93_21# 2.93e-21
C199 _20_ _50_/a_343_93# 0.00826f
C200 _06_ _17_ 0.0341f
C201 VGND net19 0.151f
C202 net4 _50_/a_27_47# 0.0239f
C203 _02_ _03_ 0.00474f
C204 _45_/a_27_47# _05_ 9.34e-23
C205 net13 _30_/a_297_297# 3.27e-20
C206 _15_ _14_ 0.148f
C207 _52_/a_93_21# net18 8.21e-21
C208 th11_0/m1_705_187# Vin 0.0585f
C209 input12/a_27_47# b[1] 0.00658f
C210 net18 b[1] 0.00134f
C211 _06_ _40_/a_109_297# 0.00175f
C212 _45_/a_193_297# net5 0.00935f
C213 _09_ _33_/a_109_93# 7.36e-20
C214 net12 _29_/a_111_297# 1.21e-19
C215 _18_ _01_ 6.1e-20
C216 _55_/a_300_47# _02_ 0.00371f
C217 input2/a_27_47# input7/a_27_47# 1.62e-19
C218 th10_0/m1_502_n495# p[9] 0.0156f
C219 _03_ _30_/a_109_53# 0.0189f
C220 p[13] _49_/a_201_297# 6.25e-20
C221 b[0] _39_/a_47_47# 2.04e-19
C222 net12 net17 2.11e-21
C223 _10_ _39_/a_285_47# 0.00289f
C224 _17_ output19/a_27_47# 0.00122f
C225 _06_ _43_/a_297_47# 4.81e-20
C226 net2 _00_ 0.00732f
C227 VGND output16/a_27_47# 0.0728f
C228 _52_/a_93_21# _45_/a_193_297# 6.01e-19
C229 _32_/a_303_47# net5 7.18e-21
C230 th03_0/m1_638_n591# th15_0/Vin 2.04e-19
C231 _10_ _07_ 2.19e-19
C232 _40_/a_297_297# _11_ 9.94e-19
C233 _04_ _18_ 1.94e-21
C234 th13_0/m1_559_n458# net16 6.79e-20
C235 _20_ _19_ 0.00734f
C236 _50_/a_27_47# _50_/a_343_93# -7.11e-33
C237 _17_ _44_/a_250_297# 0.0336f
C238 net3 net15 0.394f
C239 Vin net15 0.0041f
C240 _45_/a_27_47# input4/a_75_212# 2.18e-20
C241 _54_/a_75_212# net16 1.69e-21
C242 _25_ net18 0.0594f
C243 _22_ _53_/a_183_297# 3.71e-20
C244 _23_ _03_ 0.0564f
C245 _04_ _26_/a_29_53# 2.3e-21
C246 p[11] th09_0/m1_485_n505# 1.22e-20
C247 _45_/a_205_47# _12_ 7.46e-19
C248 _20_ net5 0.0651f
C249 p[7] _17_ 0.306f
C250 _50_/a_343_93# net8 7.25e-19
C251 VGND _32_/a_109_47# 1.05e-19
C252 net1 net14 6.64e-20
C253 net7 input7/a_27_47# 0.00318f
C254 th14_0/m1_891_419# th12_0/m1_529_n42# 0.00211f
C255 p[13] input5/a_62_47# 0.0281f
C256 _17_ th15_0/m1_849_n157# 8.52e-20
C257 p[7] _40_/a_109_297# -4.23e-19
C258 _06_ input5/a_841_47# 1.66e-19
C259 net16 _21_ 1.89e-19
C260 p[11] input14/a_27_47# 3.98e-20
C261 input5/a_381_47# th14_0/m1_891_419# 4.77e-20
C262 _14_ _49_/a_75_199# 6.79e-20
C263 p[8] net14 0.01f
C264 _07_ net9 1.39e-20
C265 _20_ b[1] 0.00465f
C266 _43_/a_297_47# p[7] -2.11e-19
C267 _02_ _00_ 0.0269f
C268 _02_ _36_/a_27_47# 9.37e-20
C269 p[7] _27_/a_277_297# -3.63e-19
C270 _34_/a_377_297# b[1] 0.00115f
C271 VGND _01_ 0.0939f
C272 th12_0/m1_394_n856# th14_0/m1_641_n318# 1.54e-19
C273 _10_ p[14] 0.00247f
C274 _15_ _20_ 0.691f
C275 _19_ net8 0.0322f
C276 p[11] b[1] 2.45e-20
C277 _33_/a_109_93# net10 0.0336f
C278 _50_/a_27_47# net5 0.0169f
C279 _34_/a_47_47# _24_ 6.84e-21
C280 _35_/a_226_47# _21_ 9.87e-19
C281 _10_ net4 0.183f
C282 net6 _13_ 0.0106f
C283 _37_/a_27_47# net14 0.0584f
C284 _40_/a_191_297# net15 8.41e-19
C285 _37_/a_109_47# net3 0.00212f
C286 _30_/a_109_53# _00_ 3.67e-20
C287 net11 _19_ 6.27e-21
C288 net4 _55_/a_80_21# 1.06e-19
C289 net8 net5 0.48f
C290 VGND _04_ 0.135f
C291 _29_/a_29_53# net5 8.1e-20
C292 th15_0/Vin input1/a_75_212# 0.00156f
C293 _15_ p[11] 0.00591f
C294 th15_0/Vin th11_0/m1_577_n654# 0.00967f
C295 th13_0/m1_831_275# p[14] 4.94e-20
C296 VGND _38_/a_109_47# 2.3e-19
C297 net11 net5 0.0129f
C298 _12_ net13 0.00632f
C299 th15_0/Vin _37_/a_303_47# 1.45e-19
C300 _07_ _05_ 1.21e-19
C301 p[0] th11_0/m1_705_187# 1.49e-19
C302 _47_/a_81_21# _01_ 6.05e-21
C303 _34_/a_47_47# input12/a_27_47# 2.17e-19
C304 th15_0/Vin th14_0/m1_641_n318# 7.77e-19
C305 net4 th13_0/m1_831_275# 3.27e-19
C306 p[7] input5/a_841_47# 0.0775f
C307 _04_ _33_/a_209_311# 0.00133f
C308 _06_ _31_/a_285_297# 1.01e-20
C309 th13_0/m1_559_n458# output16/a_27_47# 1.24e-20
C310 _23_ _36_/a_27_47# 0.00118f
C311 input5/a_381_47# net17 1.37e-20
C312 th01_0/m1_991_n1219# th15_0/Vin -8.41e-19
C313 VGND _53_/a_111_297# -2.89e-19
C314 net8 b[1] 0.0729f
C315 net7 _49_/a_544_297# 2.72e-19
C316 _06_ net2 0.0108f
C317 _29_/a_29_53# b[1] 0.0026f
C318 _52_/a_93_21# net11 2.8e-19
C319 _15_ _50_/a_27_47# 5.65e-19
C320 VGND _26_/a_183_297# 2.42e-19
C321 net14 p[10] 1.59e-20
C322 _09_ _35_/a_76_199# 0.047f
C323 _08_ _35_/a_489_413# 5.56e-19
C324 net11 b[1] 0.0777f
C325 p[2] _31_/a_285_297# 0.00165f
C326 net16 output16/a_27_47# 0.0101f
C327 net6 _50_/a_429_93# 6.18e-19
C328 _03_ net3 4.27e-20
C329 net9 net4 1.99e-22
C330 _10_ _50_/a_343_93# 0.0284f
C331 p[8] b[3] 0.0392f
C332 _52_/a_584_47# _06_ 0.00218f
C333 _15_ net8 1.79e-19
C334 _17_ _37_/a_197_47# 9.19e-21
C335 _18_ _37_/a_27_47# 3.31e-20
C336 _12_ p[12] 0.00589f
C337 net4 _53_/a_29_53# 3.26e-19
C338 _42_/a_209_311# p[14] 5.85e-22
C339 net19 p[9] 0.0767f
C340 net2 output19/a_27_47# 0.00168f
C341 _08_ _09_ 0.106f
C342 _49_/a_75_199# _20_ 0.0233f
C343 _04_ output17/a_27_47# 0.027f
C344 VGND net1 0.513f
C345 th15_0/Vin _12_ 0.00101f
C346 p[7] _31_/a_285_297# 0.013f
C347 net2 _44_/a_250_297# 0.0188f
C348 net13 _36_/a_303_47# 5.5e-20
C349 _25_ net11 0.0262f
C350 _44_/a_346_47# _44_/a_93_21# -5.12e-20
C351 _19_ _27_/a_109_297# 7.54e-21
C352 net9 _50_/a_343_93# 6.64e-19
C353 _06_ _02_ 0.85f
C354 p[7] net2 0.958f
C355 _30_/a_215_297# net5 8.27e-21
C356 p[7] th09_0/m1_962_372# 0.00391f
C357 p[7] _44_/a_256_47# -7.56e-19
C358 VGND p[8] 0.129f
C359 _22_ b[2] 0.0043f
C360 _10_ net5 0.199f
C361 _52_/a_584_47# p[7] -9.47e-19
C362 _02_ output18/a_27_47# 4.13e-19
C363 _55_/a_80_21# net5 2.78e-19
C364 th14_0/m1_891_419# input5/a_841_47# 3.61e-21
C365 net1 _47_/a_81_21# 1.58e-21
C366 _45_/a_27_47# p[12] 2.9e-19
C367 _30_/a_465_297# b[1] 4.8e-19
C368 _42_/a_368_53# net14 7.39e-19
C369 p[2] _02_ 8.49e-19
C370 _27_/a_27_297# net15 0.00888f
C371 _45_/a_109_297# net11 7.46e-20
C372 input3/a_27_47# net14 3.47e-19
C373 _06_ _30_/a_109_53# 1.96e-19
C374 _06_ input15/a_27_47# 4.73e-19
C375 _30_/a_215_297# b[1] 0.0176f
C376 _01_ _21_ 7.94e-19
C377 _52_/a_250_297# net6 0.00133f
C378 _10_ _52_/a_93_21# 0.00534f
C379 _52_/a_250_297# _13_ 5.43e-19
C380 VGND _37_/a_27_47# -0.0147f
C381 _49_/a_75_199# net8 0.00214f
C382 VGND _33_/a_296_53# -1.43e-19
C383 b[1] _27_/a_109_297# 8.35e-20
C384 _49_/a_75_199# _29_/a_29_53# 1.28e-19
C385 net3 _00_ 2.12e-19
C386 _35_/a_76_199# net10 0.0226f
C387 _10_ b[1] 2.37e-20
C388 th10_0/m1_502_n495# p[8] 1.22e-20
C389 _55_/a_80_21# b[1] 6.03e-19
C390 _38_/a_109_47# net16 4.17e-19
C391 net1 output17/a_27_47# 8.12e-19
C392 _49_/a_75_199# net11 4.49e-19
C393 net4 input4/a_75_212# 0.0178f
C394 _06_ _23_ 0.218f
C395 _43_/a_193_413# _12_ 7.94e-22
C396 VGND _47_/a_299_297# -3.63e-19
C397 _04_ _21_ 0.39f
C398 net6 _24_ 0.00121f
C399 p[7] _02_ 0.332f
C400 net9 net5 0.0368f
C401 th03_0/m1_638_n591# net7 3.67e-20
C402 input5/a_664_47# p[1] 1.21e-20
C403 net6 _14_ 2.11e-19
C404 _24_ _13_ 2.47e-19
C405 _14_ _13_ 1.47e-20
C406 _10_ _15_ 0.479f
C407 _15_ _55_/a_80_21# 0.107f
C408 th15_0/Vin input6/a_27_47# 0.00615f
C409 _08_ net10 0.194f
C410 _32_/a_27_47# _18_ 1.18e-20
C411 _04_ _35_/a_226_47# 0.00551f
C412 _32_/a_197_47# _02_ 3.78e-19
C413 _42_/a_296_53# th14_0/m1_641_n318# 8.45e-21
C414 th14_0/m1_641_n318# _16_ 2.77e-20
C415 th15_0/Vin p[13] 0.0887f
C416 p[7] _28_/a_109_297# -1.71e-19
C417 _34_/a_47_47# net11 0.0309f
C418 net19 _01_ 4.9e-19
C419 VGND p[10] 0.388f
C420 _53_/a_111_297# _21_ 4.38e-19
C421 p[7] _30_/a_109_53# 0.00151f
C422 _10_ _25_ 0.0109f
C423 p[7] input15/a_27_47# 0.0113f
C424 _42_/a_209_311# net5 3.27e-21
C425 net9 b[1] 0.0765f
C426 th14_0/m1_891_419# net2 0.011f
C427 _52_/a_93_21# _53_/a_29_53# 0.00116f
C428 _53_/a_29_53# b[1] 4.99e-19
C429 _33_/a_109_93# _03_ 2.78e-19
C430 VGND _55_/a_472_297# -0.00188f
C431 _19_ _31_/a_35_297# 1.47e-19
C432 _04_ net19 2.07e-20
C433 _22_ _50_/a_223_47# 0.031f
C434 net9 _15_ 0.00113f
C435 _15_ _50_/a_515_93# 0.00147f
C436 _09_ _38_/a_27_47# 0.00195f
C437 input3/a_27_47# b[3] 1.4e-19
C438 p[7] th10_0/m1_536_174# 0.0406f
C439 _07_ net13 0.00686f
C440 _50_/a_223_47# _11_ 0.0329f
C441 net2 _37_/a_197_47# 4.74e-20
C442 p[7] _23_ -0.00374f
C443 net6 _45_/a_193_297# 9.84e-20
C444 _31_/a_35_297# net5 2.04e-21
C445 _42_/a_209_311# b[1] 5.21e-19
C446 _10_ _45_/a_109_297# 0.00202f
C447 net1 _21_ 0.0252f
C448 p[13] input5/a_558_47# 0.00363f
C449 _19_ input5/a_62_47# 0.00159f
C450 _09_ _18_ 7.01e-21
C451 _52_/a_93_21# _05_ 1.12e-20
C452 net12 _30_/a_297_297# 7.14e-21
C453 _27_/a_27_297# _03_ 2.68e-19
C454 th01_0/m1_571_n501# Vin 0.00112f
C455 _49_/a_201_297# b[1] 0.0025f
C456 _15_ _42_/a_209_311# 0.0521f
C457 _14_ _42_/a_109_93# 0.00141f
C458 _05_ b[1] 0.0316f
C459 _32_/a_109_47# _01_ 0.00129f
C460 input5/a_62_47# net5 0.00329f
C461 _25_ _53_/a_29_53# 0.00146f
C462 net1 _35_/a_226_47# 1.3e-20
C463 _03_ _31_/a_285_47# 8.54e-19
C464 b[1] _31_/a_35_297# 0.0176f
C465 output17/a_27_47# p[10] 0.12f
C466 p[12] _39_/a_285_47# 3.03e-19
C467 net7 input1/a_75_212# 3.77e-19
C468 VGND _32_/a_27_47# 0.0233f
C469 VGND _42_/a_368_53# -4.05e-19
C470 net2 net17 0.261f
C471 VGND input3/a_27_47# 0.0414f
C472 _06_ net3 0.0072f
C473 input4/a_75_212# net5 0.0104f
C474 _06_ Vin 7.82e-20
C475 net6 _20_ 9.69e-20
C476 _20_ _13_ 7.38e-21
C477 _52_/a_93_21# _52_/a_256_47# -6.6e-20
C478 _49_/a_315_47# _02_ 0.00134f
C479 input5/a_62_47# b[1] 0.0024f
C480 _52_/a_256_47# b[1] 8.49e-20
C481 _43_/a_27_47# _00_ 0.0431f
C482 p[2] Vin 0.0232f
C483 VGND _35_/a_489_413# -8.78e-19
C484 _32_/a_27_47# _47_/a_81_21# 5.06e-21
C485 p[9] p[8] 0.11f
C486 _41_/a_59_75# _12_ 0.00101f
C487 net9 _49_/a_75_199# 0.00382f
C488 _52_/a_250_297# _24_ 3.03e-19
C489 _52_/a_346_47# _12_ 3.8e-19
C490 net4 net13 2.48e-19
C491 net3 output19/a_27_47# 0.00356f
C492 Vin output19/a_27_47# 0.00177f
C493 VGND th02_0/m1_983_133# 0.0724f
C494 net19 p[8] 0.00885f
C495 _35_/a_489_413# _33_/a_209_311# 2.77e-20
C496 _04_ _01_ 0.119f
C497 input10/a_27_47# b[1] 0.00691f
C498 _18_ _39_/a_47_47# 1.23e-19
C499 _17_ _39_/a_129_47# 1.38e-20
C500 VGND _09_ 0.397f
C501 _44_/a_93_21# net14 0.0646f
C502 _44_/a_250_297# net3 0.0088f
C503 _40_/a_297_297# net2 0.00101f
C504 net6 _50_/a_27_47# 0.0428f
C505 _22_ _12_ 0.196f
C506 _45_/a_109_297# _05_ 2.79e-22
C507 _13_ _50_/a_27_47# 0.00169f
C508 _02_ net17 0.0608f
C509 _12_ _11_ 0.195f
C510 p[7] net3 0.351f
C511 p[7] Vin 2.2f
C512 _34_/a_47_47# net9 1.41e-20
C513 p[12] p[14] 2.26e-19
C514 p[9] _37_/a_27_47# 0.0117f
C515 _18_ net10 1.47e-21
C516 _06_ _40_/a_191_297# 5.84e-19
C517 input3/a_27_47# output17/a_27_47# 3.15e-19
C518 _45_/a_205_47# net5 8.28e-20
C519 net6 _29_/a_29_53# 1.4e-20
C520 _08_ _33_/a_368_53# 5.04e-19
C521 _09_ _33_/a_209_311# 3.79e-20
C522 net2 input7/a_27_47# 3.24e-19
C523 Vin th15_0/m1_849_n157# 0.0502f
C524 net4 p[12] 0.0242f
C525 _34_/a_47_47# _53_/a_29_53# 5.88e-22
C526 net19 _37_/a_27_47# 0.0105f
C527 net6 net11 1.08e-19
C528 net11 _13_ 2.34e-19
C529 net18 _24_ 5.57e-21
C530 _26_/a_29_53# net10 3.48e-22
C531 _30_/a_109_53# net17 4.18e-20
C532 _49_/a_75_199# _31_/a_35_297# 6.24e-19
C533 th15_0/Vin p[14] 0.356f
C534 _25_ input10/a_27_47# 2.03e-20
C535 _06_ _43_/a_369_47# -2.02e-19
C536 _35_/a_76_199# _03_ 0.0733f
C537 input5/a_664_47# net8 0.0116f
C538 input13/a_27_47# _33_/a_109_93# 0.00348f
C539 net4 th15_0/Vin 3.6e-19
C540 p[11] _42_/a_109_93# 3.74e-19
C541 net12 _12_ 7.94e-21
C542 p[0] th01_0/m1_571_n501# 2.36e-19
C543 output17/a_27_47# th02_0/m1_983_133# 0.00138f
C544 _18_ _44_/a_93_21# 0.00485f
C545 net14 net15 1.07f
C546 _45_/a_465_47# _12_ 0.00211f
C547 _34_/a_47_47# _05_ 1.26e-20
C548 _36_/a_197_47# net5 0.00254f
C549 _22_ _45_/a_27_47# 0.0131f
C550 net1 _01_ 0.0509f
C551 _08_ _03_ 0.0144f
C552 net19 p[10] 1.26e-21
C553 _45_/a_27_47# _11_ 0.0703f
C554 p[7] _40_/a_191_297# -6.82e-19
C555 _19_ net13 4.45e-20
C556 VGND _39_/a_47_47# 0.0665f
C557 _02_ _53_/a_183_297# 4.14e-19
C558 _44_/a_93_21# b[3] 7.07e-20
C559 _06_ _43_/a_27_47# 0.0329f
C560 _32_/a_27_47# _21_ 8.95e-19
C561 net1 _04_ 0.018f
C562 net13 net5 0.127f
C563 th14_0/m1_641_n318# th12_0/m1_529_n42# 0.00311f
C564 VGND net10 0.446f
C565 _43_/a_369_47# p[7] -3.75e-19
C566 b[0] p[7] 0.166f
C567 th14_0/m1_891_419# net3 2.08e-19
C568 input8/a_27_47# b[1] 0.00172f
C569 th14_0/m1_891_419# Vin 0.101f
C570 _06_ _33_/a_109_93# 6.96e-19
C571 _34_/a_129_47# b[1] 3.51e-19
C572 net7 p[13] 4.55e-19
C573 th12_0/m1_394_n856# th09_0/m1_485_n505# 4.53e-19
C574 _43_/a_193_413# p[14] 1.34e-20
C575 net6 _30_/a_215_297# 3.3e-21
C576 _18_ net15 0.0382f
C577 _14_ _20_ 0.144f
C578 _52_/a_93_21# net13 7.21e-19
C579 _33_/a_209_311# net10 0.0426f
C580 net13 b[1] 0.0495f
C581 _35_/a_489_413# _21_ 0.0448f
C582 _10_ net6 0.0965f
C583 _37_/a_197_47# net3 0.0028f
C584 _37_/a_109_47# net14 1.71e-19
C585 _10_ _13_ 0.0621f
C586 net4 _55_/a_217_297# 1.13e-19
C587 _26_/a_29_53# net15 9.06e-21
C588 net12 _36_/a_303_47# 1.37e-19
C589 _09_ net16 0.00707f
C590 _14_ p[11] 1.27e-19
C591 _35_/a_76_199# _36_/a_27_47# 3.22e-19
C592 p[12] net5 0.00392f
C593 _50_/a_223_47# _17_ 5.24e-20
C594 VGND _44_/a_93_21# -0.0223f
C595 VGND _38_/a_197_47# 2.29e-19
C596 th15_0/Vin th09_0/m1_485_n505# 0.00438f
C597 _25_ _36_/a_197_47# 2.37e-21
C598 _42_/a_368_53# net19 5.12e-19
C599 b[3] net15 0.00264f
C600 VGND th11_0/m1_705_187# 0.01f
C601 _07_ _48_/a_27_47# 0.0524f
C602 p[0] p[7] 0.27f
C603 p[7] _43_/a_27_47# 0.0186f
C604 _43_/a_469_47# net15 7.41e-19
C605 _13_ th13_0/m1_831_275# 6e-20
C606 input3/a_27_47# net19 0.00105f
C607 _09_ _21_ 0.263f
C608 th15_0/Vin net5 0.00138f
C609 th15_0/Vin input14/a_27_47# 0.00489f
C610 _52_/a_250_297# net11 1.2e-19
C611 net10 output17/a_27_47# 1.31e-20
C612 p[7] _33_/a_109_93# -0.0076f
C613 _25_ net13 0.00297f
C614 _09_ _35_/a_226_47# 0.0599f
C615 _03_ net14 1.5e-19
C616 net6 _50_/a_515_93# 4.7e-19
C617 _10_ _50_/a_429_93# 0.00167f
C618 net17 net3 3.72e-19
C619 Vin net17 0.00133f
C620 _14_ net8 4.23e-19
C621 _17_ _37_/a_303_47# 1.23e-20
C622 _15_ p[12] 0.00116f
C623 net6 _53_/a_29_53# 2.11e-20
C624 _13_ _53_/a_29_53# 9.05e-19
C625 th15_0/Vin b[1] 7.03e-19
C626 p[14] _16_ 1.74e-21
C627 _55_/a_472_297# _01_ 6.28e-19
C628 _04_ p[10] 8.48e-21
C629 VGND net15 0.222f
C630 _32_/a_303_47# _20_ 1.54e-19
C631 net9 input5/a_664_47# 5.29e-19
C632 _06_ _48_/a_181_47# 6.4e-19
C633 p[7] _27_/a_27_297# 0.0329f
C634 _07_ _22_ 1.19e-20
C635 net6 _42_/a_209_311# 1.32e-20
C636 net4 _16_ 2.73e-20
C637 _49_/a_75_199# input8/a_27_47# 1.99e-20
C638 th11_0/m1_705_187# output17/a_27_47# 0.00103f
C639 _15_ th15_0/Vin 0.00389f
C640 p[7] _31_/a_285_47# -2.91e-19
C641 input12/a_27_47# net11 0.00246f
C642 net5 input5/a_558_47# 0.0597f
C643 _39_/a_47_47# net16 7.7e-20
C644 net18 net11 0.00221f
C645 _54_/a_75_212# net10 7.43e-19
C646 _43_/a_193_413# _19_ 4.85e-21
C647 _49_/a_75_199# net13 3.2e-19
C648 _13_ _05_ 2.57e-20
C649 p[7] _44_/a_346_47# -8.74e-19
C650 _18_ _03_ 7.25e-23
C651 input5/a_664_47# _42_/a_209_311# 0.0124f
C652 _40_/a_297_297# net3 2.54e-19
C653 _47_/a_81_21# net15 0.00106f
C654 _43_/a_193_413# net5 1.39e-20
C655 _55_/a_217_297# net5 8.84e-20
C656 _32_/a_27_47# _01_ 0.0266f
C657 _45_/a_109_297# p[12] 5.61e-21
C658 _26_/a_29_53# _03_ 7.93e-21
C659 b[1] input5/a_558_47# 0.00214f
C660 _41_/a_59_75# p[14] 5.52e-19
C661 _12_ _17_ 0.0109f
C662 _37_/a_27_47# p[8] 9.82e-21
C663 Vin input7/a_27_47# 0.00527f
C664 net10 _21_ 0.0275f
C665 _07_ net12 0.18f
C666 _02_ b[2] 2.81e-19
C667 p[13] th12_0/m1_529_n42# 3.34e-20
C668 _06_ _35_/a_76_199# 0.00425f
C669 _41_/a_59_75# net4 1.76e-19
C670 _34_/a_47_47# net13 1.68e-19
C671 _10_ _52_/a_250_297# 0.00368f
C672 _48_/a_181_47# p[7] -2.73e-19
C673 VGND _33_/a_368_53# 2.38e-19
C674 _15_ input5/a_558_47# 0.00166f
C675 VGND _37_/a_109_47# -7.9e-19
C676 _32_/a_303_47# net8 2.22e-34
C677 b[1] _27_/a_205_297# 1.41e-19
C678 net14 _00_ 4.11e-20
C679 _32_/a_27_47# _04_ 1.43e-19
C680 _35_/a_226_47# net10 0.018f
C681 net1 p[10] 0.00387f
C682 _38_/a_197_47# net16 5.89e-19
C683 input5/a_381_47# p[13] 0.00464f
C684 _04_ input3/a_27_47# 3.55e-19
C685 net6 input4/a_75_212# 0.0271f
C686 _11_ p[14] 4.99e-20
C687 VGND _47_/a_384_47# -2.05e-19
C688 _15_ _27_/a_205_297# 5.5e-20
C689 _15_ _43_/a_193_413# 4.86e-19
C690 _06_ _08_ 0.0343f
C691 net4 _22_ 0.0866f
C692 _10_ _24_ 0.00484f
C693 _10_ _14_ 0.0571f
C694 _20_ net8 5.07e-19
C695 net4 _11_ 0.0858f
C696 _14_ _55_/a_80_21# 0.0175f
C697 _15_ _55_/a_217_297# 0.0474f
C698 _20_ _29_/a_29_53# 0.0111f
C699 net11 _20_ 0.00128f
C700 _09_ _01_ 4.69e-21
C701 _41_/a_59_75# _50_/a_343_93# 6.13e-22
C702 _45_/a_27_47# _17_ 1.16e-20
C703 VGND _03_ 0.119f
C704 _23_ b[2] 2.87e-20
C705 _16_ net5 1.99e-20
C706 p[7] _35_/a_76_199# -0.00924f
C707 _34_/a_285_47# _07_ 0.00975f
C708 _18_ _00_ 0.157f
C709 p[14] th15_0/m1_597_n912# 4.12e-21
C710 _18_ _36_/a_27_47# 5.46e-20
C711 _33_/a_209_311# _03_ 8.38e-19
C712 _09_ _04_ 0.0904f
C713 _26_/a_111_297# _00_ 3.7e-19
C714 VGND _55_/a_300_47# -0.00109f
C715 net4 th15_0/m1_597_n912# 2.43e-20
C716 _17_ input6/a_27_47# 7.13e-22
C717 net2 th11_0/m1_577_n654# 0.0079f
C718 _22_ _50_/a_343_93# 0.0597f
C719 _15_ _50_/a_615_93# 0.00183f
C720 net4 net12 2.57e-20
C721 _26_/a_29_53# _00_ 0.0466f
C722 _26_/a_29_53# _36_/a_27_47# 1.6e-19
C723 net2 _37_/a_303_47# 4.41e-19
C724 _32_/a_27_47# net1 0.0211f
C725 net19 _44_/a_93_21# 0.0074f
C726 _50_/a_343_93# _11_ 0.0384f
C727 _29_/a_29_53# _50_/a_27_47# 1.44e-20
C728 _24_ _53_/a_29_53# 0.0835f
C729 net2 th14_0/m1_641_n318# 4.8e-19
C730 net6 _45_/a_205_47# 2.59e-20
C731 _08_ p[7] -0.0145f
C732 _42_/a_296_53# b[1] 2.38e-20
C733 _45_/a_205_47# _13_ 7.51e-20
C734 _10_ _45_/a_193_297# 0.0047f
C735 _16_ b[1] 2.21e-19
C736 _07_ _48_/a_109_47# 3.01e-19
C737 net11 _50_/a_27_47# 6.05e-21
C738 _50_/a_223_47# _02_ 2.51e-20
C739 _23_ _36_/a_109_47# 3.44e-19
C740 _09_ _53_/a_111_297# 3.4e-19
C741 _19_ input2/a_27_47# 5.26e-20
C742 _30_/a_392_297# b[1] 3.99e-19
C743 _52_/a_250_297# _05_ 8.86e-22
C744 th03_0/m1_890_n844# b[1] 0.00101f
C745 net11 net8 1.5e-19
C746 _27_/a_27_297# net17 0.00181f
C747 _14_ _42_/a_209_311# 0.00142f
C748 _15_ _42_/a_296_53# 1.28e-19
C749 net11 _29_/a_29_53# 0.00514f
C750 _15_ _16_ 0.0607f
C751 _41_/a_59_75# net5 2.41e-19
C752 _48_/a_27_47# b[1] 0.00666f
C753 _52_/a_346_47# net5 7.03e-19
C754 net18 _53_/a_29_53# 0.0118f
C755 input3/a_27_47# p[8] 6.2e-19
C756 b[1] _31_/a_117_297# 0.00281f
C757 net17 _31_/a_285_47# 0.00134f
C758 _03_ output17/a_27_47# 1.94e-19
C759 _14_ _49_/a_201_297# 4.76e-21
C760 _20_ _30_/a_215_297# 6.08e-19
C761 p[0] input7/a_27_47# 5.13e-20
C762 p[9] net15 0.00302f
C763 _06_ net14 1.94e-19
C764 net1 th02_0/m1_983_133# 4.09e-19
C765 net7 _19_ 0.0458f
C766 net6 _36_/a_197_47# 6.94e-20
C767 _52_/a_93_21# _52_/a_346_47# -5.12e-20
C768 _10_ _20_ 0.179f
C769 net19 net15 0.0501f
C770 _22_ net5 0.405f
C771 _20_ _55_/a_80_21# 0.0291f
C772 input2/a_27_47# b[1] 0.014f
C773 _09_ net1 5.26e-20
C774 _52_/a_346_47# b[1] 6.37e-20
C775 _11_ net5 0.207f
C776 VGND _00_ 0.139f
C777 net7 net5 0.195f
C778 VGND _36_/a_27_47# 0.0211f
C779 _11_ input14/a_27_47# 1.42e-19
C780 _12_ net2 1.02e-20
C781 _49_/a_208_47# _19_ 7.12e-20
C782 VGND _35_/a_226_297# -4.55e-19
C783 _10_ p[11] 9.81e-21
C784 p[11] _55_/a_80_21# 9.25e-20
C785 net9 _32_/a_303_47# 0.00218f
C786 _41_/a_59_75# _15_ 0.0143f
C787 _15_ input2/a_27_47# 3.18e-20
C788 _52_/a_93_21# _22_ 0.0347f
C789 net6 net13 0.00188f
C790 _06_ _38_/a_27_47# 0.0172f
C791 _13_ net13 4e-21
C792 net14 output19/a_27_47# 0.00142f
C793 _04_ net10 0.121f
C794 p[13] input5/a_841_47# 7.34e-19
C795 _22_ b[1] 9.74e-20
C796 _54_/a_75_212# _03_ 5.45e-21
C797 net7 b[1] 0.0783f
C798 _38_/a_27_47# output18/a_27_47# 8.6e-19
C799 _27_/a_27_297# input7/a_27_47# 0.00119f
C800 _17_ _39_/a_285_47# 7.36e-21
C801 _47_/a_81_21# _00_ 0.0258f
C802 _44_/a_250_297# net14 4.24e-20
C803 net9 _20_ 0.328f
C804 _06_ _18_ 0.54f
C805 th15_0/m1_597_n912# net5 1.17e-19
C806 _45_/a_193_297# _05_ 4.84e-22
C807 _15_ _22_ 0.0236f
C808 _10_ _50_/a_27_47# 0.0154f
C809 net12 net5 0.0674f
C810 _30_/a_215_297# net8 8.14e-21
C811 _29_/a_29_53# _30_/a_215_297# 1.72e-19
C812 _49_/a_208_47# b[1] 2.93e-19
C813 p[7] net14 0.182f
C814 _06_ _26_/a_111_297# 9e-19
C815 _15_ _11_ 0.113f
C816 net7 _15_ 8.4e-20
C817 _10_ net8 5.86e-19
C818 net11 _30_/a_215_297# 1.04e-19
C819 _06_ _26_/a_29_53# 0.0135f
C820 _03_ _21_ 0.0818f
C821 _10_ _29_/a_29_53# 5.17e-19
C822 _55_/a_80_21# net8 1.84e-21
C823 net6 p[12] 0.0439f
C824 _49_/a_75_199# th03_0/m1_890_n844# 1.69e-21
C825 _13_ p[12] 8.72e-19
C826 net19 _37_/a_109_47# 1.16e-20
C827 _12_ _02_ 0.265f
C828 _04_ _44_/a_93_21# 4.47e-21
C829 VGND input13/a_27_47# 0.0471f
C830 th03_0/m1_638_n591# Vin 5.94e-20
C831 _10_ net11 0.0109f
C832 _25_ _22_ 5.39e-19
C833 _20_ _42_/a_209_311# 1.66e-20
C834 _06_ b[3] 9.96e-21
C835 input12/a_27_47# input10/a_27_47# 0.0154f
C836 b[0] _39_/a_129_47# 2.6e-20
C837 _25_ _11_ 7.05e-19
C838 net12 b[1] 0.12f
C839 net18 input10/a_27_47# 4.16e-20
C840 _35_/a_226_47# _03_ 0.028f
C841 p[7] _38_/a_27_47# -0.0142f
C842 input13/a_27_47# _33_/a_209_311# 5.85e-20
C843 net6 th15_0/Vin 0.00781f
C844 _20_ _49_/a_201_297# 5.24e-21
C845 net2 input6/a_27_47# 0.0047f
C846 p[11] _42_/a_209_311# 4.19e-19
C847 p[10] th02_0/m1_983_133# 1.21e-20
C848 _20_ _05_ 6.79e-19
C849 VGND th01_0/m1_571_n501# 8.66e-21
C850 _01_ net15 0.0314f
C851 net1 net10 0.00388f
C852 p[7] th02_0/m1_571_144# 0.0143f
C853 net2 p[13] 0.0301f
C854 _20_ _31_/a_35_297# 1.69e-19
C855 _22_ _45_/a_109_297# 0.0426f
C856 p[7] _18_ 0.0721f
C857 _34_/a_47_47# _48_/a_27_47# 4.45e-21
C858 net9 net8 0.0605f
C859 b[3] output19/a_27_47# 0.0274f
C860 net9 _29_/a_29_53# 0.0205f
C861 b[0] b[2] 0.183f
C862 _45_/a_109_297# _11_ 0.00168f
C863 _26_/a_111_297# p[7] -5.92e-20
C864 input5/a_664_47# th15_0/Vin 2.16e-19
C865 _17_ p[14] 1.07e-19
C866 net9 net11 0.136f
C867 VGND _41_/a_145_75# 4.11e-19
C868 p[7] _26_/a_29_53# 0.0356f
C869 VGND _39_/a_377_297# -6.28e-19
C870 _12_ _23_ 0.00743f
C871 _04_ net15 0.0569f
C872 _25_ net12 4.46e-20
C873 VGND _06_ 1.1f
C874 net4 _17_ 7.52e-21
C875 _44_/a_250_297# b[3] 3.45e-19
C876 _45_/a_27_47# _02_ 0.00449f
C877 net11 _53_/a_29_53# 8.31e-19
C878 _22_ _49_/a_75_199# 9.85e-21
C879 th12_0/m1_529_n42# th09_0/m1_485_n505# 0.0107f
C880 input8/a_27_47# p[1] 5.13e-20
C881 net7 _49_/a_75_199# 0.09f
C882 p[7] b[3] 0.129f
C883 _42_/a_209_311# net8 7.7e-21
C884 VGND output18/a_27_47# 0.0581f
C885 _43_/a_469_47# p[7] -2.75e-19
C886 th14_0/m1_891_419# net14 4.02e-21
C887 net1 th11_0/m1_705_187# 5.27e-20
C888 _06_ _33_/a_209_311# 0.0187f
C889 _34_/a_285_47# b[1] 0.00368f
C890 th15_0/m1_849_n157# b[3] 2.83e-20
C891 p[11] input5/a_62_47# 0.00153f
C892 VGND p[2] 0.28f
C893 _21_ _00_ 9.26e-20
C894 input14/a_27_47# th12_0/m1_529_n42# 7.48e-19
C895 _36_/a_27_47# _21_ 0.0276f
C896 net8 _49_/a_201_297# 7.3e-19
C897 _10_ _30_/a_215_297# 5.66e-20
C898 _33_/a_296_53# net10 8.22e-20
C899 input1/a_75_212# Vin 0.01f
C900 net8 _05_ 0.0146f
C901 p[13] _02_ 2.99e-19
C902 VGND output19/a_27_47# 0.0024f
C903 _29_/a_29_53# _05_ 3.79e-20
C904 Vin th11_0/m1_577_n654# 0.0926f
C905 net6 _43_/a_193_413# 2.41e-20
C906 _43_/a_193_413# _13_ 5.58e-21
C907 _06_ _47_/a_81_21# 0.0388f
C908 _34_/a_47_47# _22_ 3.9e-21
C909 _37_/a_197_47# net14 7e-19
C910 _37_/a_303_47# net3 0.00133f
C911 net11 _49_/a_201_297# 1.42e-19
C912 net8 _31_/a_35_297# 0.0408f
C913 th15_0/Vin _42_/a_109_93# 9.71e-20
C914 input5/a_381_47# net5 0.0546f
C915 _10_ _55_/a_80_21# 5.49e-19
C916 th14_0/m1_641_n318# net3 3.58e-19
C917 Vin th14_0/m1_641_n318# 0.00276f
C918 net11 _05_ 2.76e-19
C919 _48_/a_109_47# b[1] 9.32e-20
C920 _50_/a_343_93# _17_ 0.0015f
C921 VGND _38_/a_303_47# 1.78e-19
C922 VGND _44_/a_250_297# -0.00591f
C923 input15/a_27_47# input6/a_27_47# 5.3e-19
C924 th01_0/m1_991_n1219# Vin 0.0178f
C925 _45_/a_27_47# _23_ 1.74e-19
C926 VGND p[7] 1.53f
C927 _10_ th13_0/m1_831_275# 7.72e-20
C928 net9 _30_/a_465_297# 0.00138f
C929 input5/a_62_47# net8 2.05e-19
C930 net1 net15 7.44e-20
C931 _37_/a_27_47# _44_/a_93_21# 3.19e-19
C932 input5/a_381_47# b[1] 0.0023f
C933 VGND th15_0/m1_849_n157# 0.0514f
C934 _52_/a_250_297# p[12] 1.84e-20
C935 net9 _30_/a_215_297# 0.0456f
C936 VGND _32_/a_197_47# 8.12e-20
C937 p[7] _33_/a_209_311# -0.0125f
C938 _09_ _35_/a_489_413# 0.0296f
C939 _08_ _35_/a_556_47# 7.71e-19
C940 net6 _50_/a_615_93# 1.43e-19
C941 _03_ _01_ 2.85e-19
C942 net17 net14 5.43e-19
C943 _34_/a_47_47# net12 0.0385f
C944 _10_ _50_/a_515_93# 0.00129f
C945 _10_ net9 0.0438f
C946 p[8] net15 1.73e-20
C947 _42_/a_109_93# input5/a_558_47# 1.75e-19
C948 th15_0/Vin p[1] 2.84e-19
C949 p[7] _47_/a_81_21# 0.0089f
C950 _19_ _17_ 8.82e-21
C951 _10_ _53_/a_29_53# 0.00779f
C952 p[7] th10_0/m1_502_n495# 0.0291f
C953 _12_ net3 3.09e-20
C954 _12_ Vin 2.56e-21
C955 _55_/a_300_47# _01_ 0.00113f
C956 _47_/a_81_21# th15_0/m1_849_n157# 4.9e-19
C957 _35_/a_226_47# input13/a_27_47# 3.94e-20
C958 input10/a_27_47# net11 0.112f
C959 _04_ _03_ 0.586f
C960 _17_ net5 0.00408f
C961 net6 _16_ 1.62e-20
C962 _55_/a_80_21# _42_/a_209_311# 0.0175f
C963 _54_/a_75_212# _06_ 0.00727f
C964 th11_0/m1_705_187# p[10] 0.0622f
C965 _14_ th15_0/Vin 0.00355f
C966 _37_/a_27_47# net15 0.0541f
C967 _30_/a_215_297# _05_ 0.0453f
C968 p[7] output17/a_27_47# 0.0268f
C969 _02_ _39_/a_285_47# 0.0019f
C970 _06_ net16 0.0511f
C971 _30_/a_215_297# _31_/a_35_297# 6.37e-19
C972 _54_/a_75_212# output18/a_27_47# 2.28e-19
C973 _07_ _02_ 0.0083f
C974 _10_ _05_ 9.25e-21
C975 p[7] _44_/a_584_47# -2.28e-19
C976 _32_/a_27_47# net10 2.76e-20
C977 _47_/a_299_297# net15 1.44e-20
C978 net2 p[14] 5.39e-19
C979 output18/a_27_47# net16 3.45e-19
C980 p[1] input5/a_558_47# 1.61e-21
C981 _06_ _21_ 0.143f
C982 _55_/a_80_21# _31_/a_35_297# 5.9e-21
C983 _44_/a_256_47# p[14] 6.02e-21
C984 VGND th14_0/m1_891_419# 0.00531f
C985 _45_/a_193_297# p[12] 5.2e-20
C986 input7/a_27_47# net14 3.48e-19
C987 _15_ _17_ 0.0752f
C988 _20_ net13 5.95e-19
C989 output18/a_27_47# _21_ 0.00103f
C990 p[0] input1/a_75_212# 0.0197f
C991 _06_ _35_/a_226_47# 0.00487f
C992 _41_/a_59_75# net6 0.0373f
C993 _10_ _52_/a_256_47# 1.65e-19
C994 p[10] net15 0.00989f
C995 b[1] _27_/a_277_297# 1.24e-19
C996 p[7] th13_0/m1_559_n458# 0.0186f
C997 VGND _37_/a_197_47# -4.58e-19
C998 VGND _49_/a_315_47# -0.0034f
C999 _01_ _00_ 0.00124f
C1000 _35_/a_489_413# net10 0.00225f
C1001 _54_/a_75_212# p[7] 0.0475f
C1002 net1 _03_ 0.298f
C1003 _38_/a_303_47# net16 6.47e-19
C1004 net9 _05_ 0.124f
C1005 _06_ p[9] 0.00205f
C1006 _23_ _39_/a_285_47# 1.9e-20
C1007 net3 input6/a_27_47# 2.52e-19
C1008 Vin input6/a_27_47# 0.00242f
C1009 _09_ _39_/a_47_47# 7.7e-21
C1010 th01_0/m1_991_n1219# p[0] 0.172f
C1011 _10_ input4/a_75_212# 0.00346f
C1012 p[7] net16 0.518f
C1013 input5/a_841_47# net5 0.0221f
C1014 _07_ _23_ 1.27e-19
C1015 _14_ _43_/a_193_413# 0.0297f
C1016 b[0] _12_ 2.61e-20
C1017 input5/a_664_47# input2/a_27_47# 4.47e-21
C1018 net6 _22_ 0.163f
C1019 _22_ _13_ 0.00309f
C1020 _06_ net19 0.00522f
C1021 p[13] net3 9.08e-19
C1022 Vin p[13] 0.242f
C1023 net6 _11_ 0.0257f
C1024 _14_ _55_/a_217_297# 0.0116f
C1025 _04_ _00_ 1.98e-20
C1026 _04_ _36_/a_27_47# 0.00169f
C1027 _13_ _11_ 0.164f
C1028 net2 _50_/a_343_93# 1.25e-20
C1029 _09_ net10 0.037f
C1030 VGND _29_/a_111_297# -1.9e-19
C1031 input8/a_27_47# net8 0.0181f
C1032 p[7] _21_ 0.871f
C1033 _04_ _35_/a_226_297# 4.51e-19
C1034 _50_/a_27_47# net13 7.27e-21
C1035 th12_0/m1_394_n856# p[11] 9.12e-21
C1036 net4 _02_ 0.00376f
C1037 input11/a_27_47# p[7] 0.151f
C1038 _45_/a_109_297# _17_ 4.29e-22
C1039 _34_/a_129_47# net11 0.00242f
C1040 net9 input5/a_62_47# 3.12e-19
C1041 p[9] output19/a_27_47# 0.0933f
C1042 VGND net17 0.212f
C1043 input5/a_841_47# b[1] 7.07e-19
C1044 net13 net8 7.51e-20
C1045 _29_/a_29_53# net13 0.00104f
C1046 p[7] _35_/a_226_47# 0.00194f
C1047 net7 input5/a_664_47# 0.00199f
C1048 net19 output19/a_27_47# 0.0273f
C1049 input15/a_27_47# p[14] 0.00367f
C1050 net11 net13 0.093f
C1051 _26_/a_183_297# _00_ 4.53e-19
C1052 _49_/a_201_297# _31_/a_35_297# 5.52e-20
C1053 _12_ _43_/a_27_47# 2.33e-21
C1054 _19_ _31_/a_285_297# 1.34e-19
C1055 _33_/a_209_311# net17 7.03e-21
C1056 net6 th15_0/m1_597_n912# 1.34e-20
C1057 _05_ _31_/a_35_297# 0.00649f
C1058 net6 net12 0.00643f
C1059 p[7] p[9] 0.429f
C1060 th15_0/Vin p[11] 0.186f
C1061 output18/a_27_47# output16/a_27_47# 7.85e-19
C1062 net19 _44_/a_250_297# 0.00592f
C1063 input3/a_27_47# net15 6.19e-20
C1064 net2 _19_ 0.101f
C1065 p[12] _50_/a_27_47# 1.55e-19
C1066 net6 _45_/a_465_47# 6.06e-20
C1067 _45_/a_465_47# _13_ 0.00134f
C1068 _10_ _45_/a_205_47# 6.19e-20
C1069 _12_ _33_/a_109_93# 9.75e-20
C1070 th10_0/m1_536_174# p[14] 3.8e-19
C1071 VGND input9/a_75_212# 0.063f
C1072 p[7] net19 0.189f
C1073 p[1] th03_0/m1_890_n844# 0.00745f
C1074 _50_/a_343_93# _02_ 6.94e-19
C1075 net2 net5 0.0616f
C1076 net2 input14/a_27_47# 0.0235f
C1077 net1 _00_ 9.43e-19
C1078 net1 _36_/a_27_47# 6.99e-20
C1079 _22_ _42_/a_109_93# 1.21e-19
C1080 _14_ _16_ 0.0584f
C1081 VGND _40_/a_297_297# -5.1e-19
C1082 th15_0/Vin _50_/a_27_47# 2.06e-19
C1083 _52_/a_584_47# net5 0.0022f
C1084 _03_ p[10] 8.74e-20
C1085 b[1] _31_/a_285_297# 0.0101f
C1086 _39_/a_47_47# net10 4.72e-22
C1087 output17/a_27_47# net17 0.0149f
C1088 th15_0/Vin net8 1.56e-21
C1089 VGND input7/a_27_47# 0.0575f
C1090 p[7] output16/a_27_47# 0.123f
C1091 VGND _53_/a_183_297# -4.34e-19
C1092 net2 b[1] 0.0389f
C1093 _06_ _01_ 0.00157f
C1094 _43_/a_193_413# _20_ 0.00161f
C1095 p[1] input2/a_27_47# 0.012f
C1096 _10_ _36_/a_197_47# 1.54e-19
C1097 _20_ _55_/a_217_297# 0.0013f
C1098 net13 _30_/a_465_297# 6.36e-20
C1099 _19_ _02_ 0.213f
C1100 _15_ net2 9.8e-19
C1101 _43_/a_193_413# p[11] 8.34e-20
C1102 net13 _30_/a_215_297# 0.0246f
C1103 _32_/a_109_47# p[7] 0.00124f
C1104 p[2] _01_ 0.00164f
C1105 _06_ _04_ 0.0132f
C1106 VGND _35_/a_556_47# 1.95e-19
C1107 p[11] _55_/a_217_297# 1.6e-20
C1108 _02_ net5 0.233f
C1109 _52_/a_250_297# _22_ 0.0996f
C1110 _37_/a_27_47# _00_ 6.15e-20
C1111 _10_ net13 0.00151f
C1112 p[0] p[13] 2.15e-19
C1113 net7 p[1] 0.00514f
C1114 net1 input13/a_27_47# 1.9e-19
C1115 net8 input5/a_558_47# 0.00357f
C1116 p[2] _04_ 2.84e-20
C1117 _47_/a_299_297# _00_ 7.59e-21
C1118 _52_/a_93_21# _02_ 0.0962f
C1119 _20_ _50_/a_615_93# 8.8e-19
C1120 _06_ _53_/a_111_297# 3.82e-19
C1121 _32_/a_27_47# _03_ 1.9e-19
C1122 _22_ _24_ 0.0846f
C1123 _30_/a_109_53# net5 5.84e-22
C1124 _14_ _22_ 0.00449f
C1125 _02_ b[1] 0.00718f
C1126 _24_ _11_ 7.29e-20
C1127 net9 input8/a_27_47# 3.71e-20
C1128 th10_0/m1_536_174# th09_0/m1_485_n505# 0.00429f
C1129 p[7] _01_ 0.521f
C1130 _06_ _26_/a_183_297# 3.16e-19
C1131 _14_ _11_ 0.0415f
C1132 net7 _14_ 0.00251f
C1133 _43_/a_193_413# net8 1.62e-20
C1134 p[14] net3 0.00504f
C1135 Vin p[14] 0.143f
C1136 _10_ p[12] 0.0134f
C1137 _32_/a_197_47# _01_ 0.00156f
C1138 _04_ _44_/a_250_297# 5.57e-21
C1139 _15_ _02_ 0.101f
C1140 net9 net13 0.035f
C1141 net4 net3 9.28e-21
C1142 net4 Vin 4.16e-19
C1143 net18 _22_ 1.68e-19
C1144 _39_/a_47_47# net15 9.44e-22
C1145 _20_ _16_ 0.00271f
C1146 _23_ net5 0.0052f
C1147 p[7] _04_ 0.46f
C1148 _30_/a_109_53# b[1] 0.00655f
C1149 b[0] _39_/a_285_47# 1.88e-19
C1150 p[13] _27_/a_27_297# 2.6e-19
C1151 _35_/a_489_413# _03_ 0.0205f
C1152 VGND _49_/a_544_297# -0.00256f
C1153 p[7] _38_/a_109_47# -4.66e-19
C1154 p[12] th13_0/m1_831_275# 0.00668f
C1155 _06_ net1 0.0115f
C1156 _15_ _28_/a_109_297# 0.00346f
C1157 _20_ th03_0/m1_890_n844# 3.1e-19
C1158 _10_ th15_0/Vin 0.00935f
C1159 p[11] _16_ 1.76e-19
C1160 _25_ _02_ 0.0156f
C1161 input8/a_27_47# _49_/a_201_297# 2.46e-21
C1162 _15_ input15/a_27_47# 2.15e-20
C1163 _12_ _35_/a_76_199# 6.84e-20
C1164 _52_/a_93_21# _23_ 0.0166f
C1165 input9/a_75_212# _21_ 1.17e-21
C1166 input8/a_27_47# _05_ 1.58e-19
C1167 _53_/a_111_297# p[7] 1.11e-34
C1168 _23_ b[1] 7.65e-19
C1169 _22_ _45_/a_193_297# 0.0234f
C1170 _09_ _03_ 0.326f
C1171 net1 p[2] 0.0277f
C1172 input8/a_27_47# _31_/a_35_297# 0.00955f
C1173 _45_/a_193_297# _11_ 0.0292f
C1174 net19 net17 8.84e-23
C1175 th15_0/Vin th13_0/m1_831_275# 0.00711f
C1176 _26_/a_183_297# p[7] -3.03e-19
C1177 net13 _49_/a_201_297# 3.31e-19
C1178 input12/a_27_47# net12 0.0297f
C1179 VGND _39_/a_129_47# -0.00126f
C1180 _50_/a_223_47# net14 5.89e-21
C1181 net13 _05_ 0.192f
C1182 _45_/a_109_297# _02_ 8.44e-19
C1183 net6 _17_ 3.12e-19
C1184 _41_/a_59_75# _20_ 1.78e-20
C1185 net13 _31_/a_35_297# 1.86e-20
C1186 _44_/a_93_21# net15 0.00573f
C1187 input5/a_381_47# _42_/a_109_93# 0.00763f
C1188 _32_/a_27_47# _00_ 0.00228f
C1189 net8 _16_ 0.00624f
C1190 net6 _40_/a_109_297# 2.53e-20
C1191 _32_/a_27_47# _36_/a_27_47# 0.011f
C1192 p[8] output19/a_27_47# 0.0094f
C1193 _06_ _37_/a_27_47# 2.5e-20
C1194 _06_ _33_/a_296_53# 1.11e-20
C1195 _07_ _33_/a_109_93# 3.2e-19
C1196 net1 p[7] 1.17f
C1197 _49_/a_75_199# _02_ 0.0354f
C1198 _25_ _23_ 0.00465f
C1199 th03_0/m1_890_n844# net8 3.83e-19
C1200 _22_ _20_ 0.183f
C1201 _33_/a_368_53# net10 0.00171f
C1202 VGND b[2] 0.0779f
C1203 _45_/a_27_47# _35_/a_76_199# 2.04e-21
C1204 _20_ _11_ 0.268f
C1205 net6 _43_/a_297_47# 8.23e-22
C1206 net7 _20_ 0.0257f
C1207 th01_0/m1_571_n501# p[10] 0.006f
C1208 _06_ _47_/a_299_297# 0.0174f
C1209 b[0] net4 0.0024f
C1210 _10_ _43_/a_193_413# 0.0174f
C1211 _35_/a_556_47# _21_ 2.69e-19
C1212 _37_/a_303_47# net14 0.00112f
C1213 net1 _32_/a_197_47# 0.00142f
C1214 Vin th09_0/m1_485_n505# 0.134f
C1215 _43_/a_193_413# _55_/a_80_21# 2.54e-19
C1216 net8 _31_/a_117_297# 5.91e-19
C1217 _49_/a_315_47# _01_ 1.82e-19
C1218 th15_0/Vin _42_/a_209_311# 2.47e-20
C1219 _10_ _55_/a_217_297# 1.43e-19
C1220 _19_ net3 0.0129f
C1221 th14_0/m1_641_n318# net14 0.00168f
C1222 Vin _19_ 0.00421f
C1223 p[7] p[8] 0.267f
C1224 _55_/a_80_21# _55_/a_217_297# 1.42e-32
C1225 net11 _48_/a_27_47# 0.0179f
C1226 _22_ p[11] 3.13e-20
C1227 _50_/a_223_47# _18_ 0.0367f
C1228 _41_/a_59_75# _50_/a_27_47# 9.59e-22
C1229 net3 net5 0.0365f
C1230 _34_/a_47_47# _02_ 1.09e-19
C1231 input14/a_27_47# net3 9.36e-19
C1232 Vin input14/a_27_47# 4.64e-19
C1233 _39_/a_47_47# _03_ 1.47e-19
C1234 net9 input5/a_558_47# 4.42e-19
C1235 _50_/a_223_47# _26_/a_29_53# 0.00124f
C1236 _49_/a_315_47# _04_ 7.71e-19
C1237 input2/a_27_47# net8 0.0207f
C1238 _09_ _00_ 9.35e-21
C1239 VGND _36_/a_109_47# 3.56e-19
C1240 VGND th03_0/m1_638_n591# 0.00102f
C1241 _03_ net10 0.321f
C1242 net12 _20_ 0.00437f
C1243 p[7] _33_/a_296_53# -1.15e-19
C1244 _22_ _50_/a_27_47# 0.0276f
C1245 p[7] _37_/a_27_47# -0.0178f
C1246 _17_ _42_/a_109_93# 7.83e-20
C1247 _09_ _35_/a_226_297# 4.98e-19
C1248 _50_/a_27_47# _11_ 0.0592f
C1249 net17 _01_ 0.0988f
C1250 b[1] net3 0.00334f
C1251 _34_/a_377_297# net12 0.00251f
C1252 _10_ _50_/a_615_93# 8.82e-19
C1253 Vin b[1] 0.0677f
C1254 input4/a_75_212# p[12] 0.0278f
C1255 _14_ input5/a_381_47# 5.68e-20
C1256 _22_ net8 3.3e-20
C1257 _42_/a_209_311# input5/a_558_47# 7.85e-20
C1258 _22_ _29_/a_29_53# 2.24e-21
C1259 _04_ _29_/a_111_297# 9.25e-19
C1260 _11_ net8 1.81e-20
C1261 net7 net8 0.295f
C1262 th15_0/Vin input5/a_62_47# 9.04e-19
C1263 p[7] _47_/a_299_297# 0.0643f
C1264 net7 _29_/a_29_53# 6.01e-19
C1265 _22_ net11 6.82e-21
C1266 th01_0/m1_991_n1219# th02_0/m1_571_144# 0.00603f
C1267 _15_ net3 0.224f
C1268 VGND _30_/a_297_297# -5.13e-19
C1269 net7 net11 1.77e-19
C1270 _04_ net17 0.0218f
C1271 _07_ _48_/a_181_47# 5.93e-19
C1272 _49_/a_208_47# net8 1.4e-19
C1273 th15_0/Vin input4/a_75_212# 0.00104f
C1274 _10_ _16_ 0.00486f
C1275 _55_/a_80_21# _16_ 0.0143f
C1276 p[7] p[10] 0.433f
C1277 net12 _50_/a_27_47# 7.99e-21
C1278 VGND _50_/a_223_47# 0.0159f
C1279 _06_ _32_/a_27_47# 0.00663f
C1280 _09_ input13/a_27_47# 1.27e-21
C1281 _12_ _38_/a_27_47# 0.0527f
C1282 net12 net8 0.00458f
C1283 _10_ _48_/a_27_47# 4.55e-19
C1284 net12 _29_/a_29_53# 0.0132f
C1285 _55_/a_472_297# p[7] 0.00488f
C1286 b[0] net5 3.39e-19
C1287 _04_ input9/a_75_212# 7.69e-22
C1288 net12 net11 0.358f
C1289 _39_/a_47_47# _00_ 1.85e-20
C1290 th01_0/m1_571_n501# th02_0/m1_983_133# 7.11e-20
C1291 net6 net2 0.00139f
C1292 _12_ _18_ 0.0115f
C1293 input2/a_27_47# _30_/a_215_297# 3.51e-20
C1294 _14_ _17_ 0.489f
C1295 net13 _36_/a_197_47# 1.06e-19
C1296 VGND input1/a_75_212# 0.0586f
C1297 p[1] _27_/a_277_297# 1.66e-20
C1298 _06_ _35_/a_489_413# 9.22e-19
C1299 _07_ _35_/a_76_199# 0.00226f
C1300 VGND th11_0/m1_577_n654# 0.0025f
C1301 _36_/a_27_47# net10 0.0366f
C1302 _10_ _41_/a_59_75# 0.0235f
C1303 _14_ _40_/a_109_297# -1.78e-33
C1304 _12_ _26_/a_29_53# 0.00243f
C1305 VGND _37_/a_303_47# -1.63e-19
C1306 _03_ net15 4.26e-20
C1307 input3/a_27_47# output19/a_27_47# 4.77e-21
C1308 net9 _30_/a_392_297# 9.92e-19
C1309 b[2] _21_ 2.14e-19
C1310 VGND th14_0/m1_641_n318# 0.00635f
C1311 _35_/a_226_297# net10 2.48e-19
C1312 input5/a_664_47# net2 8.11e-20
C1313 net1 net17 2.89e-19
C1314 _22_ _30_/a_215_297# 2.46e-21
C1315 _49_/a_75_199# net3 2.01e-19
C1316 net14 input6/a_27_47# 7.05e-19
C1317 th01_0/m1_991_n1219# VGND 6.29e-19
C1318 _32_/a_27_47# p[7] 0.0395f
C1319 _55_/a_300_47# net15 1.09e-19
C1320 _06_ _09_ 0.0965f
C1321 _42_/a_209_311# _16_ 0.00129f
C1322 _14_ _43_/a_297_47# 9.11e-19
C1323 input3/a_27_47# _44_/a_250_297# 2.07e-19
C1324 _07_ _08_ 0.348f
C1325 p[7] _42_/a_368_53# -3.03e-19
C1326 _10_ _22_ 0.0904f
C1327 p[13] net14 5.58e-19
C1328 p[11] th12_0/m1_529_n42# 0.0172f
C1329 _48_/a_27_47# _53_/a_29_53# 3.14e-21
C1330 _22_ _55_/a_80_21# 0.00926f
C1331 _10_ _11_ 0.176f
C1332 p[7] input3/a_27_47# 0.0688f
C1333 _10_ net7 6.22e-20
C1334 p[2] th02_0/m1_983_133# 9.44e-20
C1335 net7 _55_/a_80_21# 0.00163f
C1336 _44_/a_93_21# _00_ 4.54e-20
C1337 net6 _02_ 0.00427f
C1338 th14_0/m1_891_419# p[10] 5.19e-20
C1339 _13_ _02_ 0.0676f
C1340 _45_/a_27_47# _18_ 0.00347f
C1341 net1 input9/a_75_212# 0.002f
C1342 p[0] b[1] 0.00454f
C1343 net12 _30_/a_465_297# 8.01e-20
C1344 p[7] _35_/a_489_413# -0.00725f
C1345 _19_ _27_/a_27_297# 0.082f
C1346 input13/a_27_47# net10 8.86e-20
C1347 th03_0/m1_890_n844# _05_ 9.65e-20
C1348 input1/a_75_212# output17/a_27_47# 0.0101f
C1349 _52_/a_93_21# _33_/a_109_93# 2.89e-21
C1350 net2 _42_/a_109_93# 0.00507f
C1351 net12 _30_/a_215_297# 0.00676f
C1352 VGND _12_ 0.816f
C1353 th03_0/m1_890_n844# _31_/a_35_297# 4.56e-19
C1354 _33_/a_109_93# b[1] 0.00411f
C1355 _15_ _43_/a_27_47# 8.96e-20
C1356 input5/a_664_47# _02_ 0.00187f
C1357 p[7] th02_0/m1_983_133# 0.0376f
C1358 _27_/a_27_297# net5 3.48e-19
C1359 net6 input15/a_27_47# 0.146f
C1360 net11 _48_/a_109_47# 1.74e-19
C1361 net9 _22_ 0.0023f
C1362 _10_ net12 0.00257f
C1363 _42_/a_209_311# input2/a_27_47# 1e-22
C1364 net9 _11_ 5.39e-19
C1365 net9 net7 0.00233f
C1366 _49_/a_544_297# _01_ 0.00109f
C1367 _09_ p[7] 0.297f
C1368 _22_ _53_/a_29_53# 0.00749f
C1369 net1 input7/a_27_47# 0.0383f
C1370 _10_ _45_/a_465_47# 3.32e-19
C1371 _12_ _33_/a_209_311# 2.88e-20
C1372 input5/a_381_47# net8 7.48e-19
C1373 _50_/a_223_47# net16 4.77e-21
C1374 _11_ _53_/a_29_53# 2.33e-20
C1375 net15 _00_ 0.00147f
C1376 th13_0/m1_831_275# th15_0/m1_597_n912# 0.0186f
C1377 _20_ _17_ 0.102f
C1378 input2/a_27_47# _05_ 1.83e-19
C1379 net6 _23_ 2.13e-19
C1380 b[3] input6/a_27_47# 4.02e-19
C1381 _27_/a_27_297# b[1] 0.00644f
C1382 _23_ _13_ 2.08e-20
C1383 _06_ _39_/a_47_47# 1.44e-19
C1384 _22_ _42_/a_209_311# 1.72e-19
C1385 net11 _29_/a_183_297# 3.64e-19
C1386 _12_ _47_/a_81_21# 0.00158f
C1387 _49_/a_544_297# _04_ 0.00204f
C1388 input2/a_27_47# _31_/a_35_297# 0.00136f
C1389 _20_ _40_/a_109_297# 2.35e-20
C1390 _50_/a_223_47# _21_ 2.91e-21
C1391 b[1] _31_/a_285_47# 8.76e-19
C1392 p[11] _17_ 0.00765f
C1393 net17 p[10] 0.183f
C1394 net2 p[1] 7.54e-20
C1395 th12_0/m1_394_n856# th15_0/Vin 0.0254f
C1396 _06_ net10 0.184f
C1397 _15_ _27_/a_27_297# 9.85e-20
C1398 _22_ _49_/a_201_297# 2.45e-20
C1399 net9 net12 0.0596f
C1400 th14_0/m1_891_419# input3/a_27_47# 3.77e-20
C1401 _22_ _05_ 3.33e-21
C1402 th15_0/Vin p[12] 0.175f
C1403 net7 _49_/a_201_297# 0.00419f
C1404 VGND _45_/a_27_47# -0.029f
C1405 net7 _05_ 0.0129f
C1406 th01_0/m1_571_n501# th11_0/m1_705_187# 0.00336f
C1407 net7 _31_/a_35_297# 0.0384f
C1408 VGND _36_/a_303_47# 8.14e-19
C1409 _14_ net2 0.0104f
C1410 _50_/a_27_47# _17_ 3.93e-20
C1411 _14_ _44_/a_256_47# 0.00124f
C1412 _41_/a_59_75# input4/a_75_212# 0.00153f
C1413 VGND input6/a_27_47# -0.00236f
C1414 _17_ net8 4.52e-20
C1415 _06_ _38_/a_197_47# 4.32e-19
C1416 VGND p[13] 0.153f
C1417 p[7] _39_/a_47_47# 0.0668f
C1418 _48_/a_181_47# b[1] 3.46e-19
C1419 net7 input5/a_62_47# 2.04e-19
C1420 net12 _05_ 0.0414f
C1421 _49_/a_544_297# net1 0.00175f
C1422 _52_/a_250_297# _02_ 0.0128f
C1423 _47_/a_384_47# _00_ 5.15e-20
C1424 p[7] net10 0.393f
C1425 input7/a_27_47# p[10] 1.82e-19
C1426 _35_/a_76_199# net5 3.38e-19
C1427 net8 _27_/a_277_297# 7.99e-20
C1428 _44_/a_93_21# output19/a_27_47# 7.25e-20
C1429 p[14] net14 0.00278f
C1430 _12_ net16 0.131f
C1431 _09_ _49_/a_315_47# 1.11e-20
C1432 _10_ _29_/a_183_297# 6.24e-20
C1433 _24_ _02_ 0.0232f
C1434 _49_/a_75_199# _27_/a_27_297# 0.011f
C1435 _14_ _02_ 0.0316f
C1436 th15_0/Vin input5/a_558_47# 2.18e-19
C1437 _03_ _00_ 2.31e-20
C1438 net19 th14_0/m1_641_n318# 1.17e-19
C1439 net6 net3 0.00152f
C1440 net4 net14 2.21e-21
C1441 net6 Vin 6.97e-19
C1442 _44_/a_93_21# _44_/a_250_297# -6.97e-22
C1443 _52_/a_93_21# _35_/a_76_199# 6.83e-21
C1444 _06_ net15 0.033f
C1445 _12_ _21_ 7.99e-20
C1446 _35_/a_226_297# _03_ 0.00101f
C1447 _35_/a_76_199# b[1] 0.00458f
C1448 p[7] _38_/a_197_47# -5.24e-19
C1449 p[7] _44_/a_93_21# 0.005f
C1450 th15_0/Vin _43_/a_193_413# 5.52e-19
C1451 input4/a_75_212# th15_0/m1_597_n912# 8.81e-20
C1452 p[7] th11_0/m1_705_187# 0.0375f
C1453 input12/a_27_47# _02_ 1.88e-19
C1454 _14_ _28_/a_109_297# 5.66e-19
C1455 _04_ _36_/a_109_47# 2.39e-19
C1456 _09_ _29_/a_111_297# 5.79e-20
C1457 p[13] output17/a_27_47# 0.00118f
C1458 net18 _02_ 8.53e-20
C1459 net17 th02_0/m1_983_133# 1.59e-19
C1460 _14_ input15/a_27_47# 9.48e-21
C1461 input5/a_664_47# net3 0.00215f
C1462 input8/a_27_47# th03_0/m1_890_n844# 0.00179f
C1463 _12_ _35_/a_226_47# 8.38e-20
C1464 _52_/a_250_297# _23_ 3.17e-19
C1465 input5/a_841_47# net8 0.025f
C1466 input10/a_27_47# net12 0.00115f
C1467 _34_/a_285_47# _05_ 7.85e-21
C1468 net4 _38_/a_27_47# 0.0119f
C1469 net9 input5/a_381_47# 3.4e-19
C1470 _08_ b[1] 0.0127f
C1471 net9 _29_/a_183_297# 3.51e-19
C1472 net15 output19/a_27_47# 6.88e-19
C1473 net13 _30_/a_392_297# 6.64e-20
C1474 _20_ net2 8.83e-19
C1475 _18_ p[14] 2.75e-20
C1476 _50_/a_343_93# net14 1.07e-20
C1477 VGND _39_/a_285_47# -0.0046f
C1478 _45_/a_27_47# net16 8.68e-19
C1479 _24_ _23_ 0.012f
C1480 net4 _18_ 0.023f
C1481 _45_/a_193_297# _02_ 0.00988f
C1482 VGND _07_ 0.195f
C1483 _10_ _17_ 0.0233f
C1484 _44_/a_250_297# net15 8.86e-20
C1485 _55_/a_80_21# _17_ 7.64e-21
C1486 net2 p[11] 0.00681f
C1487 input5/a_381_47# _42_/a_209_311# 3.88e-19
C1488 net6 _40_/a_191_297# 1.16e-20
C1489 p[7] net15 0.61f
C1490 _45_/a_27_47# _21_ 1.18e-20
C1491 net4 _26_/a_29_53# 0.00412f
C1492 _06_ _33_/a_368_53# 1.7e-19
C1493 _07_ _33_/a_209_311# 0.00859f
C1494 _04_ _50_/a_223_47# 7.89e-22
C1495 p[14] b[3] 0.0451f
C1496 net18 _23_ -4.05e-24
C1497 _32_/a_303_47# _02_ 1.15e-20
C1498 _42_/a_109_93# net3 0.0435f
C1499 _45_/a_27_47# _35_/a_226_47# 5.71e-21
C1500 net6 _43_/a_369_47# 3.62e-21
C1501 _10_ _43_/a_297_47# 0.00118f
C1502 b[0] net6 2.52e-19
C1503 net8 _31_/a_285_297# 0.0215f
C1504 b[0] _13_ 0.00299f
C1505 th15_0/Vin _42_/a_296_53# 7.75e-21
C1506 th15_0/Vin _16_ 5.12e-19
C1507 net7 input8/a_27_47# 1.47e-19
C1508 _19_ net14 0.0512f
C1509 _20_ _02_ 0.1f
C1510 _50_/a_343_93# _18_ 0.0276f
C1511 net9 _17_ 2.89e-23
C1512 net2 net8 0.0525f
C1513 th14_0/m1_891_419# th11_0/m1_705_187# 1.31e-19
C1514 _09_ _53_/a_183_297# 4.18e-19
C1515 _22_ net13 4.63e-20
C1516 th15_0/Vin th03_0/m1_890_n844# 4.95e-20
C1517 _45_/a_193_297# _23_ 4.13e-19
C1518 net14 net5 0.0263f
C1519 _04_ th11_0/m1_577_n654# 4.01e-19
C1520 input14/a_27_47# net14 0.0232f
C1521 net7 net13 1.72e-19
C1522 _50_/a_343_93# _26_/a_29_53# 2.61e-19
C1523 _06_ _03_ 0.00635f
C1524 net1 _30_/a_297_297# 7.34e-20
C1525 _41_/a_59_75# p[12] 0.0048f
C1526 VGND p[14] 0.619f
C1527 _20_ _28_/a_109_297# 0.00221f
C1528 _20_ _30_/a_109_53# 8.12e-19
C1529 p[9] input6/a_27_47# 0.0756f
C1530 net10 net17 8.67e-21
C1531 p[1] net3 1.67e-20
C1532 p[7] _37_/a_109_47# -4.38e-19
C1533 _17_ _42_/a_209_311# 1.22e-19
C1534 net12 _36_/a_197_47# 4.67e-20
C1535 p[7] _33_/a_368_53# -4.26e-19
C1536 Vin p[1] 0.175f
C1537 VGND net4 0.564f
C1538 net6 _43_/a_27_47# 9.07e-20
C1539 _09_ _35_/a_556_47# 0.00122f
C1540 _43_/a_27_47# _13_ 1.66e-20
C1541 _06_ _55_/a_300_47# 2.5e-20
C1542 b[1] net14 0.00256f
C1543 p[2] _03_ 2.16e-20
C1544 net19 input6/a_27_47# 0.00574f
C1545 _38_/a_27_47# net5 1.76e-19
C1546 _41_/a_59_75# th15_0/Vin 0.00218f
C1547 _22_ p[12] 4.34e-21
C1548 p[7] _47_/a_384_47# -1.45e-19
C1549 _50_/a_27_47# _02_ 2.09e-19
C1550 p[12] _11_ 3.66e-20
C1551 net12 net13 0.363f
C1552 th14_0/m1_891_419# net15 3.54e-21
C1553 _15_ net14 0.225f
C1554 _14_ net3 0.0295f
C1555 _14_ Vin 3.46e-19
C1556 _47_/a_81_21# p[14] 1.42e-21
C1557 _18_ net5 0.0426f
C1558 _02_ net8 0.334f
C1559 _43_/a_193_413# _16_ 0.0261f
C1560 _29_/a_29_53# _02_ 6.76e-21
C1561 input9/a_75_212# net10 0.00699f
C1562 _34_/a_47_47# _08_ 0.00123f
C1563 _55_/a_217_297# _16_ 0.0017f
C1564 b[3] th09_0/m1_485_n505# 2.57e-19
C1565 th11_0/m1_705_187# net17 1.25e-19
C1566 net11 _02_ 0.0327f
C1567 net1 input1/a_75_212# 0.00208f
C1568 _39_/a_285_47# net16 1.29e-19
C1569 _26_/a_29_53# net5 0.0237f
C1570 _37_/a_197_47# net15 1.78e-19
C1571 p[7] _03_ 0.839f
C1572 net7 th15_0/Vin 1.02e-19
C1573 th15_0/Vin _11_ 0.00308f
C1574 _12_ _04_ 1.42e-19
C1575 VGND _50_/a_343_93# -3.89e-19
C1576 net9 input5/a_841_47# 2.7e-19
C1577 _52_/a_93_21# _18_ 1.97e-19
C1578 _12_ _38_/a_109_47# 0.00179f
C1579 net8 _30_/a_109_53# 1.76e-20
C1580 _29_/a_29_53# _30_/a_109_53# 0.0103f
C1581 p[12] th15_0/m1_597_n912# 0.0395f
C1582 input14/a_27_47# b[3] 0.00268f
C1583 _55_/a_300_47# p[7] -4.61e-19
C1584 input2/a_27_47# input5/a_558_47# 2.04e-20
C1585 _09_ _49_/a_544_297# 2.56e-20
C1586 _07_ _21_ 0.133f
C1587 net2 _27_/a_109_297# 7.24e-20
C1588 _06_ _00_ 0.1f
C1589 _26_/a_29_53# b[1] 9.93e-21
C1590 _06_ _36_/a_27_47# 0.0501f
C1591 _10_ net2 3.15e-19
C1592 input5/a_664_47# _27_/a_27_297# 0.0116f
C1593 _15_ _18_ 0.042f
C1594 _25_ _38_/a_27_47# 5.76e-19
C1595 _06_ _35_/a_226_297# 1.28e-19
C1596 _07_ _35_/a_226_47# 8.96e-19
C1597 _47_/a_81_21# _50_/a_343_93# 0.00282f
C1598 _47_/a_299_297# _50_/a_223_47# 2.74e-20
C1599 th15_0/Vin th15_0/m1_597_n912# 0.00183f
C1600 _34_/a_285_47# net13 4.11e-20
C1601 _14_ _40_/a_191_297# 2.4e-19
C1602 VGND th09_0/m1_485_n505# 0.00241f
C1603 net17 net15 5.19e-19
C1604 _15_ _26_/a_29_53# 0.00192f
C1605 _35_/a_556_47# net10 5.59e-19
C1606 VGND _19_ 0.379f
C1607 net11 _23_ 0.0461f
C1608 net7 input5/a_558_47# 0.00358f
C1609 _49_/a_75_199# net14 3.67e-19
C1610 VGND net5 1.2f
C1611 _22_ _43_/a_193_413# 0.00133f
C1612 VGND input14/a_27_47# 0.0389f
C1613 _14_ _43_/a_369_47# 0.00135f
C1614 th11_0/m1_705_187# input7/a_27_47# 1.5e-20
C1615 p[13] _01_ 4.28e-19
C1616 _43_/a_193_413# _11_ 5.45e-19
C1617 net7 _43_/a_193_413# 3.49e-19
C1618 net9 net2 3.64e-20
C1619 _02_ _30_/a_215_297# 3.58e-21
C1620 net7 _55_/a_217_297# 1.04e-19
C1621 _44_/a_250_297# _00_ 6.39e-20
C1622 _27_/a_27_297# _42_/a_109_93# 1.35e-20
C1623 net4 net16 0.155f
C1624 _20_ net3 4.07e-19
C1625 p[0] p[1] 0.0399f
C1626 th10_0/m1_502_n495# th09_0/m1_485_n505# 7.17e-20
C1627 VGND _52_/a_93_21# -0.0175f
C1628 _10_ _02_ 0.0537f
C1629 p[7] _00_ 0.416f
C1630 p[7] _36_/a_27_47# -0.00832f
C1631 _06_ input13/a_27_47# 4.89e-19
C1632 _55_/a_80_21# _02_ 0.164f
C1633 VGND b[1] 0.562f
C1634 _04_ p[13] 0.00111f
C1635 _09_ b[2] 4.28e-20
C1636 p[7] _35_/a_226_297# -8.38e-19
C1637 input1/a_75_212# p[10] 0.00136f
C1638 net4 _21_ 0.00535f
C1639 _47_/a_81_21# net5 4.59e-19
C1640 _40_/a_297_297# net15 4.08e-19
C1641 p[11] net3 0.00765f
C1642 p[11] Vin 0.00572f
C1643 th11_0/m1_577_n654# p[10] 4.13e-19
C1644 _52_/a_250_297# _33_/a_109_93# 5.17e-22
C1645 net2 _42_/a_209_311# 5.1e-19
C1646 _10_ _28_/a_109_297# 4.34e-19
C1647 _33_/a_209_311# b[1] 0.0129f
C1648 VGND _15_ 0.15f
C1649 th12_0/m1_394_n856# th12_0/m1_529_n42# 1.78e-33
C1650 _49_/a_315_47# _03_ 9.22e-19
C1651 _14_ _43_/a_27_47# 0.00938f
C1652 _55_/a_80_21# _28_/a_109_297# 2.05e-20
C1653 _05_ _31_/a_285_297# 6.12e-19
C1654 _19_ output17/a_27_47# 7.69e-19
C1655 input7/a_27_47# net15 1.88e-19
C1656 _10_ input15/a_27_47# 4.5e-19
C1657 net6 _35_/a_76_199# 4.6e-21
C1658 _13_ _35_/a_76_199# 3.01e-21
C1659 th01_0/m1_991_n1219# p[10] 0.00424f
C1660 net2 _05_ 4.03e-20
C1661 p[9] p[14] 0.0624f
C1662 th03_0/m1_638_n591# th02_0/m1_983_133# 0.00168f
C1663 output17/a_27_47# net5 5.01e-20
C1664 net9 _02_ 0.00611f
C1665 net2 _31_/a_35_297# 0.0635f
C1666 p[1] _27_/a_27_297# 2.87e-19
C1667 VGND _25_ 0.199f
C1668 net19 p[14] 0.06f
C1669 _03_ _29_/a_111_297# 7.48e-19
C1670 th15_0/Vin th12_0/m1_529_n42# 0.0693f
C1671 _10_ _23_ 0.00192f
C1672 _06_ _39_/a_377_297# 8.76e-20
C1673 _22_ _16_ 3.8e-19
C1674 net8 net3 9.23e-19
C1675 _02_ _53_/a_29_53# 0.0388f
C1676 Vin net8 0.0021f
C1677 _12_ _47_/a_299_297# 0.00805f
C1678 _29_/a_29_53# net3 1.68e-20
C1679 _20_ _40_/a_191_297# 2.07e-20
C1680 _15_ _47_/a_81_21# 0.00332f
C1681 _11_ _16_ 4.42e-20
C1682 net4 net19 2.65e-20
C1683 net7 _16_ 7.5e-20
C1684 p[7] input13/a_27_47# 0.0913f
C1685 _03_ net17 5.1e-19
C1686 net9 _28_/a_109_297# 3.7e-19
C1687 output17/a_27_47# b[1] 0.0373f
C1688 net2 input5/a_62_47# 0.0197f
C1689 input5/a_381_47# th15_0/Vin 3.39e-19
C1690 _14_ _27_/a_27_297# 1.66e-21
C1691 net9 _30_/a_109_53# 0.0191f
C1692 _06_ output18/a_27_47# 0.0114f
C1693 _42_/a_209_311# _02_ 9.92e-19
C1694 net1 p[13] 2.13e-19
C1695 net7 th03_0/m1_890_n844# 2.87e-19
C1696 VGND _45_/a_109_297# -0.00179f
C1697 net7 _31_/a_117_297# 0.00472f
C1698 th01_0/m1_571_n501# p[7] 0.0263f
C1699 _06_ output19/a_27_47# 1.53e-19
C1700 _42_/a_368_53# th14_0/m1_641_n318# 2.53e-20
C1701 net4 output16/a_27_47# 0.00706f
C1702 _02_ _05_ 0.00163f
C1703 _14_ _44_/a_346_47# 3.76e-19
C1704 p[13] p[8] 0.00239f
C1705 net9 _23_ 1.21e-19
C1706 input3/a_27_47# th14_0/m1_641_n318# 4.43e-19
C1707 _07_ _04_ 9.74e-20
C1708 VGND _49_/a_75_199# 5.87e-20
C1709 net16 net5 0.00476f
C1710 _02_ _31_/a_35_297# 0.00316f
C1711 input9/a_75_212# _03_ 9.32e-20
C1712 _41_/a_59_75# _22_ 6.24e-22
C1713 _41_/a_59_75# _11_ 8.7e-19
C1714 p[7] _41_/a_145_75# -2.41e-19
C1715 net7 input2/a_27_47# 0.00213f
C1716 net12 _30_/a_392_297# 2.19e-20
C1717 _06_ p[7] 1.41f
C1718 net5 _21_ 0.00784f
C1719 _54_/a_75_212# b[1] 0.0023f
C1720 _37_/a_27_47# input6/a_27_47# 9.35e-19
C1721 _30_/a_109_53# _05_ 0.033f
C1722 net12 _48_/a_27_47# 0.0126f
C1723 input1/a_75_212# th02_0/m1_983_133# 5.8e-20
C1724 _20_ _43_/a_27_47# 0.0124f
C1725 _30_/a_109_53# _31_/a_35_297# 2.89e-20
C1726 _06_ th15_0/m1_849_n157# 2.65e-19
C1727 _52_/a_256_47# _02_ 0.00344f
C1728 p[7] output18/a_27_47# 0.0689f
C1729 VGND _34_/a_47_47# 0.0892f
C1730 p[9] th09_0/m1_485_n505# 0.0164f
C1731 _22_ _11_ 0.15f
C1732 th15_0/Vin _17_ 0.00232f
C1733 net7 _22_ 2.73e-20
C1734 p[2] p[7] 0.212f
C1735 _52_/a_93_21# _21_ 9.4e-19
C1736 _44_/a_250_297# output19/a_27_47# 6.42e-20
C1737 b[1] _21_ 0.00892f
C1738 th15_0/Vin _40_/a_109_297# 7.23e-19
C1739 th01_0/m1_991_n1219# th02_0/m1_983_133# 4.16e-19
C1740 p[7] output19/a_27_47# 0.0245f
C1741 _34_/a_47_47# _33_/a_209_311# 0.017f
C1742 net3 _27_/a_109_297# 5.45e-19
C1743 Vin _27_/a_109_297# 5.3e-20
C1744 input11/a_27_47# b[1] 0.00688f
C1745 net6 net14 2.82e-21
C1746 _10_ net3 3.89e-19
C1747 input14/a_27_47# p[9] 8.53e-21
C1748 _10_ Vin 0.00189f
C1749 _52_/a_250_297# _35_/a_76_199# 3.4e-21
C1750 _52_/a_93_21# _35_/a_226_47# 4.89e-20
C1751 _55_/a_80_21# net3 2.35e-19
C1752 net7 _49_/a_208_47# 0.00312f
C1753 _54_/a_75_212# _25_ 0.0247f
C1754 _15_ _21_ 1.13e-21
C1755 _35_/a_226_47# b[1] 0.00334f
C1756 p[7] _44_/a_250_297# 0.0233f
C1757 net19 net5 0.00124f
C1758 p[7] _38_/a_303_47# -4.83e-19
C1759 net19 input14/a_27_47# 3.63e-19
C1760 _07_ net1 6.08e-22
C1761 th15_0/Vin _43_/a_297_47# 2.63e-20
C1762 net10 _30_/a_297_297# 1.68e-19
C1763 _25_ net16 1.16e-19
C1764 p[13] p[10] 0.00616f
C1765 input15/a_27_47# input4/a_75_212# 1.1e-21
C1766 _20_ _27_/a_27_297# 3.14e-20
C1767 _22_ net12 5.73e-20
C1768 Vin th13_0/m1_831_275# 0.0354f
C1769 input5/a_664_47# net14 0.0179f
C1770 _52_/a_256_47# _23_ 6.66e-19
C1771 p[7] th15_0/m1_849_n157# 0.0316f
C1772 net12 _11_ 3.82e-21
C1773 net7 net12 1.57e-19
C1774 net4 _38_/a_109_47# 7.32e-19
C1775 _17_ input5/a_558_47# 2.13e-21
C1776 _13_ _38_/a_27_47# 4.58e-19
C1777 _34_/a_285_47# _48_/a_27_47# 6.66e-20
C1778 _25_ _21_ 0.00164f
C1779 p[7] _32_/a_197_47# 0.00146f
C1780 input8/a_27_47# _31_/a_285_297# 1.04e-19
C1781 net19 b[1] 1e-19
C1782 output16/a_27_47# net5 4.14e-19
C1783 _15_ p[9] 2.06e-19
C1784 net9 net3 5.09e-20
C1785 _50_/a_343_93# _01_ 0.0131f
C1786 _50_/a_429_93# net14 6.04e-21
C1787 _45_/a_109_297# net16 5.1e-20
C1788 net4 _53_/a_111_297# 2.09e-19
C1789 _09_ _12_ 0.00526f
C1790 _43_/a_193_413# _17_ 0.0503f
C1791 net6 _18_ 0.166f
C1792 _13_ _18_ 0.019f
C1793 net13 _31_/a_285_297# 3.85e-20
C1794 _15_ net19 0.166f
C1795 net11 _33_/a_109_93# 5.14e-19
C1796 _26_/a_111_297# net6 1.12e-19
C1797 th15_0/Vin input5/a_841_47# 9.9e-20
C1798 net6 _26_/a_29_53# 0.0032f
C1799 _32_/a_109_47# net5 5.69e-21
C1800 _49_/a_544_297# _03_ 0.00568f
C1801 _42_/a_209_311# net3 0.029f
C1802 _42_/a_109_93# net14 0.00351f
C1803 input5/a_664_47# _18_ 1.09e-20
C1804 _27_/a_27_297# net8 0.0108f
C1805 net6 b[3] 8.06e-19
C1806 _32_/a_27_47# p[13] 6.49e-20
C1807 _45_/a_27_47# _35_/a_489_413# 3.89e-21
C1808 _45_/a_109_297# _35_/a_226_47# 1.59e-21
C1809 net6 _43_/a_469_47# 4.85e-21
C1810 _10_ _43_/a_369_47# 0.00199f
C1811 _49_/a_75_199# _21_ 6.64e-19
C1812 net8 _31_/a_285_47# 0.00129f
C1813 net11 _27_/a_27_297# 1.58e-20
C1814 _19_ _01_ 0.031f
C1815 p[13] input3/a_27_47# 0.00527f
C1816 _49_/a_315_47# p[2] 8.45e-20
C1817 input9/a_75_212# input13/a_27_47# 0.00732f
C1818 _06_ _29_/a_111_297# 6.74e-20
C1819 Vin _31_/a_35_297# 3.35e-20
C1820 p[14] p[8] 1.91e-20
C1821 _49_/a_75_199# _35_/a_226_47# 8.73e-20
C1822 _01_ net5 0.0779f
C1823 input8/a_27_47# _02_ 5.08e-20
C1824 th14_0/m1_891_419# p[7] 0.049f
C1825 _09_ _45_/a_27_47# 0.00823f
C1826 input1/a_75_212# th11_0/m1_705_187# 5.25e-20
C1827 _04_ _19_ 0.356f
C1828 _34_/a_47_47# _21_ 8.93e-19
C1829 th11_0/m1_705_187# th11_0/m1_577_n654# -1.6e-19
C1830 net13 _02_ 0.00154f
C1831 p[1] net14 0.0025f
C1832 _12_ _39_/a_47_47# 0.0317f
C1833 _17_ _16_ 0.242f
C1834 p[7] _37_/a_197_47# -3.27e-19
C1835 input5/a_62_47# net3 0.00164f
C1836 _04_ net5 0.00476f
C1837 _20_ _35_/a_76_199# 3.21e-20
C1838 VGND net6 0.512f
C1839 _49_/a_315_47# p[7] 3.4e-19
C1840 th15_0/Vin net2 0.0484f
C1841 VGND _13_ 0.363f
C1842 _10_ _43_/a_27_47# 0.0279f
C1843 th15_0/Vin _44_/a_256_47# 1.36e-19
C1844 _43_/a_27_47# _55_/a_80_21# 1.56e-19
C1845 _34_/a_285_47# net12 8.07e-20
C1846 b[1] _01_ 0.00233f
C1847 _30_/a_215_297# _33_/a_109_93# 0.00104f
C1848 p[14] _37_/a_27_47# 3.97e-19
C1849 th01_0/m1_991_n1219# th11_0/m1_705_187# 7.73e-20
C1850 _12_ net10 7.82e-20
C1851 net7 input5/a_381_47# 4.91e-19
C1852 net13 _30_/a_109_53# 1.05e-19
C1853 _52_/a_93_21# _04_ 2.35e-19
C1854 _14_ net14 0.184f
C1855 _15_ _01_ 0.007f
C1856 VGND input5/a_664_47# 0.0136f
C1857 _04_ b[1] 0.0568f
C1858 p[7] _29_/a_111_297# -5.85e-19
C1859 p[12] _02_ 8.05e-19
C1860 net6 _47_/a_81_21# 2.14e-19
C1861 net4 _47_/a_299_297# 3.28e-19
C1862 _06_ _40_/a_297_297# 1.64e-19
C1863 p[2] input9/a_75_212# 5.13e-20
C1864 p[1] th02_0/m1_571_144# 1.08e-20
C1865 _37_/a_303_47# net15 0.00118f
C1866 p[7] net17 0.037f
C1867 _15_ _04_ 3.61e-20
C1868 VGND _50_/a_429_93# 4.71e-19
C1869 th14_0/m1_641_n318# net15 4.16e-20
C1870 _27_/a_27_297# _27_/a_109_297# -3.68e-20
C1871 _23_ net13 4.11e-19
C1872 _41_/a_59_75# _17_ 0.00149f
C1873 _52_/a_250_297# _18_ 1.77e-19
C1874 net2 input5/a_558_47# 5.99e-21
C1875 _12_ _38_/a_197_47# 0.00173f
C1876 _45_/a_27_47# _39_/a_47_47# 1.31e-19
C1877 _06_ _53_/a_183_297# 0.00146f
C1878 net1 _19_ 2.86e-19
C1879 th15_0/Vin _02_ 7.82e-21
C1880 input15/a_27_47# p[12] 3.73e-19
C1881 _29_/a_29_53# _35_/a_76_199# 9.88e-19
C1882 net9 _33_/a_109_93# 0.00211f
C1883 _39_/a_129_47# _00_ 1.63e-20
C1884 net1 net5 0.0772f
C1885 _43_/a_193_413# net2 1.52e-19
C1886 net11 _35_/a_76_199# 4e-19
C1887 p[8] th09_0/m1_485_n505# 0.00223f
C1888 VGND _42_/a_109_93# -0.0045f
C1889 p[2] input7/a_27_47# 0.0023f
C1890 _22_ _17_ 0.00334f
C1891 input5/a_841_47# _16_ 8.62e-19
C1892 _14_ _18_ 0.243f
C1893 _10_ _44_/a_346_47# 9.13e-21
C1894 net18 _38_/a_27_47# 0.00997f
C1895 _17_ _11_ 0.197f
C1896 p[7] input9/a_75_212# 0.0822f
C1897 _07_ _35_/a_489_413# 0.00429f
C1898 th15_0/Vin input15/a_27_47# 0.00696f
C1899 _03_ _30_/a_297_297# 0.00117f
C1900 _24_ _26_/a_29_53# 2.11e-20
C1901 _14_ _26_/a_29_53# 3.67e-19
C1902 _11_ _40_/a_109_297# 0.00522f
C1903 input14/a_27_47# p[8] 0.0132f
C1904 _40_/a_297_297# p[7] -5.42e-19
C1905 _08_ net11 8.83e-19
C1906 net1 b[1] 0.0593f
C1907 _49_/a_75_199# _01_ 0.009f
C1908 _12_ net15 8.14e-21
C1909 th15_0/Vin th10_0/m1_536_174# 0.0771f
C1910 _14_ _43_/a_469_47# 0.00259f
C1911 _07_ _09_ 0.0416f
C1912 _50_/a_223_47# _03_ 1.41e-21
C1913 _33_/a_109_93# _05_ 0.0206f
C1914 p[7] input7/a_27_47# 0.0772f
C1915 net18 _26_/a_29_53# 2.57e-21
C1916 _37_/a_27_47# net5 1.13e-20
C1917 _20_ net14 8.01e-20
C1918 _49_/a_75_199# _04_ 0.0782f
C1919 _27_/a_27_297# _42_/a_209_311# 4.7e-20
C1920 net6 net16 8.27e-20
C1921 _43_/a_193_413# _02_ 9.4e-21
C1922 VGND p[1] 0.197f
C1923 p[0] input5/a_62_47# 1.39e-19
C1924 _13_ net16 0.0198f
C1925 VGND _52_/a_250_297# -0.00314f
C1926 _44_/a_93_21# input6/a_27_47# 8.53e-19
C1927 _55_/a_217_297# _02_ 6.01e-19
C1928 _42_/a_109_93# output17/a_27_47# 8.6e-21
C1929 p[7] _35_/a_556_47# -6.9e-19
C1930 _47_/a_299_297# net5 0.00198f
C1931 net6 _21_ 2.92e-20
C1932 _13_ _21_ 1.69e-19
C1933 p[11] net14 4.35e-19
C1934 th11_0/m1_705_187# p[13] 0.0061f
C1935 net2 _16_ 0.00654f
C1936 th03_0/m1_890_n844# _31_/a_285_297# 3.4e-20
C1937 VGND _24_ -0.00863f
C1938 net13 net3 3.25e-21
C1939 VGND _14_ 0.226f
C1940 _33_/a_296_53# b[1] 2.69e-20
C1941 _19_ p[10] 9.65e-20
C1942 _43_/a_193_413# input15/a_27_47# 1.62e-20
C1943 _05_ _31_/a_285_47# 5.61e-19
C1944 _34_/a_47_47# _04_ 1.17e-20
C1945 net7 input5/a_841_47# 0.00193f
C1946 _10_ _35_/a_76_199# 7.19e-20
C1947 _13_ _35_/a_226_47# 5.62e-21
C1948 input5/a_664_47# _21_ 9.42e-22
C1949 net5 p[10] 5.12e-21
C1950 _15_ _37_/a_27_47# 1.11e-19
C1951 VGND input12/a_27_47# 0.0405f
C1952 _32_/a_27_47# _50_/a_343_93# 6.48e-20
C1953 VGND net18 0.255f
C1954 _20_ _18_ 0.0151f
C1955 net6 p[9] 0.139f
C1956 th12_0/m1_394_n856# Vin 8.07e-19
C1957 net8 net14 0.0516f
C1958 input6/a_27_47# net15 0.00115f
C1959 _12_ _47_/a_384_47# 9.51e-20
C1960 _09_ net4 0.00262f
C1961 _10_ _08_ 1.51e-19
C1962 _29_/a_29_53# net14 1.61e-20
C1963 _14_ _47_/a_81_21# 6.24e-20
C1964 _15_ _47_/a_299_297# 0.0103f
C1965 net6 net19 0.00346f
C1966 Vin p[12] 0.0619f
C1967 _20_ _26_/a_29_53# 0.00447f
C1968 _49_/a_75_199# net1 0.00799f
C1969 b[1] p[10] 0.114f
C1970 p[11] _18_ 1.24e-19
C1971 net11 net14 9.95e-19
C1972 p[13] net15 0.00241f
C1973 _50_/a_223_47# _00_ 0.00738f
C1974 _50_/a_223_47# _36_/a_27_47# 1.27e-20
C1975 net2 input2/a_27_47# 0.024f
C1976 _07_ net10 0.0605f
C1977 _49_/a_544_297# p[7] 0.00504f
C1978 _02_ _16_ 0.00564f
C1979 _50_/a_27_47# _38_/a_27_47# 2.37e-20
C1980 VGND _45_/a_193_297# -0.00241f
C1981 _12_ _03_ 2.76e-20
C1982 th15_0/Vin net3 0.00715f
C1983 input5/a_664_47# net19 1.38e-21
C1984 th15_0/Vin Vin 0.999f
C1985 _06_ b[2] 0.0116f
C1986 net7 _31_/a_285_297# 0.00227f
C1987 _17_ th12_0/m1_529_n42# 1.35e-20
C1988 net6 output16/a_27_47# 1.5e-19
C1989 _22_ net2 1.93e-20
C1990 _13_ output16/a_27_47# 4.58e-19
C1991 _50_/a_27_47# _18_ 0.0665f
C1992 _16_ _28_/a_109_297# 1.26e-19
C1993 _48_/a_27_47# _02_ 0.00435f
C1994 net11 _38_/a_27_47# 1.68e-20
C1995 net7 net2 0.00234f
C1996 net2 _11_ 0.234f
C1997 VGND _32_/a_303_47# -4.83e-19
C1998 output18/a_27_47# b[2] 0.0141f
C1999 _32_/a_27_47# net5 0.0961f
C2000 _08_ net9 7.71e-21
C2001 input15/a_27_47# _16_ 7.13e-19
C2002 _55_/a_472_297# _15_ 0.00626f
C2003 _52_/a_584_47# _22_ 6.24e-19
C2004 _18_ net8 1.15e-21
C2005 _50_/a_27_47# _26_/a_29_53# 5.56e-19
C2006 p[7] _39_/a_129_47# -9.47e-19
C2007 input3/a_27_47# input14/a_27_47# 5.08e-20
C2008 VGND _20_ 0.471f
C2009 _29_/a_29_53# _26_/a_29_53# 0.00121f
C2010 _35_/a_76_199# _05_ 0.00238f
C2011 _52_/a_346_47# _02_ 0.00526f
C2012 _32_/a_27_47# b[1] 6.39e-19
C2013 net4 _39_/a_47_47# 0.0202f
C2014 _06_ _36_/a_109_47# 0.00168f
C2015 net11 _26_/a_29_53# 1.08e-20
C2016 VGND _34_/a_377_297# -0.00102f
C2017 _42_/a_368_53# b[1] 5.32e-20
C2018 net3 input5/a_558_47# 0.0137f
C2019 _42_/a_109_93# net19 0.0448f
C2020 input7/a_27_47# net17 4.99e-20
C2021 _45_/a_27_47# _03_ 2.06e-20
C2022 input3/a_27_47# b[1] 2.97e-19
C2023 VGND p[11] 0.224f
C2024 p[7] b[2] 0.262f
C2025 _24_ net16 6.93e-19
C2026 net4 net10 8.28e-22
C2027 th15_0/Vin _40_/a_191_297# 3.41e-19
C2028 _09_ _19_ 4.8e-21
C2029 _32_/a_27_47# _15_ 1.19e-19
C2030 _22_ _02_ 0.552f
C2031 _08_ _05_ 0.00897f
C2032 input2/a_27_47# _30_/a_109_53# 1.54e-20
C2033 net14 _27_/a_109_297# 1.32e-19
C2034 net3 _27_/a_205_297# 4.37e-19
C2035 _41_/a_59_75# input15/a_27_47# 3.96e-20
C2036 _43_/a_193_413# net3 5.65e-20
C2037 Vin _27_/a_205_297# 2.93e-20
C2038 _11_ _02_ 0.0621f
C2039 _10_ net14 2.4e-19
C2040 _52_/a_250_297# _35_/a_226_47# 2.63e-20
C2041 net7 _02_ 0.445f
C2042 _55_/a_80_21# net14 4.7e-19
C2043 _55_/a_217_297# net3 5.78e-20
C2044 _15_ input3/a_27_47# 7.53e-19
C2045 _47_/a_81_21# _20_ 0.0457f
C2046 _09_ net5 5.18e-19
C2047 _54_/a_75_212# net18 0.0143f
C2048 _24_ _21_ 0.0388f
C2049 _35_/a_489_413# b[1] 0.00104f
C2050 net13 _33_/a_109_93# 0.0254f
C2051 th15_0/Vin _43_/a_369_47# 1.11e-19
C2052 _12_ _00_ 0.00396f
C2053 _12_ _36_/a_27_47# 0.00178f
C2054 net18 net16 0.00585f
C2055 _49_/a_208_47# _02_ 0.00193f
C2056 VGND _50_/a_27_47# -0.00432f
C2057 p[14] _44_/a_93_21# 2.07e-19
C2058 _11_ _28_/a_109_297# 6.29e-19
C2059 _22_ _30_/a_109_53# 3.67e-21
C2060 net6 _04_ 2.61e-20
C2061 b[1] th02_0/m1_983_133# 7.26e-20
C2062 _04_ _13_ 1.17e-21
C2063 _12_ _35_/a_226_297# 3.35e-20
C2064 _06_ _50_/a_223_47# 0.0481f
C2065 _52_/a_93_21# _09_ 0.0227f
C2066 input15/a_27_47# _11_ 4.4e-19
C2067 _17_ _40_/a_109_297# 9.67e-19
C2068 input12/a_27_47# _21_ 2.32e-19
C2069 VGND net8 0.405f
C2070 net4 _38_/a_197_47# 7.64e-19
C2071 VGND _29_/a_29_53# 0.0544f
C2072 _10_ _38_/a_27_47# 0.0133f
C2073 th03_0/m1_638_n591# p[7] 0.0124f
C2074 net18 _21_ 0.00215f
C2075 p[7] _36_/a_109_47# -4.66e-19
C2076 _09_ b[1] 0.00408f
C2077 VGND net11 0.475f
C2078 net12 _02_ 2.28e-19
C2079 _14_ p[9] 2.62e-21
C2080 net9 net14 7.12e-20
C2081 _50_/a_515_93# net14 1.39e-20
C2082 _45_/a_193_297# net16 0.00187f
C2083 input5/a_664_47# _04_ 6.73e-21
C2084 _22_ _23_ 0.0187f
C2085 _43_/a_297_47# _17_ 5.72e-20
C2086 _10_ _18_ 0.133f
C2087 _23_ _11_ 2e-20
C2088 _14_ net19 0.00714f
C2089 net11 _33_/a_209_311# 2.49e-19
C2090 _55_/a_80_21# _18_ 1.44e-20
C2091 p[0] th15_0/Vin 0.336f
C2092 th15_0/Vin _43_/a_27_47# 1.9e-19
C2093 _10_ _26_/a_111_297# 7.13e-20
C2094 p[7] _30_/a_297_297# -4.92e-19
C2095 _47_/a_81_21# net8 2.08e-21
C2096 _10_ _26_/a_29_53# 0.0265f
C2097 net12 _30_/a_109_53# 4.25e-20
C2098 p[14] net15 0.00328f
C2099 _45_/a_27_47# _00_ 4.84e-20
C2100 _42_/a_209_311# net14 0.0238f
C2101 _42_/a_296_53# net3 1.81e-19
C2102 _16_ net3 1.77e-19
C2103 Vin _16_ 6.65e-20
C2104 _09_ _25_ 1.49e-19
C2105 _10_ b[3] 6.63e-21
C2106 _39_/a_47_47# net5 0.0389f
C2107 _45_/a_193_297# _35_/a_226_47# 8.15e-21
C2108 _43_/a_193_413# _43_/a_369_47# -1.25e-19
C2109 net4 net15 8.68e-19
C2110 net2 th12_0/m1_529_n42# 0.0122f
C2111 p[7] _50_/a_223_47# -0.00601f
C2112 _10_ _43_/a_469_47# 0.00124f
C2113 _38_/a_27_47# _53_/a_29_53# 1.29e-19
C2114 Vin th03_0/m1_890_n844# 2.47e-19
C2115 _49_/a_201_297# net14 1.52e-19
C2116 net8 output17/a_27_47# 0.0043f
C2117 net12 _23_ 2.28e-21
C2118 net10 net5 0.0316f
C2119 _04_ _42_/a_109_93# 5.77e-22
C2120 net9 _18_ 1.51e-19
C2121 input5/a_381_47# net2 0.0138f
C2122 _52_/a_93_21# _39_/a_47_47# 1.44e-20
C2123 _34_/a_285_47# _02_ 7.14e-19
C2124 VGND _30_/a_465_297# 6.42e-19
C2125 _20_ _21_ 0.191f
C2126 net9 _26_/a_29_53# 0.00343f
C2127 net6 p[8] 1.3e-20
C2128 _07_ _03_ 0.0113f
C2129 input5/a_664_47# net1 2.41e-19
C2130 _34_/a_377_297# _21_ 2.37e-19
C2131 VGND _30_/a_215_297# 0.00687f
C2132 _52_/a_93_21# net10 7.84e-20
C2133 p[7] input1/a_75_212# 0.0788f
C2134 p[7] th11_0/m1_577_n654# -4.9e-19
C2135 VGND _27_/a_109_297# -6.15e-19
C2136 _18_ _42_/a_209_311# 3.21e-19
C2137 net10 b[1] 0.117f
C2138 _12_ _39_/a_377_297# 6.77e-19
C2139 p[7] _37_/a_303_47# -3.13e-19
C2140 input5/a_62_47# net14 5.28e-20
C2141 Vin input2/a_27_47# 0.00133f
C2142 _20_ _35_/a_226_47# 5.19e-20
C2143 VGND _10_ 1.15f
C2144 p[7] th14_0/m1_641_n318# 0.00238f
C2145 _09_ _49_/a_75_199# 2.93e-19
C2146 _06_ _12_ 0.136f
C2147 th15_0/Vin _44_/a_346_47# 1.88e-19
C2148 VGND _55_/a_80_21# 0.00281f
C2149 _43_/a_27_47# _55_/a_217_297# 2.18e-19
C2150 _44_/a_93_21# net5 3.61e-20
C2151 _30_/a_215_297# _33_/a_209_311# 1.56e-19
C2152 th01_0/m1_991_n1219# p[7] 0.0681f
C2153 _50_/a_27_47# net16 2.35e-20
C2154 net6 _37_/a_27_47# 4.3e-20
C2155 _04_ p[1] 9.99e-21
C2156 _52_/a_250_297# _04_ 3.98e-21
C2157 VGND th13_0/m1_831_275# 0.0456f
C2158 _14_ _01_ 0.0193f
C2159 _22_ net3 9.39e-20
C2160 _35_/a_76_199# net13 0.0337f
C2161 _54_/a_75_212# net11 0.00956f
C2162 _11_ net3 0.165f
C2163 _27_/a_27_297# input5/a_558_47# 1.57e-19
C2164 net7 net3 7.45e-20
C2165 Vin _11_ 1.06e-19
C2166 _20_ net19 1.29e-19
C2167 net7 Vin 0.00115f
C2168 _50_/a_27_47# _21_ 3.38e-21
C2169 _34_/a_129_47# _08_ 3.29e-19
C2170 p[11] p[9] 0.00354f
C2171 net6 _47_/a_299_297# 3.63e-19
C2172 net11 net16 4.43e-22
C2173 _10_ _47_/a_81_21# 0.0061f
C2174 net2 _17_ 0.181f
C2175 _25_ net10 2.66e-19
C2176 th11_0/m1_705_187# b[1] 0.00504f
C2177 net8 _21_ 0.00656f
C2178 _29_/a_29_53# _21_ 0.0775f
C2179 VGND _50_/a_515_93# -4.75e-19
C2180 _14_ _04_ 2.04e-21
C2181 VGND net9 0.372f
C2182 p[11] net19 0.00647f
C2183 _19_ net15 0.00628f
C2184 net2 _40_/a_109_297# 0.0011f
C2185 _08_ net13 1.82e-19
C2186 _12_ _38_/a_303_47# 0.00153f
C2187 net11 _21_ 0.586f
C2188 _15_ _44_/a_93_21# 0.0168f
C2189 VGND _53_/a_29_53# -0.0168f
C2190 _12_ p[7] 0.28f
C2191 _06_ _45_/a_27_47# 0.0021f
C2192 net5 net15 0.0226f
C2193 input11/a_27_47# net11 0.00318f
C2194 _29_/a_29_53# _35_/a_226_47# 2.64e-19
C2195 net9 _33_/a_209_311# 4.33e-20
C2196 Vin th15_0/m1_597_n912# 7.85e-19
C2197 _39_/a_285_47# _00_ 1.47e-21
C2198 input4/a_75_212# _18_ 4.36e-19
C2199 _12_ th15_0/m1_849_n157# 2.47e-21
C2200 net11 _35_/a_226_47# 3.21e-19
C2201 _53_/a_111_297# _24_ 9.08e-21
C2202 _06_ _36_/a_303_47# 5.3e-19
C2203 VGND _42_/a_209_311# -0.008f
C2204 _10_ _44_/a_584_47# 1.14e-20
C2205 _43_/a_27_47# _16_ 2.47e-19
C2206 th14_0/m1_891_419# th11_0/m1_577_n654# 0.0383f
C2207 _26_/a_183_297# _14_ 6.98e-22
C2208 net9 _47_/a_81_21# 3.49e-19
C2209 _06_ input6/a_27_47# 2.85e-19
C2210 net19 net8 1.15e-19
C2211 b[1] net15 0.00314f
C2212 VGND _49_/a_201_297# -0.00403f
C2213 _11_ _40_/a_191_297# 0.00207f
C2214 net1 p[1] 0.0291f
C2215 _42_/a_109_93# _37_/a_27_47# 2.55e-20
C2216 _17_ _02_ 0.00482f
C2217 VGND _05_ 0.754f
C2218 _32_/a_303_47# _01_ 8.58e-19
C2219 VGND _31_/a_35_297# -0.00828f
C2220 _15_ net15 0.156f
C2221 _33_/a_209_311# _05_ 0.0311f
C2222 input6/a_27_47# output19/a_27_47# 0.107f
C2223 _45_/a_27_47# p[7] -0.00418f
C2224 input15/a_27_47# _17_ 6.14e-19
C2225 _20_ _01_ 0.161f
C2226 _27_/a_27_297# _16_ 3.74e-22
C2227 _34_/a_47_47# net10 0.0507f
C2228 _10_ net16 0.0338f
C2229 VGND _52_/a_256_47# -0.00161f
C2230 VGND input5/a_62_47# 0.0499f
C2231 p[7] _36_/a_303_47# -4.83e-19
C2232 _30_/a_215_297# _21_ 1.48e-19
C2233 _42_/a_109_93# p[10] 1.82e-21
C2234 input12/a_27_47# net1 7.44e-20
C2235 p[7] input6/a_27_47# 0.00129f
C2236 _47_/a_384_47# net5 0.00129f
C2237 p[13] _44_/a_250_297# 4.09e-20
C2238 _10_ _21_ 0.00421f
C2239 VGND input4/a_75_212# 0.0528f
C2240 _20_ _04_ 0.0677f
C2241 _32_/a_109_47# net8 0.0011f
C2242 th13_0/m1_831_275# net16 1.81e-20
C2243 net4 _00_ 0.0166f
C2244 net13 net14 2.21e-21
C2245 net4 _36_/a_27_47# 0.0103f
C2246 p[7] p[13] 0.318f
C2247 _33_/a_368_53# b[1] 4.19e-19
C2248 _22_ _43_/a_27_47# 0.091f
C2249 _19_ _03_ 0.0019f
C2250 _34_/a_377_297# _04_ 1.7e-20
C2251 _43_/a_27_47# _11_ 4.27e-19
C2252 VGND input10/a_27_47# 0.00285f
C2253 p[0] net7 1.36e-19
C2254 _05_ output17/a_27_47# 1.12e-19
C2255 net7 _43_/a_27_47# 6.31e-19
C2256 _10_ _35_/a_226_47# 1.25e-19
C2257 _03_ net5 1.04e-19
C2258 net3 th12_0/m1_529_n42# 3.65e-21
C2259 Vin th12_0/m1_529_n42# 0.0341f
C2260 _14_ _37_/a_27_47# 0.00137f
C2261 _22_ _33_/a_109_93# 1.34e-22
C2262 input5/a_841_47# _02_ 0.00591f
C2263 _27_/a_27_297# input2/a_27_47# 1.16e-19
C2264 _10_ p[9] 0.00225f
C2265 _53_/a_29_53# net16 2.04e-20
C2266 input5/a_381_47# net3 0.0299f
C2267 _06_ _39_/a_285_47# 1.23e-20
C2268 net8 _01_ 0.0802f
C2269 _09_ net6 5.43e-20
C2270 _49_/a_75_199# net15 5.13e-20
C2271 p[1] p[10] 9.56e-19
C2272 _09_ _13_ 0.0927f
C2273 _15_ _47_/a_384_47# 0.00112f
C2274 net9 _21_ 0.0282f
C2275 _29_/a_29_53# _01_ 8.33e-20
C2276 _29_/a_183_297# net3 7.38e-21
C2277 _06_ _07_ 0.185f
C2278 _52_/a_93_21# _03_ 0.00985f
C2279 input5/a_62_47# output17/a_27_47# 1.02e-19
C2280 _10_ net19 3.43e-19
C2281 _55_/a_80_21# net19 0.00423f
C2282 _32_/a_303_47# net1 1.45e-19
C2283 net11 _01_ 3.82e-20
C2284 _04_ _50_/a_27_47# 2.07e-21
C2285 _50_/a_343_93# _00_ 0.102f
C2286 _03_ b[1] 0.0738f
C2287 _53_/a_29_53# _21_ 0.00959f
C2288 _18_ net13 1.06e-20
C2289 net9 _35_/a_226_47# 1.22e-20
C2290 net7 _27_/a_27_297# 1.22e-19
C2291 VGND _45_/a_205_47# -2.47e-19
C2292 _04_ net8 0.02f
C2293 input3/a_27_47# _42_/a_109_93# 0.00249f
C2294 _04_ _29_/a_29_53# 0.0408f
C2295 input1/a_75_212# input7/a_27_47# 3.2e-20
C2296 th15_0/Vin net14 0.0111f
C2297 _15_ _03_ 7.39e-20
C2298 net12 _33_/a_109_93# 0.0435f
C2299 _55_/a_300_47# b[1] 1.1e-19
C2300 net7 _31_/a_285_47# 0.00132f
C2301 net13 _26_/a_29_53# 2.23e-20
C2302 net1 _20_ 0.363f
C2303 net11 _04_ 0.078f
C2304 _02_ _31_/a_285_297# 5.86e-20
C2305 _55_/a_472_297# _14_ 0.00192f
C2306 _55_/a_300_47# _15_ 1.42e-20
C2307 _05_ _21_ 0.0104f
C2308 th14_0/m1_891_419# p[13] 0.0575f
C2309 _25_ _03_ 0.00422f
C2310 p[7] _39_/a_285_47# -9.53e-19
C2311 p[12] _18_ 2.17e-19
C2312 th13_0/m1_831_275# output16/a_27_47# 7.67e-22
C2313 _07_ p[7] 0.0761f
C2314 p[14] _41_/a_145_75# 1.12e-19
C2315 _17_ net3 0.0698f
C2316 _35_/a_226_47# _49_/a_201_297# 1.66e-20
C2317 Vin _17_ 3.65e-19
C2318 _42_/a_209_311# p[9] 5.51e-21
C2319 net5 _00_ 0.00954f
C2320 _35_/a_226_47# _05_ 0.0134f
C2321 VGND _36_/a_197_47# -3.75e-19
C2322 _06_ p[14] 2.49e-19
C2323 _36_/a_27_47# net5 0.0163f
C2324 _52_/a_584_47# _02_ 0.00389f
C2325 p[11] p[8] 0.00322f
C2326 th15_0/Vin th02_0/m1_571_144# 8.16e-21
C2327 VGND input8/a_27_47# 0.0574f
C2328 net4 _39_/a_377_297# 8.88e-19
C2329 net6 _39_/a_47_47# 0.0249f
C2330 _40_/a_109_297# net3 3.14e-19
C2331 VGND _34_/a_129_47# -8.76e-20
C2332 _13_ _39_/a_47_47# 0.00117f
C2333 net14 input5/a_558_47# 0.0325f
C2334 _42_/a_209_311# net19 0.0766f
C2335 _06_ net4 0.281f
C2336 th15_0/Vin _18_ 6.4e-19
C2337 net2 input15/a_27_47# 0.00296f
C2338 _54_/a_75_212# input10/a_27_47# 1.17e-22
C2339 net6 net10 1.35e-20
C2340 net1 net8 0.381f
C2341 _13_ net10 4.52e-21
C2342 VGND net13 0.142f
C2343 net1 _29_/a_29_53# 9.76e-19
C2344 _43_/a_193_413# net14 1.11e-19
C2345 net3 _27_/a_277_297# 2.71e-19
C2346 net14 _27_/a_205_297# 3.63e-19
C2347 _08_ _48_/a_27_47# 2.58e-19
C2348 Vin _27_/a_277_297# 1.98e-20
C2349 _36_/a_27_47# b[1] 7.95e-19
C2350 _10_ _01_ 2.22e-19
C2351 net11 net1 1.13e-19
C2352 p[14] output19/a_27_47# 0.0459f
C2353 _55_/a_80_21# _01_ 0.0121f
C2354 _55_/a_217_297# net14 2.1e-19
C2355 _47_/a_299_297# _20_ 0.002f
C2356 _49_/a_75_199# _03_ 0.0849f
C2357 net9 _32_/a_109_47# 6.44e-19
C2358 _35_/a_226_297# b[1] 1.03e-19
C2359 th15_0/Vin b[3] 0.106f
C2360 net13 _33_/a_209_311# 0.0227f
C2361 _04_ _30_/a_215_297# 0.00225f
C2362 th15_0/Vin _43_/a_469_47# 2.09e-19
C2363 p[1] th02_0/m1_983_133# 0.122f
C2364 _15_ _00_ 0.207f
C2365 p[13] net17 8.11e-20
C2366 p[14] _44_/a_250_297# 7.34e-21
C2367 _04_ _27_/a_109_297# 7.2e-20
C2368 input11/a_27_47# input10/a_27_47# 5.3e-19
C2369 _10_ _04_ 9.24e-20
C2370 _22_ _35_/a_76_199# 6.58e-21
C2371 _06_ _50_/a_343_93# 0.0376f
C2372 VGND th12_0/m1_394_n856# 0.0134f
C2373 p[7] p[14] 0.0553f
C2374 _17_ _40_/a_191_297# 4.35e-19
C2375 _52_/a_250_297# _09_ 1.97e-20
C2376 net6 _44_/a_93_21# 1.08e-20
C2377 net4 _38_/a_303_47# 5.95e-19
C2378 _35_/a_76_199# _11_ 6.99e-22
C2379 net7 _35_/a_76_199# 1.79e-20
C2380 _10_ _38_/a_109_47# 5.44e-19
C2381 VGND p[12] 0.359f
C2382 net4 p[7] 1.07f
C2383 th15_0/m1_849_n157# p[14] 0.0846f
C2384 _34_/a_47_47# _03_ 4.5e-20
C2385 _02_ _30_/a_109_53# 5.03e-22
C2386 _25_ _36_/a_27_47# 2.34e-20
C2387 _50_/a_615_93# net14 1.69e-20
C2388 net9 _01_ 0.157f
C2389 p[11] p[10] 0.00389f
C2390 net8 _37_/a_27_47# 6.66e-21
C2391 _09_ _24_ 0.0202f
C2392 _43_/a_193_413# _18_ 0.0413f
C2393 _43_/a_369_47# _17_ 5.87e-19
C2394 _55_/a_472_297# _20_ 0.00212f
C2395 _10_ _53_/a_111_297# 2.06e-19
C2396 input5/a_664_47# _44_/a_93_21# 1.88e-20
C2397 VGND th15_0/Vin 1.04f
C2398 _08_ net7 9.54e-25
C2399 input13/a_27_47# b[1] 0.00624f
C2400 _10_ _26_/a_183_297# 5.74e-19
C2401 _23_ _02_ 0.0648f
C2402 net9 _04_ 0.0213f
C2403 _45_/a_109_297# _00_ 4.86e-20
C2404 net12 _35_/a_76_199# 0.0132f
C2405 _16_ net14 0.00266f
C2406 _42_/a_209_311# _01_ 1.58e-19
C2407 _42_/a_296_53# net14 2.18e-19
C2408 _09_ net18 1.97e-21
C2409 input5/a_381_47# _27_/a_27_297# 1.47e-19
C2410 _39_/a_377_297# net5 0.00234f
C2411 net1 _30_/a_215_297# 0.00375f
C2412 net6 net15 0.0664f
C2413 _06_ net5 0.41f
C2414 p[7] _50_/a_343_93# -0.0126f
C2415 net8 p[10] 0.00619f
C2416 _49_/a_201_297# _01_ 0.0105f
C2417 p[2] _19_ 1.1e-21
C2418 _10_ net1 4.34e-19
C2419 th15_0/Vin _47_/a_81_21# 6.76e-20
C2420 _32_/a_27_47# _20_ 0.0069f
C2421 _05_ _01_ 5.03e-19
C2422 _50_/a_343_93# th15_0/m1_849_n157# 2.76e-21
C2423 _43_/a_27_47# _17_ 0.00131f
C2424 net1 _55_/a_80_21# 1.8e-19
C2425 th15_0/Vin th10_0/m1_502_n495# 0.0036f
C2426 _04_ _42_/a_209_311# 9.84e-22
C2427 _08_ net12 0.0269f
C2428 Vin _31_/a_285_297# 7.71e-20
C2429 _01_ _31_/a_35_297# 4.27e-19
C2430 _42_/a_109_93# _44_/a_93_21# 1.25e-19
C2431 _09_ _45_/a_193_297# 0.00961f
C2432 input5/a_664_47# net15 0.0216f
C2433 VGND input5/a_558_47# -0.00104f
C2434 _52_/a_93_21# _06_ 0.0584f
C2435 _04_ _49_/a_201_297# 0.0253f
C2436 net2 net3 0.519f
C2437 _06_ b[1] 0.0885f
C2438 net2 Vin 0.0131f
C2439 Vin th09_0/m1_962_372# 0.00142f
C2440 _44_/a_256_47# net3 0.00101f
C2441 _04_ _05_ 0.0352f
C2442 _52_/a_250_297# net10 2.86e-21
C2443 input14/a_27_47# output19/a_27_47# 0.0101f
C2444 th15_0/Vin output17/a_27_47# 1.87e-20
C2445 p[11] input3/a_27_47# 0.0153f
C2446 _04_ _31_/a_35_297# 1.89e-20
C2447 VGND _27_/a_205_297# -3.36e-19
C2448 input2/a_27_47# net14 0.0102f
C2449 p[7] th09_0/m1_485_n505# 0.0937f
C2450 _12_ _39_/a_129_47# 0.00175f
C2451 VGND _43_/a_193_413# -0.0147f
C2452 _18_ _16_ 0.144f
C2453 output18/a_27_47# b[1] 9.26e-19
C2454 p[7] _19_ 0.0335f
C2455 _06_ _15_ 0.22f
C2456 th15_0/Vin _44_/a_584_47# 2.71e-19
C2457 VGND _55_/a_217_297# -0.00342f
C2458 th03_0/m1_890_n844# th02_0/m1_571_144# 1.09e-20
C2459 net13 _21_ 0.13f
C2460 _44_/a_250_297# net5 3.11e-20
C2461 p[2] b[1] 0.00237f
C2462 p[14] _37_/a_197_47# 1.52e-19
C2463 input14/a_27_47# _44_/a_250_297# 8.25e-21
C2464 net9 net1 0.47f
C2465 p[12] th13_0/m1_559_n458# 2.29e-19
C2466 _17_ _27_/a_27_297# 6.78e-22
C2467 p[7] net5 0.613f
C2468 p[7] input14/a_27_47# 0.0739f
C2469 _04_ input5/a_62_47# 0.00345f
C2470 _22_ net14 2.23e-19
C2471 _09_ _20_ 7.11e-19
C2472 _35_/a_226_47# net13 0.00709f
C2473 _32_/a_27_47# net8 0.0275f
C2474 _11_ net14 5e-19
C2475 th01_0/m1_991_n1219# th03_0/m1_638_n591# 2.42e-20
C2476 _06_ _25_ 0.144f
C2477 net7 net14 2.23e-19
C2478 _42_/a_109_93# net15 4.62e-19
C2479 _12_ b[2] 3.89e-20
C2480 _32_/a_197_47# net5 5.61e-21
C2481 _34_/a_285_47# _08_ 0.00414f
C2482 input12/a_27_47# net10 0.00182f
C2483 th15_0/Vin th13_0/m1_559_n458# 1.16e-21
C2484 _10_ _47_/a_299_297# 0.0134f
C2485 _52_/a_93_21# p[7] -0.00838f
C2486 net18 net10 3.35e-20
C2487 _17_ _44_/a_346_47# 7.2e-19
C2488 _02_ net3 9.52e-20
C2489 _25_ output18/a_27_47# 0.072f
C2490 Vin _02_ 3.16e-21
C2491 p[7] b[1] 1.09f
C2492 VGND _50_/a_615_93# -5.19e-19
C2493 net2 _40_/a_191_297# 0.00143f
C2494 _14_ _44_/a_93_21# 0.04f
C2495 _15_ _44_/a_250_297# 0.00517f
C2496 _22_ _38_/a_27_47# 2.86e-19
C2497 net1 _49_/a_201_297# 0.00304f
C2498 _45_/a_193_297# _39_/a_47_47# 1.4e-20
C2499 _11_ _38_/a_27_47# 0.071f
C2500 net1 _05_ 0.151f
C2501 _06_ _45_/a_109_297# 0.0023f
C2502 _15_ p[7] 0.912f
C2503 net6 _03_ 2.9e-20
C2504 _13_ _03_ 1.74e-20
C2505 net1 _31_/a_35_297# 0.0111f
C2506 input15/a_27_47# net3 8.74e-20
C2507 input15/a_27_47# Vin 0.00251f
C2508 _15_ th15_0/m1_849_n157# 2.53e-19
C2509 _09_ _50_/a_27_47# 1.3e-19
C2510 _22_ _18_ 0.0211f
C2511 VGND _16_ -0.00582f
C2512 th12_0/m1_394_n856# p[9] 1.33e-19
C2513 _18_ _11_ 0.484f
C2514 net7 _18_ 2.58e-20
C2515 _26_/a_111_297# _22_ 0.00137f
C2516 _07_ _35_/a_556_47# 0.00128f
C2517 p[1] net15 1.8e-19
C2518 p[12] p[9] 1.02e-19
C2519 _10_ _55_/a_472_297# 7.35e-21
C2520 _25_ p[7] 0.0829f
C2521 _55_/a_472_297# _55_/a_80_21# 1.78e-33
C2522 VGND _30_/a_392_297# 3.41e-19
C2523 _09_ _29_/a_29_53# 0.00488f
C2524 VGND th03_0/m1_890_n844# 0.0199f
C2525 _22_ _26_/a_29_53# 0.09f
C2526 net1 input5/a_62_47# 7.59e-20
C2527 Vin th10_0/m1_536_174# 0.102f
C2528 _42_/a_209_311# _37_/a_27_47# 1.59e-20
C2529 _11_ _26_/a_29_53# 1.09e-19
C2530 _09_ net11 0.0262f
C2531 VGND _48_/a_27_47# 0.0548f
C2532 VGND _31_/a_117_297# -0.00177f
C2533 _20_ _39_/a_47_47# 2.3e-20
C2534 th14_0/m1_891_419# net5 0.00243f
C2535 _49_/a_75_199# p[2] 2.21e-19
C2536 th11_0/m1_577_n654# th14_0/m1_641_n318# 2.63e-20
C2537 _14_ net15 0.0538f
C2538 th15_0/Vin p[9] 0.228f
C2539 _49_/a_315_47# _19_ 1.33e-19
C2540 _33_/a_296_53# _05_ 4.53e-19
C2541 input5/a_62_47# p[8] 1.22e-19
C2542 _34_/a_47_47# _06_ 0.0391f
C2543 _43_/a_27_47# net2 0.01f
C2544 _20_ net10 3.23e-19
C2545 _45_/a_109_297# p[7] -0.011f
C2546 th15_0/Vin net19 0.00574f
C2547 net12 _18_ 2.25e-21
C2548 _34_/a_377_297# net10 1.62e-19
C2549 VGND _41_/a_59_75# 0.0205f
C2550 VGND input2/a_27_47# -0.0137f
C2551 _12_ _50_/a_223_47# 0.00327f
C2552 VGND _52_/a_346_47# -0.00175f
C2553 _10_ _32_/a_27_47# 0.00217f
C2554 input8/a_27_47# _01_ 1.43e-19
C2555 _42_/a_209_311# p[10] 2.37e-20
C2556 net12 _26_/a_29_53# 6.55e-19
C2557 _49_/a_75_199# p[7] 0.0154f
C2558 net6 _36_/a_27_47# 5.1e-19
C2559 net6 _00_ 0.00178f
C2560 net13 _01_ 0.00228f
C2561 _13_ _00_ 3.77e-20
C2562 VGND _22_ 0.0404f
C2563 _49_/a_315_47# b[1] 5.66e-19
C2564 input8/a_27_47# _04_ 2.36e-22
C2565 _19_ net17 0.0211f
C2566 VGND _11_ 0.091f
C2567 VGND net7 0.421f
C2568 _05_ p[10] 6.39e-20
C2569 _10_ _35_/a_489_413# 3.41e-19
C2570 _41_/a_59_75# _47_/a_81_21# 1.5e-19
C2571 _31_/a_35_297# p[10] 3.66e-19
C2572 net2 _27_/a_27_297# 0.0131f
C2573 _50_/a_27_47# net10 3.78e-21
C2574 net14 th12_0/m1_529_n42# 3.01e-19
C2575 net19 input5/a_558_47# 2.24e-20
C2576 net17 net5 4.21e-21
C2577 _15_ _37_/a_197_47# 3.02e-19
C2578 _43_/a_27_47# _02_ 1.88e-21
C2579 p[11] _44_/a_93_21# 7.91e-19
C2580 net9 _32_/a_27_47# 0.0136f
C2581 _34_/a_47_47# p[7] 0.0389f
C2582 VGND _49_/a_208_47# -0.00164f
C2583 _04_ net13 0.569f
C2584 net8 net10 2.05e-21
C2585 _43_/a_193_413# p[9] 1.09e-19
C2586 _29_/a_29_53# net10 1.77e-19
C2587 input5/a_381_47# net14 0.00479f
C2588 _10_ _09_ 0.0222f
C2589 _43_/a_193_413# net19 3.31e-19
C2590 _22_ _47_/a_81_21# 7.25e-19
C2591 net11 net10 0.592f
C2592 _02_ _33_/a_109_93# 1.54e-21
C2593 net2 _44_/a_346_47# 1.64e-19
C2594 input2/a_27_47# output17/a_27_47# 0.107f
C2595 _47_/a_81_21# _11_ 0.0454f
C2596 VGND th15_0/m1_597_n912# 0.051f
C2597 net17 b[1] 0.0287f
C2598 Vin net3 0.00372f
C2599 VGND net12 0.344f
C2600 VGND _45_/a_465_47# -8.14e-19
C2601 _20_ net15 0.0021f
C2602 input3/a_27_47# _42_/a_209_311# 1.56e-19
C2603 _24_ _03_ 9.46e-20
C2604 net12 _33_/a_209_311# 0.0769f
C2605 _18_ th12_0/m1_529_n42# 1.01e-20
C2606 _27_/a_27_297# _02_ 0.00179f
C2607 th11_0/m1_705_187# net8 0.00167f
C2608 net7 output17/a_27_47# 0.0018f
C2609 _32_/a_27_47# _05_ 2.2e-20
C2610 net1 input8/a_27_47# 0.0347f
C2611 _19_ input7/a_27_47# 3.12e-21
C2612 p[11] net15 1.71e-19
C2613 _32_/a_27_47# _31_/a_35_297# 9.17e-20
C2614 _09_ net9 2.62e-19
C2615 input9/a_75_212# b[1] 0.00598f
C2616 _55_/a_300_47# _14_ 8.09e-19
C2617 net18 _03_ 2.07e-21
C2618 _48_/a_27_47# _21_ 0.0121f
C2619 _09_ _53_/a_29_53# 0.00642f
C2620 net1 net13 3.51e-19
C2621 _17_ net14 0.104f
C2622 input1/a_75_212# p[13] 4.16e-19
C2623 p[13] th11_0/m1_577_n654# 0.029f
C2624 _30_/a_465_297# net10 0.00106f
C2625 _40_/a_191_297# net3 1.89e-19
C2626 net6 _39_/a_377_297# 0.00143f
C2627 VGND _34_/a_285_47# -0.00301f
C2628 _10_ _39_/a_47_47# 0.00824f
C2629 p[13] th14_0/m1_641_n318# 0.00188f
C2630 _01_ input5/a_558_47# 3.97e-20
C2631 input3/a_27_47# input5/a_62_47# 0.00179f
C2632 _42_/a_296_53# net19 2.71e-19
C2633 net19 _16_ 0.206f
C2634 _06_ net6 0.308f
C2635 input7/a_27_47# b[1] 0.00663f
C2636 _06_ _13_ 0.00188f
C2637 _30_/a_215_297# net10 0.0512f
C2638 net8 net15 0.2f
C2639 _45_/a_193_297# _03_ 2.57e-20
C2640 _54_/a_75_212# _11_ 3.22e-20
C2641 _09_ _49_/a_201_297# 1.74e-20
C2642 _22_ net16 0.00606f
C2643 _10_ net10 4.45e-19
C2644 _48_/a_181_47# _02_ 3.9e-19
C2645 _09_ _05_ 0.0683f
C2646 _11_ net16 0.172f
C2647 net14 _27_/a_277_297# 5.1e-19
C2648 _43_/a_193_413# _01_ 8.16e-19
C2649 _43_/a_297_47# net14 1.09e-21
C2650 b[0] Vin 1.65e-19
C2651 _04_ input5/a_558_47# 1.25e-20
C2652 _45_/a_27_47# _12_ 0.0867f
C2653 VGND _48_/a_109_47# 9.44e-19
C2654 _55_/a_217_297# _01_ 0.00112f
C2655 _47_/a_384_47# _20_ 1.72e-19
C2656 _06_ input5/a_664_47# 3.21e-19
C2657 _22_ _21_ 0.00314f
C2658 _49_/a_75_199# net17 0.00127f
C2659 _35_/a_556_47# b[1] 3.23e-19
C2660 VGND th12_0/m1_529_n42# 0.00796f
C2661 net13 _33_/a_296_53# 3.71e-20
C2662 net6 output19/a_27_47# 0.00112f
C2663 th12_0/m1_394_n856# p[8] 0.00768f
C2664 _11_ _21_ 9.98e-20
C2665 net7 _21_ 3e-19
C2666 _14_ _00_ 0.133f
C2667 _17_ _18_ 0.271f
C2668 _41_/a_59_75# p[9] 1.02e-19
C2669 _04_ _27_/a_205_297# 6.42e-19
C2670 _43_/a_193_413# _04_ 5.67e-21
C2671 th15_0/Vin net1 4.02e-19
C2672 _22_ _35_/a_226_47# 1.39e-20
C2673 _06_ _50_/a_429_93# 0.00169f
C2674 VGND input5/a_381_47# -0.00305f
C2675 net19 input2/a_27_47# 2.9e-23
C2676 _41_/a_59_75# net19 1.97e-20
C2677 _20_ _03_ 0.0794f
C2678 VGND _29_/a_183_297# 4.41e-19
C2679 _10_ _38_/a_197_47# 6.29e-19
C2680 _10_ _44_/a_93_21# 2.48e-19
C2681 net7 _35_/a_226_47# 2.93e-20
C2682 net6 p[7] 0.999f
C2683 net9 net10 0.111f
C2684 _34_/a_377_297# _03_ 3.13e-20
C2685 p[7] _13_ 0.0804f
C2686 p[0] Vin 0.134f
C2687 th15_0/Vin p[8] 0.167f
C2688 _17_ b[3] 5.76e-20
C2689 _35_/a_76_199# _02_ 5.73e-19
C2690 net6 th15_0/m1_849_n157# 3.87e-20
C2691 _53_/a_29_53# net10 7.88e-22
C2692 _11_ p[9] 1.01e-19
C2693 _43_/a_469_47# _17_ 0.00177f
C2694 net12 _21_ 0.23f
C2695 _06_ _42_/a_109_93# 5.53e-20
C2696 _22_ net19 2.17e-19
C2697 _11_ net19 2.19e-19
C2698 input5/a_664_47# p[7] 0.00488f
C2699 net1 input5/a_558_47# 1.1e-19
C2700 _49_/a_544_297# b[1] 8.23e-19
C2701 _08_ _02_ 2.26e-20
C2702 _45_/a_193_297# _00_ 4.38e-20
C2703 net12 _35_/a_226_47# 8.29e-19
C2704 _16_ _01_ 3.24e-19
C2705 th15_0/Vin _37_/a_27_47# 0.00332f
C2706 _39_/a_129_47# net5 0.00344f
C2707 _10_ net15 0.0101f
C2708 p[7] _50_/a_429_93# -3.61e-19
C2709 _44_/a_584_47# th12_0/m1_529_n42# 1.38e-20
C2710 _55_/a_80_21# net15 0.00759f
C2711 _05_ net10 0.457f
C2712 _42_/a_109_93# output19/a_27_47# 1.56e-20
C2713 net8 _03_ 0.0287f
C2714 _27_/a_27_297# net3 0.0166f
C2715 input5/a_381_47# output17/a_27_47# 6.6e-20
C2716 Vin _27_/a_27_297# 2.78e-19
C2717 net10 _31_/a_35_297# 3.95e-20
C2718 th15_0/Vin _47_/a_299_297# 8.81e-20
C2719 _29_/a_29_53# _03_ 0.0414f
C2720 VGND _17_ 0.313f
C2721 Vin _31_/a_285_47# 2.61e-20
C2722 net11 _03_ 0.0952f
C2723 net4 _50_/a_223_47# 0.0107f
C2724 VGND _40_/a_109_297# -0.00181f
C2725 _42_/a_209_311# _44_/a_93_21# 2.21e-19
C2726 _42_/a_109_93# _44_/a_250_297# 6.38e-19
C2727 _52_/a_250_297# _06_ 0.0058f
C2728 net2 net14 0.151f
C2729 p[7] _42_/a_109_93# -0.00115f
C2730 b[2] net5 7.33e-20
C2731 _44_/a_256_47# net14 0.00379f
C2732 _44_/a_346_47# net3 8.04e-19
C2733 _20_ _00_ 0.271f
C2734 _34_/a_285_47# _21_ 6.94e-20
C2735 _52_/a_256_47# net10 8.13e-20
C2736 _20_ _36_/a_27_47# 0.00148f
C2737 th15_0/Vin p[10] 0.185f
C2738 input4/a_75_212# _39_/a_47_47# 3.1e-19
C2739 VGND _27_/a_277_297# -4.65e-19
C2740 _08_ _23_ 1.81e-19
C2741 _12_ _39_/a_285_47# 0.0221f
C2742 VGND _43_/a_297_47# -1.33e-19
C2743 p[2] p[1] 0.0489f
C2744 net9 net15 8.49e-20
C2745 _47_/a_81_21# _17_ 0.0456f
C2746 _06_ _24_ 0.113f
C2747 _07_ _12_ 2.94e-23
C2748 _06_ _14_ 0.0556f
C2749 th11_0/m1_705_187# _31_/a_35_297# 9e-21
C2750 _52_/a_93_21# b[2] 1.63e-19
C2751 b[2] b[1] 5.48e-19
C2752 _43_/a_193_413# _37_/a_27_47# 0.0102f
C2753 _04_ input2/a_27_47# 4.5e-21
C2754 input10/a_27_47# net10 0.00321f
C2755 _22_ _01_ 0.15f
C2756 input5/a_664_47# th14_0/m1_891_419# 2.08e-20
C2757 _35_/a_489_413# net13 7.36e-20
C2758 _06_ input12/a_27_47# 5.3e-22
C2759 net7 _01_ 0.233f
C2760 _06_ net18 0.0211f
C2761 _42_/a_209_311# net15 0.0157f
C2762 input5/a_62_47# _44_/a_93_21# 5.05e-20
C2763 _36_/a_109_47# net5 0.00144f
C2764 _14_ output19/a_27_47# 1.43e-19
C2765 p[7] p[1] 0.135f
C2766 _52_/a_250_297# p[7] 0.019f
C2767 net2 _18_ 0.00181f
C2768 _10_ _47_/a_384_47# 3.53e-19
C2769 _50_/a_27_47# _36_/a_27_47# 6.08e-19
C2770 _50_/a_27_47# _00_ 0.00197f
C2771 input5/a_558_47# p[10] 1.09e-19
C2772 _30_/a_465_297# _03_ 7.72e-19
C2773 _02_ net14 0.00952f
C2774 net18 output18/a_27_47# 0.0106f
C2775 VGND input5/a_841_47# 0.0943f
C2776 _49_/a_208_47# _01_ 2.13e-19
C2777 _22_ _04_ 1.76e-20
C2778 _49_/a_201_297# net15 1.41e-19
C2779 net8 _00_ 3.23e-19
C2780 _36_/a_27_47# net8 1.52e-19
C2781 _09_ net13 0.0379f
C2782 net7 _04_ 0.0602f
C2783 _30_/a_215_297# _03_ 0.0393f
C2784 net1 th03_0/m1_890_n844# 2.78e-20
C2785 _14_ _44_/a_250_297# 4.82e-19
C2786 _29_/a_29_53# _36_/a_27_47# 6.92e-20
C2787 _25_ b[2] 0.0015f
C2788 th03_0/m1_638_n591# b[1] 1.59e-19
C2789 th15_0/Vin _42_/a_368_53# 1.2e-20
C2790 _06_ _45_/a_193_297# 0.00201f
C2791 _24_ p[7] 0.0129f
C2792 _07_ _45_/a_27_47# 1.02e-20
C2793 _03_ _27_/a_109_297# 1.97e-20
C2794 net11 _36_/a_27_47# 0.0717f
C2795 _14_ p[7] 0.186f
C2796 _10_ _03_ 0.00244f
C2797 _52_/a_584_47# _26_/a_29_53# 7.45e-20
C2798 net2 b[3] 0.00419f
C2799 th15_0/Vin input3/a_27_47# 0.00105f
C2800 net12 _01_ 1.67e-21
C2801 net19 th12_0/m1_529_n42# 4.2e-21
C2802 th14_0/m1_891_419# _42_/a_109_93# 1.58e-19
C2803 _22_ _53_/a_111_297# 4.7e-20
C2804 _02_ _38_/a_27_47# 0.00103f
C2805 net4 _12_ 0.105f
C2806 _50_/a_223_47# net5 0.00202f
C2807 _26_/a_183_297# _22_ 0.00184f
C2808 input12/a_27_47# p[7] 0.0892f
C2809 net18 p[7] 0.104f
C2810 _30_/a_297_297# b[1] 3.14e-19
C2811 input5/a_381_47# net19 0.00173f
C2812 net1 input2/a_27_47# 4.81e-19
C2813 _37_/a_27_47# _16_ 2.07e-19
C2814 net12 _04_ 0.267f
C2815 _18_ _02_ 2.96e-20
C2816 _25_ _36_/a_109_47# 3.76e-21
C2817 VGND _31_/a_285_297# -0.00136f
C2818 th15_0/Vin th02_0/m1_983_133# 0.0143f
C2819 _06_ _20_ 0.133f
C2820 _19_ th11_0/m1_577_n654# 3.11e-19
C2821 _26_/a_29_53# _02_ 0.0466f
C2822 net9 _03_ 0.149f
C2823 _33_/a_368_53# _05_ 9.2e-19
C2824 VGND net2 0.852f
C2825 _34_/a_377_297# _06_ 0.00427f
C2826 _22_ net1 0.0129f
C2827 net6 _40_/a_297_297# 7.47e-22
C2828 _45_/a_193_297# p[7] -0.00859f
C2829 VGND _44_/a_256_47# -0.00184f
C2830 net7 net1 0.0712f
C2831 input15/a_27_47# _18_ 8.27e-21
C2832 _34_/a_129_47# net10 0.003f
C2833 _12_ _50_/a_343_93# 5.63e-20
C2834 p[2] _20_ 3.01e-20
C2835 VGND _52_/a_584_47# -0.00112f
C2836 _15_ _50_/a_223_47# 0.00698f
C2837 net4 _45_/a_27_47# 0.024f
C2838 _42_/a_109_93# net17 3.1e-21
C2839 _32_/a_303_47# p[7] 6.03e-19
C2840 _30_/a_215_297# _36_/a_27_47# 7.13e-20
C2841 _11_ p[8] 6.68e-20
C2842 net13 net10 0.375f
C2843 input1/a_75_212# b[1] 0.0074f
C2844 _17_ p[9] 1.03e-20
C2845 p[14] input6/a_27_47# 0.0235f
C2846 _47_/a_81_21# net2 4.95e-19
C2847 input15/a_27_47# b[3] 1.77e-19
C2848 _10_ _00_ 0.301f
C2849 _49_/a_201_297# _03_ 0.00842f
C2850 _10_ _36_/a_27_47# 0.00109f
C2851 _55_/a_80_21# _00_ 5.5e-19
C2852 _06_ _50_/a_27_47# 0.00972f
C2853 _17_ net19 0.0269f
C2854 _55_/a_472_297# _16_ 3.71e-19
C2855 input5/a_664_47# input7/a_27_47# 1.08e-21
C2856 _03_ _05_ 0.135f
C2857 _41_/a_59_75# _47_/a_299_297# 0.00146f
C2858 _31_/a_117_297# p[10] 1.09e-19
C2859 net12 net1 1.17e-19
C2860 p[7] _20_ 0.341f
C2861 _03_ _31_/a_35_297# 0.00749f
C2862 _06_ net8 0.00282f
C2863 p[12] _39_/a_47_47# 0.00138f
C2864 _06_ _29_/a_29_53# 0.00111f
C2865 VGND _02_ 1.63f
C2866 th10_0/m1_536_174# b[3] 0.00833f
C2867 _34_/a_377_297# p[7] -0.00132f
C2868 p[11] _44_/a_250_297# 0.00177f
C2869 _20_ th15_0/m1_849_n157# 2.76e-21
C2870 _11_ _37_/a_27_47# 0.0018f
C2871 _06_ net11 0.546f
C2872 net2 output17/a_27_47# 0.0285f
C2873 p[7] p[11] 0.401f
C2874 input5/a_841_47# _21_ 1.59e-21
C2875 p[2] net8 0.0146f
C2876 _12_ net5 0.983f
C2877 input2/a_27_47# p[10] 0.0095f
C2878 net2 _44_/a_584_47# 0.0053f
C2879 p[1] net17 8.41e-20
C2880 th15_0/Vin _39_/a_47_47# 8.52e-22
C2881 net11 output18/a_27_47# 6.84e-20
C2882 _47_/a_299_297# _11_ 0.00738f
C2883 VGND _28_/a_109_297# -9.87e-19
C2884 net9 _00_ 0.00501f
C2885 net9 _36_/a_27_47# 0.00493f
C2886 VGND _30_/a_109_53# -0.0072f
C2887 net3 net14 0.689f
C2888 VGND input15/a_27_47# 0.0158f
C2889 Vin net14 0.00129f
C2890 _47_/a_81_21# _02_ 1.59e-20
C2891 _52_/a_93_21# _12_ 0.0157f
C2892 _04_ _29_/a_183_297# 0.0015f
C2893 p[7] _50_/a_27_47# -0.00335f
C2894 _12_ b[1] 3.18e-21
C2895 _14_ net17 2.4e-20
C2896 net12 _33_/a_296_53# 1.23e-20
C2897 net7 p[10] 0.00695f
C2898 _35_/a_76_199# _33_/a_109_93# 3.08e-19
C2899 VGND th10_0/m1_536_174# 0.0658f
C2900 p[7] net8 0.702f
C2901 VGND _23_ 0.16f
C2902 p[7] _29_/a_29_53# 0.0303f
C2903 Vin _38_/a_27_47# 5.31e-19
C2904 _15_ _12_ 0.00833f
C2905 net11 p[7] 1.14f
C2906 net13 net15 8.84e-19
C2907 _32_/a_197_47# net8 3.39e-20
C2908 _45_/a_27_47# net5 0.0288f
C2909 th15_0/Vin _44_/a_93_21# 0.00197f
C2910 Vin th02_0/m1_571_144# 8.17e-20
C2911 _36_/a_27_47# _05_ 3.67e-21
C2912 _05_ _00_ 5.03e-22
C2913 _17_ _01_ 1.46e-20
C2914 _18_ net3 7.34e-20
C2915 th15_0/Vin th11_0/m1_705_187# 0.0346f
C2916 Vin _18_ 3.79e-21
C2917 _36_/a_303_47# net5 0.00256f
C2918 net9 input13/a_27_47# 2.42e-19
C2919 _06_ _30_/a_215_297# 2.03e-20
C2920 _25_ _12_ 1.23e-20
C2921 p[1] input7/a_27_47# 0.0164f
C2922 net6 _39_/a_129_47# 6.91e-19
C2923 net4 _39_/a_285_47# 9.71e-19
C2924 _10_ _41_/a_145_75# 0.00148f
C2925 _19_ p[13] 0.00101f
C2926 _10_ _39_/a_377_297# 7.42e-19
C2927 th03_0/m1_890_n844# th02_0/m1_983_133# 0.0135f
C2928 _26_/a_29_53# net3 2.83e-21
C2929 _52_/a_93_21# _45_/a_27_47# 1.18e-19
C2930 _10_ _06_ 1.14f
C2931 _14_ _40_/a_297_297# 1.58e-19
C2932 th14_0/m1_891_419# p[11] 0.0117f
C2933 _06_ _55_/a_80_21# 5.15e-19
C2934 p[12] net15 1.84e-19
C2935 _04_ _17_ 4.34e-19
C2936 input5/a_381_47# net1 1.27e-19
C2937 p[13] net5 0.012f
C2938 _32_/a_27_47# _22_ 1.76e-19
C2939 p[13] input14/a_27_47# 3.88e-19
C2940 b[3] net3 2.43e-20
C2941 Vin b[3] 0.0166f
C2942 p[8] th12_0/m1_529_n42# 0.00973f
C2943 _43_/a_369_47# net14 6.79e-21
C2944 _09_ _48_/a_27_47# 0.00541f
C2945 _32_/a_27_47# _11_ 1.65e-20
C2946 net7 _32_/a_27_47# 0.00559f
C2947 _54_/a_75_212# _02_ 6.6e-20
C2948 _45_/a_109_297# _12_ 0.00587f
C2949 _22_ input3/a_27_47# 5.13e-20
C2950 net2 p[9] 0.00112f
C2951 p[9] th09_0/m1_962_372# 5.57e-19
C2952 _44_/a_93_21# input5/a_558_47# 2.71e-19
C2953 _02_ net16 8.94e-19
C2954 net13 _33_/a_368_53# 2.1e-20
C2955 th15_0/Vin net15 0.00757f
C2956 _10_ output19/a_27_47# 2.79e-20
C2957 p[7] _30_/a_465_297# -4.57e-19
C2958 net2 net19 0.599f
C2959 input13/a_27_47# _05_ 3.93e-19
C2960 p[13] b[1] 0.00201f
C2961 _04_ _27_/a_277_297# 0.00113f
C2962 th14_0/m1_891_419# net8 2.46e-21
C2963 _06_ net9 0.0505f
C2964 _06_ _50_/a_515_93# 0.00244f
C2965 _43_/a_193_413# _44_/a_93_21# 0.0161f
C2966 _15_ input6/a_27_47# 4.43e-19
C2967 _02_ _21_ 0.397f
C2968 p[7] _30_/a_215_297# -0.00497f
C2969 _10_ _38_/a_303_47# 7.36e-19
C2970 _20_ net17 4e-20
C2971 p[7] _27_/a_109_297# -2.45e-19
C2972 _06_ _53_/a_29_53# 0.0709f
C2973 _10_ p[7] 0.577f
C2974 _32_/a_27_47# net12 1.52e-19
C2975 VGND net3 0.323f
C2976 p[7] _55_/a_80_21# 0.0289f
C2977 _25_ _36_/a_303_47# 2.03e-21
C2978 VGND Vin 0.768f
C2979 _43_/a_27_47# net14 4.87e-20
C2980 _35_/a_226_47# _02_ 2.21e-19
C2981 net9 p[2] 1.4e-20
C2982 _10_ th15_0/m1_849_n157# 1.54e-19
C2983 _43_/a_369_47# _18_ 1.49e-19
C2984 _09_ _22_ 0.0279f
C2985 _53_/a_29_53# output18/a_27_47# 9.46e-19
C2986 _30_/a_109_53# _21_ 3.31e-20
C2987 _06_ _42_/a_209_311# 1.66e-19
C2988 _09_ _11_ 0.0665f
C2989 net13 _03_ 0.271f
C2990 _09_ net7 0.00258f
C2991 p[7] th13_0/m1_831_275# 0.0295f
C2992 input5/a_558_47# net15 0.00672f
C2993 th13_0/m1_831_275# th15_0/m1_849_n157# 5.99e-19
C2994 net12 _35_/a_489_413# 3.97e-20
C2995 _09_ _49_/a_208_47# 5.43e-21
C2996 _02_ net19 0.0474f
C2997 th15_0/Vin _37_/a_109_47# 5.47e-20
C2998 _06_ _05_ 0.00724f
C2999 _47_/a_81_21# net3 6.66e-19
C3000 net10 _30_/a_392_297# 3.4e-19
C3001 _23_ _21_ 0.0217f
C3002 Vin th10_0/m1_502_n495# 9.53e-19
C3003 _39_/a_285_47# net5 0.05f
C3004 _43_/a_193_413# net15 0.00169f
C3005 net9 p[7] 0.535f
C3006 _40_/a_297_297# _20_ 9.18e-21
C3007 p[7] _50_/a_515_93# -5.03e-19
C3008 _55_/a_217_297# net15 7.79e-19
C3009 p[0] th02_0/m1_571_144# 0.0179f
C3010 _48_/a_27_47# net10 0.00377f
C3011 net11 _29_/a_111_297# 8.27e-19
C3012 _27_/a_27_297# net14 0.0118f
C3013 p[2] _49_/a_201_297# 8.68e-20
C3014 net8 net17 0.18f
C3015 input15/a_27_47# p[9] 0.0194f
C3016 p[7] _53_/a_29_53# 0.00821f
C3017 _43_/a_27_47# _18_ 0.0201f
C3018 p[2] _05_ 5.07e-19
C3019 _09_ net12 0.0374f
C3020 _23_ _35_/a_226_47# 4.21e-19
C3021 net9 _32_/a_197_47# 6.06e-19
C3022 _08_ _35_/a_76_199# 0.0061f
C3023 _01_ _31_/a_285_297# 1.92e-19
C3024 net11 net17 3.19e-20
C3025 input15/a_27_47# net19 0.00231f
C3026 p[2] _31_/a_35_297# 0.00277f
C3027 net6 _50_/a_223_47# 0.0194f
C3028 net4 _50_/a_343_93# 0.00124f
C3029 _44_/a_93_21# _16_ 0.00354f
C3030 VGND _40_/a_191_297# -9.29e-19
C3031 _13_ _50_/a_223_47# 8.2e-20
C3032 output17/a_27_47# net3 0.00248f
C3033 Vin output17/a_27_47# 0.00661f
C3034 _09_ _45_/a_465_47# 2.77e-19
C3035 _52_/a_256_47# _06_ 0.00207f
C3036 p[7] _42_/a_209_311# -0.00753f
C3037 _17_ _37_/a_27_47# 0.00277f
C3038 th10_0/m1_536_174# p[9] 0.185f
C3039 net2 _01_ 2.72e-19
C3040 _07_ b[1] 0.0417f
C3041 _49_/a_75_199# p[13] 1.23e-19
C3042 _44_/a_346_47# net14 0.00464f
C3043 input2/a_27_47# net10 1.17e-20
C3044 _06_ input4/a_75_212# 0.00205f
C3045 VGND _43_/a_369_47# -8.43e-19
C3046 VGND b[0] 0.181f
C3047 p[7] _49_/a_201_297# 0.0175f
C3048 _29_/a_29_53# input9/a_75_212# 9.7e-21
C3049 _11_ _39_/a_47_47# 3.9e-19
C3050 p[7] _05_ 0.118f
C3051 _32_/a_109_47# _02_ 3.98e-19
C3052 net1 input5/a_841_47# 1.33e-19
C3053 p[14] th09_0/m1_485_n505# 1.95e-20
C3054 _52_/a_250_297# b[2] 1.6e-19
C3055 _04_ net2 0.158f
C3056 net11 input9/a_75_212# 1.1e-20
C3057 p[7] _31_/a_35_297# 0.0284f
C3058 net13 _36_/a_27_47# 0.0488f
C3059 net7 net10 1.65e-36
C3060 _52_/a_584_47# _04_ 2.5e-19
C3061 Vin th13_0/m1_559_n458# 2.77e-19
C3062 _35_/a_226_297# net13 6.88e-19
C3063 input5/a_62_47# _44_/a_250_297# 2.45e-20
C3064 _16_ net15 0.214f
C3065 _24_ b[2] 1.85e-19
C3066 th11_0/m1_705_187# input2/a_27_47# 3e-19
C3067 input7/a_27_47# net8 2.03e-21
C3068 net4 net5 0.0447f
C3069 _52_/a_256_47# p[7] -9.47e-19
C3070 p[7] input5/a_62_47# 0.0601f
C3071 Vin net16 3.38e-19
C3072 _02_ _01_ 0.106f
C3073 p[0] VGND 0.423f
C3074 VGND _43_/a_27_47# -0.0153f
C3075 th03_0/m1_638_n591# p[1] 0.135f
C3076 _30_/a_215_297# net17 4.69e-20
C3077 p[7] input4/a_75_212# 0.0608f
C3078 net18 b[2] 0.0131f
C3079 _52_/a_93_21# net4 7.93e-20
C3080 _11_ _44_/a_93_21# 4.78e-20
C3081 _03_ _27_/a_205_297# 1.46e-20
C3082 VGND _33_/a_109_93# -0.0132f
C3083 input5/a_841_47# _37_/a_27_47# 4.64e-20
C3084 net12 net10 0.539f
C3085 net7 th11_0/m1_705_187# 1.13e-19
C3086 net1 _31_/a_285_297# 5.85e-19
C3087 _04_ _02_ 0.0541f
C3088 input10/a_27_47# p[7] 0.0547f
C3089 _15_ p[14] 0.00339f
C3090 _02_ _38_/a_109_47# 1.63e-19
C3091 th14_0/m1_891_419# _42_/a_209_311# 6.86e-21
C3092 input13/a_27_47# net13 0.00139f
C3093 net1 net2 1.64e-19
C3094 th15_0/Vin _00_ 1.03e-19
C3095 net6 _12_ 0.0891f
C3096 _50_/a_343_93# net5 0.00124f
C3097 net4 _15_ 0.00427f
C3098 _12_ _13_ 0.462f
C3099 _41_/a_59_75# net15 1.16e-20
C3100 input2/a_27_47# net15 1.61e-19
C3101 _07_ _49_/a_75_199# 4.05e-21
C3102 _09_ _29_/a_183_297# 4.51e-20
C3103 input9/a_75_212# _30_/a_215_297# 6.24e-21
C3104 _04_ _30_/a_109_53# 9.19e-21
C3105 p[9] net3 1.63e-19
C3106 VGND _27_/a_27_297# -0.0157f
C3107 Vin p[9] 0.112f
C3108 _53_/a_111_297# _02_ 9.57e-20
C3109 net9 _29_/a_111_297# 8.06e-21
C3110 _42_/a_109_93# th14_0/m1_641_n318# 1.75e-19
C3111 net2 p[8] 0.0279f
C3112 _20_ _39_/a_129_47# 1.71e-20
C3113 _10_ input9/a_75_212# 5.49e-21
C3114 net19 net3 0.611f
C3115 Vin net19 1.54e-19
C3116 p[0] output17/a_27_47# 0.00839f
C3117 _06_ _36_/a_197_47# 6.18e-19
C3118 _22_ net15 2.74e-19
C3119 b[0] th13_0/m1_559_n458# 5.75e-19
C3120 net9 net17 1.26e-20
C3121 _11_ net15 0.145f
C3122 net7 net15 2.91e-19
C3123 _34_/a_47_47# _07_ 0.011f
C3124 _34_/a_129_47# _06_ 5.3e-19
C3125 VGND _44_/a_346_47# -0.00198f
C3126 _45_/a_205_47# p[7] -1.62e-19
C3127 _34_/a_285_47# net10 0.0454f
C3128 b[0] net16 0.0306f
C3129 _35_/a_76_199# _18_ 6.82e-21
C3130 th14_0/m1_891_419# input5/a_62_47# 0.00116f
C3131 _19_ net5 6.41e-21
C3132 _15_ _50_/a_343_93# 0.0098f
C3133 _06_ net13 0.0758f
C3134 net2 _37_/a_27_47# 0.0692f
C3135 p[2] input8/a_27_47# 0.0217f
C3136 net1 _02_ 0.00251f
C3137 _10_ _53_/a_183_297# 2.86e-19
C3138 input1/a_75_212# p[1] 0.0023f
C3139 Vin output16/a_27_47# 3.69e-19
C3140 net4 _45_/a_109_297# 6.43e-20
C3141 net6 _45_/a_27_47# 0.021f
C3142 _42_/a_209_311# net17 1.04e-21
C3143 _45_/a_27_47# _13_ 0.0703f
C3144 net9 input9/a_75_212# 0.0245f
C3145 _43_/a_193_413# _00_ 0.00721f
C3146 _47_/a_299_297# net2 1.18e-19
C3147 VGND _48_/a_181_47# 3.03e-19
C3148 _03_ _30_/a_392_297# 6.33e-19
C3149 net6 _36_/a_303_47# 1.25e-19
C3150 th03_0/m1_890_n844# _03_ 3.64e-21
C3151 _19_ b[1] 0.00967f
C3152 _05_ net17 0.0111f
C3153 net1 _30_/a_109_53# 0.0297f
C3154 th01_0/m1_991_n1219# p[1] 5.78e-20
C3155 net6 input6/a_27_47# 0.00208f
C3156 _31_/a_285_297# p[10] 4.45e-20
C3157 _52_/a_93_21# net5 0.0124f
C3158 _03_ _31_/a_117_297# 5.32e-19
C3159 p[12] _41_/a_145_75# 4.82e-19
C3160 p[7] _36_/a_197_47# -5.24e-19
C3161 p[12] _39_/a_377_297# 4.68e-19
C3162 net17 _31_/a_35_297# 0.0514f
C3163 th15_0/Vin th01_0/m1_571_n501# 0.00971f
C3164 b[1] net5 0.00349f
C3165 _06_ p[12] 0.0132f
C3166 input8/a_27_47# p[7] 0.0886f
C3167 _34_/a_129_47# p[7] -9.23e-19
C3168 _15_ _19_ 1.46e-20
C3169 net2 p[10] 0.0373f
C3170 _15_ net5 0.0352f
C3171 input2/a_27_47# _03_ 2.71e-19
C3172 p[7] net13 0.615f
C3173 th15_0/Vin _41_/a_145_75# 1.73e-19
C3174 _52_/a_93_21# b[1] 2.82e-19
C3175 _47_/a_384_47# _11_ 7.23e-20
C3176 input9/a_75_212# _05_ 1.24e-21
C3177 _06_ th15_0/Vin 0.00739f
C3178 input5/a_664_47# p[13] 0.0024f
C3179 _44_/a_93_21# th12_0/m1_529_n42# 7.97e-20
C3180 net3 _01_ 1.16e-19
C3181 Vin _01_ 5.85e-20
C3182 _33_/a_109_93# _21_ 1.62e-20
C3183 VGND _35_/a_76_199# -0.0034f
C3184 th10_0/m1_536_174# p[8] 0.0134f
C3185 net11 b[2] 1.46e-19
C3186 _52_/a_250_297# _12_ 0.0139f
C3187 _25_ net5 6.42e-19
C3188 _22_ _03_ 2.55e-20
C3189 th15_0/Vin p[2] 1.51e-21
C3190 net12 _33_/a_368_53# 2.63e-19
C3191 _15_ b[1] 1.19e-19
C3192 input15/a_27_47# _37_/a_27_47# 3.27e-19
C3193 net7 _03_ 0.078f
C3194 _35_/a_76_199# _33_/a_209_311# 9.95e-21
C3195 _35_/a_226_47# _33_/a_109_93# 4.9e-19
C3196 _04_ net3 0.113f
C3197 _04_ Vin 0.00376f
C3198 th12_0/m1_394_n856# p[7] 0.00333f
C3199 b[0] output16/a_27_47# 0.014f
C3200 _16_ _00_ 0.00613f
C3201 _17_ _39_/a_47_47# 1.47e-20
C3202 th15_0/Vin output19/a_27_47# 0.0163f
C3203 VGND _08_ 0.161f
C3204 p[7] p[12] 0.144f
C3205 _12_ _24_ 1.67e-19
C3206 _20_ _50_/a_223_47# 1.71e-19
C3207 _14_ _12_ 1.98e-20
C3208 _55_/a_300_47# _22_ 2.08e-19
C3209 _49_/a_208_47# _03_ 3.86e-19
C3210 p[12] th15_0/m1_849_n157# 0.0103f
C3211 _25_ b[1] 0.0015f
C3212 _45_/a_109_297# net5 0.0184f
C3213 th15_0/Vin _44_/a_250_297# 7.01e-19
C3214 _06_ input5/a_558_47# 3.55e-19
C3215 _08_ _33_/a_209_311# 0.0122f
C3216 _18_ net14 0.0147f
C3217 net2 input3/a_27_47# 0.0229f
C3218 th12_0/m1_529_n42# net15 2.01e-21
C3219 _49_/a_75_199# _19_ 0.0206f
C3220 _55_/a_472_297# _02_ 1.25e-19
C3221 th15_0/Vin p[7] 0.945f
C3222 net18 _12_ 8.24e-19
C3223 net6 _39_/a_285_47# 1.53e-19
C3224 net12 _03_ 0.0268f
C3225 th15_0/Vin th15_0/m1_849_n157# 0.173f
C3226 _10_ _39_/a_129_47# 2.51e-19
C3227 _13_ _39_/a_285_47# 0.00451f
C3228 _06_ _43_/a_193_413# 0.0138f
C3229 _26_/a_29_53# net14 1.33e-20
C3230 _07_ _13_ 3.22e-23
C3231 input5/a_381_47# net15 7.15e-19
C3232 net8 _30_/a_297_297# 2.42e-21
C3233 _06_ _55_/a_217_297# 3.46e-19
C3234 _41_/a_59_75# _00_ 2.43e-20
C3235 b[3] net14 8.65e-19
C3236 _17_ _44_/a_93_21# 0.0646f
C3237 _27_/a_27_297# net19 1.98e-19
C3238 _43_/a_469_47# net14 1.44e-20
C3239 _45_/a_27_47# _24_ 4.57e-19
C3240 _45_/a_193_297# _12_ 0.0103f
C3241 net2 th02_0/m1_983_133# 3.55e-19
C3242 net1 net3 4.25e-20
C3243 net1 Vin 0.00771f
C3244 _29_/a_29_53# _50_/a_223_47# 1.45e-20
C3245 p[11] th14_0/m1_641_n318# 0.114f
C3246 _49_/a_75_199# b[1] 0.00805f
C3247 _32_/a_27_47# _02_ 0.00247f
C3248 _22_ _00_ 0.477f
C3249 _22_ _36_/a_27_47# 2.82e-20
C3250 p[7] input5/a_558_47# 0.0083f
C3251 _44_/a_346_47# net19 0.00124f
C3252 _11_ _00_ 0.238f
C3253 net7 _00_ 8.12e-21
C3254 _06_ _50_/a_615_93# 0.00264f
C3255 p[8] net3 1.87e-19
C3256 Vin p[8] 0.564f
C3257 _14_ input6/a_27_47# 3.75e-21
C3258 _18_ _26_/a_29_53# 5.26e-20
C3259 p[7] _27_/a_205_297# 1.05e-19
C3260 _43_/a_193_413# p[7] 0.0063f
C3261 _32_/a_27_47# _30_/a_109_53# 1.51e-19
C3262 _34_/a_47_47# b[1] 0.0197f
C3263 VGND net14 0.441f
C3264 p[7] _55_/a_217_297# -0.00133f
C3265 _43_/a_27_47# _01_ 9.77e-20
C3266 _35_/a_489_413# _02_ 3.86e-19
C3267 net6 p[14] 0.00518f
C3268 _12_ _20_ 3.9e-19
C3269 _17_ net15 0.195f
C3270 _43_/a_469_47# _18_ 1.59e-19
C3271 _06_ _16_ 0.00162f
C3272 th15_0/Vin th14_0/m1_891_419# 0.0726f
C3273 net4 net6 0.713f
C3274 _35_/a_76_199# _21_ 0.0175f
C3275 net13 net17 5.21e-20
C3276 net4 _13_ 0.212f
C3277 _40_/a_109_297# net15 0.0016f
C3278 _37_/a_27_47# net3 0.094f
C3279 Vin _37_/a_27_47# 2.88e-19
C3280 net12 _36_/a_27_47# 0.0185f
C3281 _53_/a_29_53# b[2] 6.22e-19
C3282 _09_ _02_ 0.297f
C3283 VGND _38_/a_27_47# 0.00767f
C3284 _30_/a_215_297# _30_/a_297_297# -8.88e-34
C3285 input8/a_27_47# input9/a_75_212# 3.09e-20
C3286 _35_/a_76_199# _35_/a_226_47# -2.84e-32
C3287 th15_0/Vin _37_/a_197_47# 1.87e-19
C3288 _47_/a_299_297# net3 2.55e-19
C3289 _06_ _48_/a_27_47# 0.0251f
C3290 Vin 0 11.5f
C3291 th11_0/m1_705_187# 0 0.602f
C3292 p[10] 0 0.502f
C3293 th11_0/m1_577_n654# 0 0.286f
C3294 th13_0/m1_831_275# 0 1.05f
C3295 p[12] 0 0.639f
C3296 th13_0/m1_559_n458# 0 0.286f
C3297 _03_ 0 0.36f
C3298 net10 0 0.418f
C3299 _30_/a_109_53# 0 0.159f
C3300 _30_/a_215_297# 0 0.142f
C3301 p[14] 0 0.608f
C3302 th15_0/m1_849_n157# 0 1.28f
C3303 th15_0/m1_597_n912# 0 0.19f
C3304 _05_ 0 0.152f
C3305 _31_/a_285_297# 0 0.00137f
C3306 _31_/a_35_297# 0 0.255f
C3307 _32_/a_27_47# 0 0.175f
C3308 _50_/a_343_93# 0 0.172f
C3309 _50_/a_223_47# 0 0.141f
C3310 _50_/a_27_47# 0 0.259f
C3311 _07_ 0 0.285f
C3312 _06_ 0 0.779f
C3313 _33_/a_209_311# 0 0.143f
C3314 _33_/a_109_93# 0 0.158f
C3315 _34_/a_285_47# 0 0.0174f
C3316 _34_/a_47_47# 0 0.199f
C3317 _23_ 0 0.106f
C3318 _09_ 0 0.142f
C3319 _08_ 0 0.128f
C3320 _35_/a_489_413# 0 0.0254f
C3321 _35_/a_226_47# 0 0.162f
C3322 _35_/a_76_199# 0 0.141f
C3323 input15/a_27_47# 0 0.208f
C3324 _24_ 0 0.135f
C3325 _12_ 0 0.378f
C3326 _52_/a_250_297# 0 0.0278f
C3327 _52_/a_93_21# 0 0.151f
C3328 _10_ 0 0.624f
C3329 _36_/a_27_47# 0 0.175f
C3330 _53_/a_29_53# 0 0.18f
C3331 input14/a_27_47# 0 0.208f
C3332 VGND 0 23.7f
C3333 p[0] 0 0.808f
C3334 th01_0/m1_991_n1219# 0 1.24f
C3335 th01_0/m1_571_n501# 0 0.194f
C3336 th15_0/Vin 0 6.95f
C3337 _11_ 0 0.265f
C3338 _37_/a_27_47# 0 0.175f
C3339 net13 0 0.377f
C3340 input13/a_27_47# 0 0.208f
C3341 net18 0 0.207f
C3342 _25_ 0 0.191f
C3343 _54_/a_75_212# 0 0.21f
C3344 _38_/a_27_47# 0 0.175f
C3345 net19 0 0.165f
C3346 _22_ 0 0.215f
C3347 _14_ 0 0.225f
C3348 _15_ 0 0.331f
C3349 _55_/a_217_297# 0 0.00117f
C3350 _55_/a_80_21# 0 0.21f
C3351 input12/a_27_47# 0 0.208f
C3352 net9 0 0.285f
C3353 input9/a_75_212# 0 0.21f
C3354 _39_/a_285_47# 0 0.0174f
C3355 _39_/a_47_47# 0 0.199f
C3356 input11/a_27_47# 0 0.208f
C3357 net8 0 0.386f
C3358 input8/a_27_47# 0 0.208f
C3359 p[2] 0 0.644f
C3360 th03_0/m1_890_n844# 0 1.05f
C3361 th03_0/m1_638_n591# 0 0.224f
C3362 input10/a_27_47# 0 0.208f
C3363 net7 0 0.449f
C3364 input7/a_27_47# 0 0.208f
C3365 p[9] 0 0.698f
C3366 th10_0/m1_536_174# 0 0.825f
C3367 th10_0/m1_502_n495# 0 0.146f
C3368 input6/a_27_47# 0 0.208f
C3369 net5 0 0.817f
C3370 input5/a_841_47# 0 0.0929f
C3371 input5/a_664_47# 0 0.13f
C3372 input5/a_558_47# 0 0.164f
C3373 input5/a_381_47# 0 0.11f
C3374 input5/a_62_47# 0 0.169f
C3375 input4/a_75_212# 0 0.21f
C3376 th12_0/m1_529_n42# 0 0.861f
C3377 p[11] 0 0.505f
C3378 th12_0/m1_394_n856# 0 0.215f
C3379 input3/a_27_47# 0 0.208f
C3380 net2 0 0.68f
C3381 input2/a_27_47# 0 0.208f
C3382 net1 0 0.337f
C3383 input1/a_75_212# 0 0.21f
C3384 th14_0/m1_891_419# 0 1.48f
C3385 p[13] 0 0.763f
C3386 th14_0/m1_641_n318# 0 0.241f
C3387 b[3] 0 0.136f
C3388 output19/a_27_47# 0 0.543f
C3389 th09_0/m1_485_n505# 0 1.18f
C3390 p[8] 0 0.623f
C3391 th09_0/m1_962_372# 0 0.118f
C3392 b[2] 0 0.515f
C3393 output18/a_27_47# 0 0.543f
C3394 b[1] 0 0.281f
C3395 net17 0 0.169f
C3396 output17/a_27_47# 0 0.543f
C3397 _41_/a_59_75# 0 0.177f
C3398 b[0] 0 0.501f
C3399 output16/a_27_47# 0 0.543f
C3400 _16_ 0 0.125f
C3401 _42_/a_209_311# 0 0.143f
C3402 _42_/a_109_93# 0 0.158f
C3403 net6 0 0.533f
C3404 net4 0 0.315f
C3405 _26_/a_29_53# 0 0.18f
C3406 _43_/a_193_413# 0 0.136f
C3407 _43_/a_27_47# 0 0.224f
C3408 _01_ 0 0.15f
C3409 net14 0 0.502f
C3410 net3 0 0.453f
C3411 net15 0 0.446f
C3412 _27_/a_27_297# 0 0.163f
C3413 _18_ 0 0.143f
C3414 _17_ 0 0.242f
C3415 _44_/a_250_297# 0 0.0278f
C3416 _44_/a_93_21# 0 0.151f
C3417 net16 0 0.23f
C3418 _13_ 0 0.133f
C3419 _45_/a_193_297# 0 0.0011f
C3420 _45_/a_109_297# 0 7.11e-19
C3421 _45_/a_27_47# 0 0.216f
C3422 _00_ 0 0.377f
C3423 net11 0 0.755f
C3424 net12 0 0.511f
C3425 _29_/a_29_53# 0 0.18f
C3426 _19_ 0 0.113f
C3427 _04_ 0 0.334f
C3428 p[1] 0 0.451f
C3429 th02_0/m1_983_133# 0 1.44f
C3430 th02_0/m1_571_144# 0 0.252f
C3431 _47_/a_299_297# 0 0.0348f
C3432 _47_/a_81_21# 0 0.147f
C3433 p[7] 0 84.2f
C3434 _48_/a_27_47# 0 0.177f
C3435 _21_ 0 0.29f
C3436 _20_ 0 0.237f
C3437 _02_ 0 0.449f
C3438 _49_/a_201_297# 0 0.00345f
C3439 _49_/a_75_199# 0 0.205f
.ends

