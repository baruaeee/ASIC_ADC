* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : inv02f                                       *
* Netlisted  : Sun Dec  8 23:16:33 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733696178270                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733696178270 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.5e-07 W=8e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733696178270

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733696178271                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733696178271 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=2.85e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733696178271

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv02f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv02f 3 1 4 2
** N=9 EP=4 FDC=2
X0 1 2 3 pfet_01v8_CDNS_733696178270 $T=335 2855 0 0 $X=-110 $Y=2675
X1 4 2 3 nfet_01v8_CDNS_733696178271 $T=315 640 0 0 $X=-90 $Y=490
.ends inv02f
