magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 2432 29 2438
rect -29 2398 -17 2432
rect -29 2392 29 2398
rect -29 -2398 29 -2392
rect -29 -2432 -17 -2398
rect -29 -2438 29 -2432
<< pwell >>
rect -211 -2570 211 2570
<< nmos >>
rect -15 -2360 15 2360
<< ndiff >>
rect -73 2348 -15 2360
rect -73 -2348 -61 2348
rect -27 -2348 -15 2348
rect -73 -2360 -15 -2348
rect 15 2348 73 2360
rect 15 -2348 27 2348
rect 61 -2348 73 2348
rect 15 -2360 73 -2348
<< ndiffc >>
rect -61 -2348 -27 2348
rect 27 -2348 61 2348
<< psubdiff >>
rect -175 2500 -79 2534
rect 79 2500 175 2534
rect -175 2438 -141 2500
rect 141 2438 175 2500
rect -175 -2500 -141 -2438
rect 141 -2500 175 -2438
rect -175 -2534 -79 -2500
rect 79 -2534 175 -2500
<< psubdiffcont >>
rect -79 2500 79 2534
rect -175 -2438 -141 2438
rect 141 -2438 175 2438
rect -79 -2534 79 -2500
<< poly >>
rect -33 2432 33 2448
rect -33 2398 -17 2432
rect 17 2398 33 2432
rect -33 2382 33 2398
rect -15 2360 15 2382
rect -15 -2382 15 -2360
rect -33 -2398 33 -2382
rect -33 -2432 -17 -2398
rect 17 -2432 33 -2398
rect -33 -2448 33 -2432
<< polycont >>
rect -17 2398 17 2432
rect -17 -2432 17 -2398
<< locali >>
rect -175 2500 -79 2534
rect 79 2500 175 2534
rect -175 2438 -141 2500
rect 141 2438 175 2500
rect -33 2398 -17 2432
rect 17 2398 33 2432
rect -61 2348 -27 2364
rect -61 -2364 -27 -2348
rect 27 2348 61 2364
rect 27 -2364 61 -2348
rect -33 -2432 -17 -2398
rect 17 -2432 33 -2398
rect -175 -2500 -141 -2438
rect 141 -2500 175 -2438
rect -175 -2534 -79 -2500
rect 79 -2534 175 -2500
<< viali >>
rect -17 2398 17 2432
rect -61 -2348 -27 2348
rect 27 -2348 61 2348
rect -17 -2432 17 -2398
<< metal1 >>
rect -29 2432 29 2438
rect -29 2398 -17 2432
rect 17 2398 29 2432
rect -29 2392 29 2398
rect -67 2348 -21 2360
rect -67 -2348 -61 2348
rect -27 -2348 -21 2348
rect -67 -2360 -21 -2348
rect 21 2348 67 2360
rect 21 -2348 27 2348
rect 61 -2348 67 2348
rect 21 -2360 67 -2348
rect -29 -2398 29 -2392
rect -29 -2432 -17 -2398
rect 17 -2432 29 -2398
rect -29 -2438 29 -2432
<< properties >>
string FIXED_BBOX -158 -2517 158 2517
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 23.6 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
