* NGSPICE file created from adc.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_D7Y3TR a_n63_n101# a_n33_n75# a_n249_n145# a_63_n75#
+ a_n125_n75#
X0 a_63_n75# a_n63_n101# a_n33_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.233 pd=2.12 as=0.124 ps=1.08 w=0.75 l=0.15
X1 a_n33_n75# a_n63_n101# a_n125_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.08 as=0.233 ps=2.12 w=0.75 l=0.15
C0 a_n33_n75# a_63_n75# 0.113f
C1 a_n33_n75# a_n125_n75# 0.113f
C2 a_63_n75# a_n63_n101# 0.0104f
C3 a_n33_n75# a_n63_n101# 0.0186f
C4 a_n63_n101# a_n125_n75# 0.00451f
C5 a_63_n75# a_n249_n145# 0.0963f
C6 a_n33_n75# a_n249_n145# 0.0361f
C7 a_n125_n75# a_n249_n145# 0.105f
C8 a_n63_n101# a_n249_n145# 0.294f
.ends

.subckt sky130_fd_pr__pfet_01v8_2ZD99F w_n349_n261# a_n153_n139# a_n211_n42# a_153_n42#
+ VSUBS
X0 a_153_n42# a_n153_n139# a_n211_n42# w_n349_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.53
C0 a_n211_n42# a_153_n42# 0.0169f
C1 a_153_n42# a_n153_n139# 0.0177f
C2 a_n211_n42# a_n153_n139# 0.0177f
C3 a_153_n42# w_n349_n261# 0.0179f
C4 a_n211_n42# w_n349_n261# 0.034f
C5 w_n349_n261# a_n153_n139# 0.388f
C6 a_153_n42# VSUBS 0.0558f
C7 a_n211_n42# VSUBS 0.0456f
C8 a_n153_n139# VSUBS 0.556f
C9 w_n349_n261# VSUBS 1.16f
.ends

.subckt sky130_fd_pr__nfet_01v8_2BW22M a_154_n42# a_n154_n130# a_n314_n182# a_n212_n42#
X0 a_154_n42# a_n154_n130# a_n212_n42# a_n314_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.54
C0 a_154_n42# a_n212_n42# 0.0169f
C1 a_154_n42# a_n154_n130# 0.0178f
C2 a_n154_n130# a_n212_n42# 0.0178f
C3 a_154_n42# a_n314_n182# 0.0737f
C4 a_n212_n42# a_n314_n182# 0.0816f
C5 a_n154_n130# a_n314_n182# 0.924f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJP3BL a_15_n150# w_n211_n369# a_n73_n150# a_n33_n247#
+ VSUBS
X0 a_15_n150# a_n33_n247# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.15
C0 a_n73_n150# a_15_n150# 0.242f
C1 a_15_n150# a_n33_n247# 0.0267f
C2 a_n73_n150# a_n33_n247# 0.0267f
C3 a_15_n150# w_n211_n369# 0.0292f
C4 a_n73_n150# w_n211_n369# 0.0292f
C5 w_n211_n369# a_n33_n247# 0.19f
C6 a_15_n150# VSUBS 0.126f
C7 a_n73_n150# VSUBS 0.126f
C8 a_n33_n247# VSUBS 0.146f
C9 w_n211_n369# VSUBS 1.02f
.ends

.subckt sky130_fd_pr__nfet_01v8_LH5FDA a_n150_n130# a_276_n182# a_n208_n42# a_150_n42#
X0 a_150_n42# a_n150_n130# a_n208_n42# a_276_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.5
C0 a_150_n42# a_n208_n42# 0.0172f
C1 a_150_n42# a_n150_n130# 0.0176f
C2 a_n150_n130# a_n208_n42# 0.0176f
C3 a_150_n42# a_276_n182# 0.0815f
C4 a_n208_n42# a_276_n182# 0.0736f
C5 a_n150_n130# a_276_n182# 0.904f
.ends

.subckt th02 Vin V02 Vp m1_983_133# m1_571_144# Vn
XXM0 Vin Vn Vn m1_983_133# m1_983_133# sky130_fd_pr__nfet_01v8_D7Y3TR
XXM1 Vp Vin m1_571_144# m1_983_133# Vn sky130_fd_pr__pfet_01v8_2ZD99F
XXM2 m1_571_144# Vp Vn Vp sky130_fd_pr__nfet_01v8_2BW22M
XXM3 V02 Vp Vp m1_983_133# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_983_133# Vn V02 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 m1_571_144# Vn 0.00115f
C1 Vp V02 0.118f
C2 m1_983_133# V02 0.155f
C3 Vn Vin 0.0263f
C4 Vp m1_983_133# 0.366f
C5 m1_571_144# V02 0.011f
C6 m1_571_144# Vp 0.176f
C7 m1_571_144# m1_983_133# 0.0183f
C8 V02 Vin 0.00845f
C9 Vp Vin 0.25f
C10 m1_983_133# Vin 0.279f
C11 m1_571_144# Vin 0.332f
C12 V02 Vn 0.00239f
C13 Vp Vn 0.0235f
C14 m1_983_133# Vn 0.216f
C15 Vn 0 0.263f
C16 V02 0 0.334f
C17 m1_983_133# 0 1.44f
C18 Vp 0 3.16f
C19 m1_571_144# 0 0.252f
C20 Vin 0 0.949f
.ends

.subckt sky130_fd_pr__nfet_01v8_2V6S9N a_n216_n42# a_158_n42# a_n158_n130# a_n284_n216#
X0 a_158_n42# a_n158_n130# a_n216_n42# a_n284_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.58
C0 a_n216_n42# a_158_n42# 0.0165f
C1 a_n158_n130# a_158_n42# 0.018f
C2 a_n158_n130# a_n216_n42# 0.018f
C3 a_158_n42# a_n284_n216# 0.0746f
C4 a_n216_n42# a_n284_n216# 0.0746f
C5 a_n158_n130# a_n284_n216# 0.981f
.ends

.subckt sky130_fd_pr__pfet_01v8_XYZSMQ a_n33_n255# a_15_n158# w_n211_n377# a_n73_n158#
+ VSUBS
X0 a_15_n158# a_n33_n255# a_n73_n158# w_n211_n377# sky130_fd_pr__pfet_01v8 ad=0.458 pd=3.74 as=0.458 ps=3.74 w=1.58 l=0.15
C0 a_n33_n255# a_n73_n158# 0.0271f
C1 a_15_n158# a_n33_n255# 0.0271f
C2 w_n211_n377# a_n73_n158# 0.0299f
C3 a_15_n158# w_n211_n377# 0.0299f
C4 a_15_n158# a_n73_n158# 0.254f
C5 w_n211_n377# a_n33_n255# 0.191f
C6 a_15_n158# VSUBS 0.132f
C7 a_n73_n158# VSUBS 0.132f
C8 a_n33_n255# VSUBS 0.146f
C9 w_n211_n377# VSUBS 1.04f
.ends

.subckt sky130_fd_pr__pfet_01v8_AZD9DW w_n353_n261# a_n157_n139# a_n215_n42# a_157_n42#
+ VSUBS
X0 a_157_n42# a_n157_n139# a_n215_n42# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.57
C0 a_n157_n139# a_n215_n42# 0.0179f
C1 a_157_n42# a_n157_n139# 0.0179f
C2 w_n353_n261# a_n215_n42# 0.0179f
C3 a_157_n42# w_n353_n261# 0.0323f
C4 a_157_n42# a_n215_n42# 0.0166f
C5 w_n353_n261# a_n157_n139# 0.396f
C6 a_157_n42# VSUBS 0.0468f
C7 a_n215_n42# VSUBS 0.0559f
C8 a_n157_n139# VSUBS 0.569f
C9 w_n353_n261# VSUBS 1.17f
.ends

.subckt sky130_fd_pr__nfet_01v8_T8HSQ7 a_n175_n297# a_15_n157# a_n33_n245# a_n73_n157#
X0 a_15_n157# a_n33_n245# a_n73_n157# a_n175_n297# sky130_fd_pr__nfet_01v8 ad=0.455 pd=3.72 as=0.455 ps=3.72 w=1.57 l=0.15
C0 a_n73_n157# a_15_n157# 0.253f
C1 a_n33_n245# a_15_n157# 0.0289f
C2 a_n33_n245# a_n73_n157# 0.0289f
C3 a_15_n157# a_n175_n297# 0.161f
C4 a_n73_n157# a_n175_n297# 0.188f
C5 a_n33_n245# a_n175_n297# 0.322f
.ends

.subckt th09 V09 Vin Vn m1_485_n505# Vp m1_962_372#
XXM0 m1_485_n505# Vn Vin Vn sky130_fd_pr__nfet_01v8_2V6S9N
XXM1 Vin m1_485_n505# Vp Vp Vn sky130_fd_pr__pfet_01v8_XYZSMQ
XXM2 Vp m1_485_n505# Vp m1_962_372# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM3 Vp m1_485_n505# V09 m1_962_372# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM4 Vn V09 m1_485_n505# Vn sky130_fd_pr__nfet_01v8_T8HSQ7
C0 Vin V09 2.77e-19
C1 Vin Vn 0.0386f
C2 Vp m1_962_372# 0.0579f
C3 Vp Vin 0.187f
C4 m1_485_n505# m1_962_372# 0.0822f
C5 V09 Vn 0.00364f
C6 m1_485_n505# Vin 0.372f
C7 Vp V09 0.0743f
C8 Vp Vn 0.0176f
C9 Vin m1_962_372# 0.00821f
C10 m1_485_n505# V09 0.104f
C11 m1_485_n505# Vn 0.0846f
C12 m1_485_n505# Vp 0.372f
C13 V09 m1_962_372# 0.00205f
C14 Vn m1_962_372# 6.71e-21
C15 Vin 0 1.1f
C16 m1_485_n505# 0 1.18f
C17 V09 0 0.27f
C18 Vn 0 0.344f
C19 Vp 0 3.27f
C20 m1_962_372# 0 0.118f
.ends

.subckt sky130_fd_pr__pfet_01v8_HPNF99 a_n33_n147# a_23_n50# a_n81_n50# w_n219_n269#
+ VSUBS
X0 a_23_n50# a_n33_n147# a_n81_n50# w_n219_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.23
C0 w_n219_n269# a_23_n50# 0.0185f
C1 a_n81_n50# a_23_n50# 0.07f
C2 w_n219_n269# a_n33_n147# 0.173f
C3 a_n33_n147# a_n81_n50# 0.00814f
C4 w_n219_n269# a_n81_n50# 0.0419f
C5 a_n33_n147# a_23_n50# 0.00814f
C6 a_23_n50# VSUBS 0.0578f
C7 a_n81_n50# VSUBS 0.0428f
C8 a_n33_n147# VSUBS 0.157f
C9 w_n219_n269# VSUBS 0.779f
.ends

.subckt sky130_fd_pr__nfet_01v8_JZU22M a_n213_n42# a_155_n42# a_n155_n130# a_281_n238#
X0 a_155_n42# a_n155_n130# a_n213_n42# a_281_n238# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.55
C0 a_n155_n130# a_n213_n42# 0.0178f
C1 a_n213_n42# a_155_n42# 0.0168f
C2 a_n155_n130# a_155_n42# 0.0178f
C3 a_155_n42# a_281_n238# 0.0816f
C4 a_n213_n42# a_281_n238# 0.0737f
C5 a_n155_n130# a_281_n238# 0.928f
.ends

.subckt sky130_fd_pr__pfet_01v8_TM5S5A a_n80_n147# a_n138_n50# a_80_n50# w_n276_n269#
+ VSUBS
X0 a_80_n50# a_n80_n147# a_n138_n50# w_n276_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.8
C0 w_n276_n269# a_80_n50# 0.0231f
C1 a_n138_n50# a_80_n50# 0.0335f
C2 w_n276_n269# a_n80_n147# 0.297f
C3 a_n80_n147# a_n138_n50# 0.0141f
C4 w_n276_n269# a_n138_n50# 0.0231f
C5 a_n80_n147# a_80_n50# 0.0141f
C6 a_80_n50# VSUBS 0.0565f
C7 a_n138_n50# VSUBS 0.0565f
C8 a_n80_n147# VSUBS 0.296f
C9 w_n276_n269# VSUBS 1.01f
.ends

.subckt sky130_fd_pr__pfet_01v8_AM8GZ5 w_n526_n261# a_n330_n139# a_330_n42# a_n388_n42#
+ VSUBS
X0 a_330_n42# a_n330_n139# a_n388_n42# w_n526_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.3
C0 w_n526_n261# a_330_n42# 0.0408f
C1 a_n388_n42# a_330_n42# 0.00853f
C2 w_n526_n261# a_n330_n139# 0.719f
C3 a_n330_n139# a_n388_n42# 0.0223f
C4 w_n526_n261# a_n388_n42# 0.0179f
C5 a_n330_n139# a_330_n42# 0.0223f
C6 a_330_n42# VSUBS 0.0435f
C7 a_n388_n42# VSUBS 0.0585f
C8 a_n330_n139# VSUBS 1.13f
C9 w_n526_n261# VSUBS 1.76f
.ends

.subckt sky130_fd_pr__nfet_01v8_H7HSAV a_n73_n250# a_15_n250# a_n33_n338# a_n141_n424#
X0 a_15_n250# a_n33_n338# a_n73_n250# a_n141_n424# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.15
C0 a_n33_n338# a_n73_n250# 0.0337f
C1 a_n73_n250# a_15_n250# 0.401f
C2 a_n33_n338# a_15_n250# 0.0337f
C3 a_15_n250# a_n141_n424# 0.24f
C4 a_n73_n250# a_n141_n424# 0.24f
C5 a_n33_n338# a_n141_n424# 0.327f
.ends

.subckt th14 V14 Vin Vn m1_641_n318# Vp m1_891_419#
XXM0 Vn Vn m1_641_n318# Vp Vn sky130_fd_pr__pfet_01v8_HPNF99
XXM1 m1_641_n318# m1_891_419# Vin Vn sky130_fd_pr__nfet_01v8_JZU22M
XXM2 Vin Vp m1_891_419# Vp Vn sky130_fd_pr__pfet_01v8_TM5S5A
XXM3 Vp m1_891_419# V14 Vp Vn sky130_fd_pr__pfet_01v8_AM8GZ5
XXM4 Vn V14 m1_891_419# Vn sky130_fd_pr__nfet_01v8_H7HSAV
C0 m1_641_n318# m1_891_419# 0.00289f
C1 Vp m1_891_419# 0.227f
C2 V14 Vp 0.082f
C3 m1_641_n318# Vin 0.229f
C4 Vin Vp 0.201f
C5 V14 m1_891_419# 0.249f
C6 m1_641_n318# Vp 0.0629f
C7 Vin m1_891_419# 0.132f
C8 Vin V14 0.00516f
C9 V14 Vn 0.273f
C10 m1_891_419# Vn 1.7f
C11 Vp Vn 3.39f
C12 m1_641_n318# Vn 0.313f
C13 Vin Vn 1.76f
.ends

.subckt sky130_fd_pr__nfet_01v8_VGVEGU a_n142_n216# a_n74_n42# a_n33_n130# a_16_n42#
X0 a_16_n42# a_n33_n130# a_n74_n42# a_n142_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.16
C0 a_n33_n130# a_n74_n42# 0.0191f
C1 a_n33_n130# a_16_n42# 0.0191f
C2 a_n74_n42# a_16_n42# 0.0684f
C3 a_16_n42# a_n142_n216# 0.0652f
C4 a_n74_n42# a_n142_n216# 0.0652f
C5 a_n33_n130# a_n142_n216# 0.317f
.ends

.subckt sky130_fd_pr__pfet_01v8_EDPLE3 a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 w_n211_n261# a_n33_n139# 0.187f
C1 w_n211_n261# a_15_n42# 0.0197f
C2 w_n211_n261# a_n73_n42# 0.0197f
C3 a_n33_n139# a_15_n42# 0.0192f
C4 a_n33_n139# a_n73_n42# 0.0192f
C5 a_n73_n42# a_15_n42# 0.0699f
C6 a_15_n42# VSUBS 0.0445f
C7 a_n73_n42# VSUBS 0.0445f
C8 a_n33_n139# VSUBS 0.143f
C9 w_n211_n261# VSUBS 0.749f
.ends

.subckt sky130_fd_pr__pfet_01v8_JM8GTH a_50_n42# w_n246_n261# a_n50_n139# a_n108_n42#
+ VSUBS
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 w_n246_n261# a_n50_n139# 0.223f
C1 w_n246_n261# a_50_n42# 0.0224f
C2 w_n246_n261# a_n108_n42# 0.0224f
C3 a_n50_n139# a_50_n42# 0.00909f
C4 a_n50_n139# a_n108_n42# 0.00909f
C5 a_n108_n42# a_50_n42# 0.0391f
C6 a_50_n42# VSUBS 0.0488f
C7 a_n108_n42# VSUBS 0.0488f
C8 a_n50_n139# VSUBS 0.209f
C9 w_n246_n261# VSUBS 0.88f
.ends

.subckt sky130_fd_pr__nfet_01v8_MYA4RC a_n73_n46# a_n33_n134# a_15_n46# a_n175_n186#
X0 a_15_n46# a_n33_n134# a_n73_n46# a_n175_n186# sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.5 as=0.133 ps=1.5 w=0.46 l=0.15
C0 a_n33_n134# a_n73_n46# 0.0212f
C1 a_n33_n134# a_15_n46# 0.0212f
C2 a_n73_n46# a_15_n46# 0.0763f
C3 a_15_n46# a_n175_n186# 0.0671f
C4 a_n73_n46# a_n175_n186# 0.0756f
C5 a_n33_n134# a_n175_n186# 0.314f
.ends

.subckt th07 Vin V07 Vp m1_808_n892# Vn
XXM0 Vn m1_808_n892# Vin Vn sky130_fd_pr__nfet_01v8_VGVEGU
XXM1 m1_808_n892# Vp Vin Vp Vn sky130_fd_pr__pfet_01v8_EDPLE3
XXM2 V07 Vp m1_808_n892# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM3 V07 m1_808_n892# Vn Vn sky130_fd_pr__nfet_01v8_MYA4RC
C0 Vp V07 0.0569f
C1 Vin Vp 0.157f
C2 Vin V07 0.00135f
C3 m1_808_n892# Vp 0.209f
C4 m1_808_n892# V07 0.112f
C5 m1_808_n892# Vin 0.365f
C6 Vin Vn 0.524f
C7 Vp Vn 1.57f
C8 m1_808_n892# Vn 0.596f
C9 V07 Vn 0.276f
.ends

.subckt sky130_fd_pr__pfet_01v8_P28Q2U a_n33_n232# a_15_n135# w_n211_n354# a_n73_n135#
+ VSUBS
X0 a_15_n135# a_n33_n232# a_n73_n135# w_n211_n354# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.28 as=0.391 ps=3.28 w=1.35 l=0.15
C0 w_n211_n354# a_15_n135# 0.0279f
C1 w_n211_n354# a_n73_n135# 0.0279f
C2 a_n73_n135# a_15_n135# 0.218f
C3 w_n211_n354# a_n33_n232# 0.19f
C4 a_15_n135# a_n33_n232# 0.0258f
C5 a_n73_n135# a_n33_n232# 0.0258f
C6 a_15_n135# VSUBS 0.115f
C7 a_n73_n135# VSUBS 0.115f
C8 a_n33_n232# VSUBS 0.146f
C9 w_n211_n354# VSUBS 0.983f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZMY3VB a_n348_n42# a_n290_n130# a_n450_n182# a_290_n42#
X0 a_290_n42# a_n290_n130# a_n348_n42# a_n450_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.9
C0 a_n290_n130# a_290_n42# 0.0217f
C1 a_n290_n130# a_n348_n42# 0.0217f
C2 a_290_n42# a_n348_n42# 0.00961f
C3 a_290_n42# a_n450_n182# 0.076f
C4 a_n348_n42# a_n450_n182# 0.0839f
C5 a_n290_n130# a_n450_n182# 1.6f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 w_n211_n319# a_15_n100# 0.0248f
C1 w_n211_n319# a_n73_n100# 0.0248f
C2 a_n73_n100# a_15_n100# 0.162f
C3 w_n211_n319# a_n33_n197# 0.189f
C4 a_15_n100# a_n33_n197# 0.0236f
C5 a_n73_n100# a_n33_n197# 0.0236f
C6 a_15_n100# VSUBS 0.0885f
C7 a_n73_n100# VSUBS 0.0885f
C8 a_n33_n197# VSUBS 0.145f
C9 w_n211_n319# VSUBS 0.894f
.ends

.subckt sky130_fd_pr__pfet_01v8_WV9GCW a_n158_n42# w_n296_n261# a_n100_n139# a_100_n42#
+ VSUBS
X0 a_100_n42# a_n100_n139# a_n158_n42# w_n296_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1
C0 w_n296_n261# a_100_n42# 0.0224f
C1 w_n296_n261# a_n158_n42# 0.0224f
C2 a_n158_n42# a_100_n42# 0.024f
C3 w_n296_n261# a_n100_n139# 0.346f
C4 a_100_n42# a_n100_n139# 0.0144f
C5 a_n158_n42# a_n100_n139# 0.0144f
C6 a_100_n42# VSUBS 0.0504f
C7 a_n158_n42# VSUBS 0.0504f
C8 a_n100_n139# VSUBS 0.353f
C9 w_n296_n261# VSUBS 1.06f
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n141_240# a_n33_n188# a_15_n100#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n141_240# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n33_n188# a_15_n100# 0.0254f
C1 a_n33_n188# a_n73_n100# 0.0254f
C2 a_15_n100# a_n73_n100# 0.162f
C3 a_15_n100# a_n141_240# 0.113f
C4 a_n73_n100# a_n141_240# 0.113f
C5 a_n33_n188# a_n141_240# 0.322f
.ends

.subckt th12 Vp V12 Vin m1_394_n856# Vn m1_529_n42#
XXM0 Vn Vn Vp m1_394_n856# Vn sky130_fd_pr__pfet_01v8_P28Q2U
XXM1 m1_529_n42# Vin Vn m1_394_n856# sky130_fd_pr__nfet_01v8_ZMY3VB
XXM2 m1_529_n42# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM3 Vp Vp m1_529_n42# V12 Vn sky130_fd_pr__pfet_01v8_WV9GCW
XXM4 V12 Vn m1_529_n42# Vn sky130_fd_pr__nfet_01v8_648S5X
C0 Vp V12 0.0454f
C1 Vn V12 0.0234f
C2 Vin Vp 0.238f
C3 m1_529_n42# m1_394_n856# 0.0134f
C4 Vin Vn 0.135f
C5 Vp m1_529_n42# 0.322f
C6 Vn m1_529_n42# 0.254f
C7 Vin V12 0.00205f
C8 Vp m1_394_n856# 0.04f
C9 Vn m1_394_n856# 0.0338f
C10 V12 m1_529_n42# 0.0929f
C11 Vin m1_529_n42# 0.0965f
C12 Vp Vn 0.132f
C13 V12 m1_394_n856# 4.74e-19
C14 Vin m1_394_n856# 0.321f
C15 Vn 0 0.29f
C16 Vp 0 2.88f
C17 m1_529_n42# 0 0.861f
C18 V12 0 0.359f
C19 Vin 0 1.9f
C20 m1_394_n856# 0 0.215f
.ends

.subckt sky130_fd_pr__nfet_01v8_Q7AWK3 a_n180_n340# a_20_n200# a_n78_n200# a_n33_n288#
X0 a_20_n200# a_n33_n288# a_n78_n200# a_n180_n340# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
C0 a_n33_n288# a_n78_n200# 0.024f
C1 a_n33_n288# a_20_n200# 0.024f
C2 a_20_n200# a_n78_n200# 0.288f
C3 a_20_n200# a_n180_n340# 0.202f
C4 a_n78_n200# a_n180_n340# 0.237f
C5 a_n33_n288# a_n180_n340# 0.325f
.ends

.subckt sky130_fd_pr__pfet_01v8_EXJYQP w_n359_n261# a_n163_n139# a_n221_n42# a_163_n42#
+ VSUBS
X0 a_163_n42# a_n163_n139# a_n221_n42# w_n359_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.63
C0 a_163_n42# w_n359_n261# 0.0408f
C1 a_163_n42# a_n163_n139# 0.0182f
C2 a_163_n42# a_n221_n42# 0.0161f
C3 w_n359_n261# a_n163_n139# 0.413f
C4 w_n359_n261# a_n221_n42# 0.0179f
C5 a_n221_n42# a_n163_n139# 0.0182f
C6 a_163_n42# VSUBS 0.041f
C7 a_n221_n42# VSUBS 0.056f
C8 a_n163_n139# VSUBS 0.584f
C9 w_n359_n261# VSUBS 1.24f
.ends

.subckt sky130_fd_pr__pfet_01v8_HJHF6N a_n170_n50# w_n308_n269# a_n112_n147# a_112_n50#
+ VSUBS
X0 a_112_n50# a_n112_n147# a_n170_n50# w_n308_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1.12
C0 a_112_n50# w_n308_n269# 0.0232f
C1 a_112_n50# a_n112_n147# 0.0172f
C2 a_112_n50# a_n170_n50# 0.0259f
C3 w_n308_n269# a_n112_n147# 0.378f
C4 w_n308_n269# a_n170_n50# 0.0232f
C5 a_n170_n50# a_n112_n147# 0.0172f
C6 a_112_n50# VSUBS 0.0577f
C7 a_n170_n50# VSUBS 0.0577f
C8 a_n112_n147# VSUBS 0.389f
C9 w_n308_n269# VSUBS 1.14f
.ends

.subckt sky130_fd_pr__nfet_01v8_N39H2X a_n76_n100# a_n33_n188# a_18_n100# a_144_n240#
X0 a_18_n100# a_n33_n188# a_n76_n100# a_144_n240# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.18
C0 a_n33_n188# a_n76_n100# 0.0205f
C1 a_n33_n188# a_18_n100# 0.0205f
C2 a_18_n100# a_n76_n100# 0.152f
C3 a_18_n100# a_144_n240# 0.133f
C4 a_n76_n100# a_144_n240# 0.115f
C5 a_n33_n188# a_144_n240# 0.32f
.ends

.subckt th05 Vp V05 Vin m1_752_n794# Vn
XXM0 Vn m1_752_n794# Vn Vin sky130_fd_pr__nfet_01v8_Q7AWK3
XXM1 Vp Vin m1_752_n794# Vp Vn sky130_fd_pr__pfet_01v8_EXJYQP
XXM2 Vp Vp m1_752_n794# V05 Vn sky130_fd_pr__pfet_01v8_HJHF6N
XXM3 Vn m1_752_n794# V05 Vn sky130_fd_pr__nfet_01v8_N39H2X
C0 V05 Vp 0.0548f
C1 m1_752_n794# Vn 0.136f
C2 Vin Vn 0.041f
C3 m1_752_n794# V05 0.0855f
C4 Vin V05 0.00406f
C5 m1_752_n794# Vp 0.198f
C6 Vin Vp 0.139f
C7 V05 Vn 0.0364f
C8 m1_752_n794# Vin 0.2f
C9 Vp Vn 0.0115f
C10 m1_752_n794# 0 0.788f
C11 Vp 0 2.28f
C12 V05 0 0.314f
C13 Vin 0 0.905f
C14 Vn 0 0.547f
.ends

.subckt sky130_fd_pr__nfet_01v8_4L9AWD a_n206_n182# a_n46_n130# a_n104_n42# a_46_n42#
X0 a_46_n42# a_n46_n130# a_n104_n42# a_n206_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.46
C0 a_n46_n130# a_n104_n42# 0.00852f
C1 a_n104_n42# a_46_n42# 0.0412f
C2 a_n46_n130# a_46_n42# 0.00852f
C3 a_46_n42# a_n206_n182# 0.0705f
C4 a_n104_n42# a_n206_n182# 0.0784f
C5 a_n46_n130# a_n206_n182# 0.388f
.ends

.subckt sky130_fd_pr__pfet_01v8_EZD9Q7 w_n224_n261# a_28_n42# a_n33_n139# a_n86_n42#
+ VSUBS
X0 a_28_n42# a_n33_n139# a_n86_n42# w_n224_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.28
C0 w_n224_n261# a_n33_n139# 0.183f
C1 a_n33_n139# a_n86_n42# 0.00625f
C2 a_n33_n139# a_28_n42# 0.00625f
C3 w_n224_n261# a_n86_n42# 0.0224f
C4 w_n224_n261# a_28_n42# 0.0224f
C5 a_n86_n42# a_28_n42# 0.0541f
C6 a_28_n42# VSUBS 0.0479f
C7 a_n86_n42# VSUBS 0.0479f
C8 a_n33_n139# VSUBS 0.155f
C9 w_n224_n261# VSUBS 0.799f
.ends

.subckt sky130_fd_pr__pfet_01v8_M479BZ a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 w_n211_n261# a_n33_n139# 0.182f
C1 a_n33_n139# a_n73_n42# 0.0192f
C2 a_n33_n139# a_15_n42# 0.0192f
C3 w_n211_n261# a_n73_n42# 0.016f
C4 w_n211_n261# a_15_n42# 0.0389f
C5 a_n73_n42# a_15_n42# 0.0699f
C6 a_15_n42# VSUBS 0.0328f
C7 a_n73_n42# VSUBS 0.0478f
C8 a_n33_n139# VSUBS 0.145f
C9 w_n211_n261# VSUBS 0.785f
.ends

.subckt sky130_fd_pr__nfet_01v8_4BNSKG a_n144_n216# a_18_n42# a_n33_n130# a_n76_n42#
X0 a_18_n42# a_n33_n130# a_n76_n42# a_n144_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.18
C0 a_n33_n130# a_n76_n42# 0.0154f
C1 a_n76_n42# a_18_n42# 0.0655f
C2 a_n33_n130# a_18_n42# 0.0154f
C3 a_18_n42# a_n144_n216# 0.0668f
C4 a_n76_n42# a_n144_n216# 0.0668f
C5 a_n33_n130# a_n144_n216# 0.319f
.ends

.subckt th10 Vp V10 Vin Vn m1_502_n495# m1_536_174#
XXM0 m1_502_n495# Vn Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vn Vin m1_536_174# m1_502_n495# sky130_fd_pr__nfet_01v8_4L9AWD
XXM2 Vp m1_536_174# Vin Vp Vn sky130_fd_pr__pfet_01v8_EZD9Q7
XXM3 Vp Vp m1_536_174# V10 Vn sky130_fd_pr__pfet_01v8_M479BZ
XXM4 Vn V10 m1_536_174# Vn sky130_fd_pr__nfet_01v8_4BNSKG
C0 Vin Vn 0.114f
C1 m1_536_174# m1_502_n495# 0.00612f
C2 Vp m1_536_174# 0.172f
C3 Vp m1_502_n495# 0.0256f
C4 Vin V10 0.0187f
C5 m1_536_174# Vn 0.233f
C6 Vn m1_502_n495# 0.0348f
C7 Vp Vn 0.102f
C8 m1_536_174# V10 0.177f
C9 V10 m1_502_n495# 0.042f
C10 Vp V10 0.0702f
C11 Vn V10 0.0577f
C12 m1_536_174# Vin 0.0971f
C13 Vin m1_502_n495# 0.0207f
C14 Vp Vin 0.175f
C15 Vin 0 0.664f
C16 m1_536_174# 0 0.825f
C17 Vp 0 2.17f
C18 V10 0 0.249f
C19 Vn 0 0.463f
C20 m1_502_n495# 0 0.146f
.ends

.subckt sky130_fd_pr__nfet_01v8_X33H33 a_n73_n110# a_n175_n250# a_n33_n198# a_15_n110#
X0 a_15_n110# a_n33_n198# a_n73_n110# a_n175_n250# sky130_fd_pr__nfet_01v8 ad=0.319 pd=2.78 as=0.319 ps=2.78 w=1.1 l=0.15
C0 a_n73_n110# a_n33_n198# 0.0261f
C1 a_n33_n198# a_15_n110# 0.0261f
C2 a_n73_n110# a_15_n110# 0.178f
C3 a_15_n110# a_n175_n250# 0.121f
C4 a_n73_n110# a_n175_n250# 0.141f
C5 a_n33_n198# a_n175_n250# 0.32f
.ends

.subckt sky130_fd_pr__pfet_01v8_AMA9E4 a_n194_n44# a_n136_n141# w_n332_n263# a_136_n44#
+ VSUBS
X0 a_136_n44# a_n136_n141# a_n194_n44# w_n332_n263# sky130_fd_pr__pfet_01v8 ad=0.128 pd=1.46 as=0.128 ps=1.46 w=0.44 l=1.36
C0 a_n136_n141# w_n332_n263# 0.434f
C1 a_136_n44# a_n194_n44# 0.0196f
C2 w_n332_n263# a_n194_n44# 0.0226f
C3 a_n136_n141# a_n194_n44# 0.0174f
C4 a_136_n44# w_n332_n263# 0.0226f
C5 a_136_n44# a_n136_n141# 0.0174f
C6 a_136_n44# VSUBS 0.0532f
C7 a_n194_n44# VSUBS 0.0532f
C8 a_n136_n141# VSUBS 0.457f
C9 w_n332_n263# VSUBS 1.2f
.ends

.subckt sky130_fd_pr__pfet_01v8_8DZSNJ a_n74_n100# a_16_n100# w_n212_n319# a_n33_n197#
+ VSUBS
X0 a_16_n100# a_n33_n197# a_n74_n100# w_n212_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.16
C0 a_n33_n197# w_n212_n319# 0.189f
C1 a_16_n100# a_n74_n100# 0.159f
C2 w_n212_n319# a_n74_n100# 0.0252f
C3 a_n33_n197# a_n74_n100# 0.0223f
C4 a_16_n100# w_n212_n319# 0.0252f
C5 a_16_n100# a_n33_n197# 0.0223f
C6 a_16_n100# VSUBS 0.089f
C7 a_n74_n100# VSUBS 0.089f
C8 a_n33_n197# VSUBS 0.146f
C9 w_n212_n319# VSUBS 0.899f
.ends

.subckt th03 Vp V03 Vin m1_890_n844# m1_638_n591# Vn
XXM0 Vn Vn Vin m1_890_n844# sky130_fd_pr__nfet_01v8_X33H33
XXM1 m1_638_n591# Vin Vp m1_890_n844# Vn sky130_fd_pr__pfet_01v8_AMA9E4
XXM2 Vp Vn Vp m1_638_n591# sky130_fd_pr__nfet_01v8_LH5FDA
XXM3 Vp V03 Vp m1_890_n844# Vn sky130_fd_pr__pfet_01v8_8DZSNJ
XXM4 m1_890_n844# Vn Vn V03 sky130_fd_pr__nfet_01v8_LH5FDA
C0 Vp V03 0.0492f
C1 m1_638_n591# m1_890_n844# 0.0187f
C2 m1_638_n591# Vin 0.0439f
C3 Vn m1_890_n844# 0.183f
C4 Vp m1_638_n591# 0.169f
C5 Vn Vin 0.105f
C6 Vn V03 0.0337f
C7 Vp Vn 0.023f
C8 m1_890_n844# Vin 0.188f
C9 m1_890_n844# V03 0.129f
C10 Vp m1_890_n844# 0.459f
C11 Vn m1_638_n591# 0.0097f
C12 Vin V03 0.0036f
C13 Vp Vin 0.313f
C14 Vp 0 3.07f
C15 Vn 0 0.446f
C16 m1_890_n844# 0 1.05f
C17 V03 0 0.308f
C18 m1_638_n591# 0 0.224f
C19 Vin 0 0.924f
.ends

.subckt sky130_fd_pr__nfet_01v8_SHU4BF a_n73_n353# a_n141_493# a_15_n353# a_n33_n441#
X0 a_15_n353# a_n33_n441# a_n73_n353# a_n141_493# sky130_fd_pr__nfet_01v8 ad=1.02 pd=7.64 as=1.02 ps=7.64 w=3.53 l=0.15
C0 a_n33_n441# a_n73_n353# 0.0384f
C1 a_15_n353# a_n73_n353# 0.564f
C2 a_n33_n441# a_15_n353# 0.0384f
C3 a_15_n353# a_n141_493# 0.327f
C4 a_n73_n353# a_n141_493# 0.327f
C5 a_n33_n441# a_n141_493# 0.329f
.ends

.subckt sky130_fd_pr__pfet_01v8_HE9GT9 a_n408_n42# a_350_n42# w_n546_n261# a_n350_n139#
+ VSUBS
X0 a_350_n42# a_n350_n139# a_n408_n42# w_n546_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 w_n546_n261# a_350_n42# 0.0179f
C1 w_n546_n261# a_n350_n139# 0.756f
C2 a_n408_n42# a_350_n42# 0.00807f
C3 a_n408_n42# a_n350_n139# 0.0226f
C4 w_n546_n261# a_n408_n42# 0.0408f
C5 a_n350_n139# a_350_n42# 0.0226f
C6 a_350_n42# VSUBS 0.0587f
C7 a_n408_n42# VSUBS 0.0437f
C8 a_n350_n139# VSUBS 1.19f
C9 w_n546_n261# VSUBS 1.83f
.ends

.subckt sky130_fd_pr__nfet_01v8_LHD8GA a_n408_n42# a_350_n42# a_n350_n130# a_n510_n182#
X0 a_350_n42# a_n350_n130# a_n408_n42# a_n510_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 a_n350_n130# a_n408_n42# 0.0226f
C1 a_350_n42# a_n408_n42# 0.00807f
C2 a_n350_n130# a_350_n42# 0.0226f
C3 a_350_n42# a_n510_n182# 0.0766f
C4 a_n408_n42# a_n510_n182# 0.0845f
C5 a_n350_n130# a_n510_n182# 1.9f
.ends

.subckt th01 Vp Vin V01 m1_991_n1219# Vn m1_571_n501#
XXM0 Vn Vn m1_991_n1219# Vin sky130_fd_pr__nfet_01v8_SHU4BF
XXM1 m1_571_n501# m1_991_n1219# Vp Vin Vn sky130_fd_pr__pfet_01v8_HE9GT9
XXM2 Vp m1_571_n501# Vp Vn sky130_fd_pr__nfet_01v8_LHD8GA
XXM3 Vp Vp V01 m1_991_n1219# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_991_n1219# Vn V01 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 V01 Vp 0.0684f
C1 V01 m1_571_n501# 2.16e-20
C2 Vn Vin 0.0582f
C3 m1_991_n1219# Vp 0.423f
C4 m1_991_n1219# m1_571_n501# 0.0899f
C5 V01 m1_991_n1219# 0.0901f
C6 Vin Vp 0.354f
C7 Vn Vp 0.0233f
C8 Vin m1_571_n501# 0.274f
C9 Vn m1_571_n501# 2.57e-20
C10 V01 Vin 0.00412f
C11 Vn V01 0.0149f
C12 m1_991_n1219# Vin 0.208f
C13 Vn m1_991_n1219# 0.0569f
C14 Vp m1_571_n501# 0.32f
C15 Vn 0 0.633f
C16 V01 0 0.373f
C17 m1_991_n1219# 0 1.24f
C18 Vp 0 4.41f
C19 m1_571_n501# 0 0.194f
C20 Vin 0 1.87f
.ends

.subckt sky130_fd_pr__pfet_01v8_MWHFPY a_n73_n63# a_n33_n160# w_n211_n282# a_15_n63#
+ VSUBS
X0 a_15_n63# a_n33_n160# a_n73_n63# w_n211_n282# sky130_fd_pr__pfet_01v8 ad=0.183 pd=1.84 as=0.183 ps=1.84 w=0.63 l=0.15
C0 a_n33_n160# a_n73_n63# 0.021f
C1 w_n211_n282# a_15_n63# 0.0591f
C2 w_n211_n282# a_n33_n160# 0.237f
C3 a_n33_n160# a_15_n63# 0.021f
C4 w_n211_n282# a_n73_n63# 0.0591f
C5 a_n73_n63# a_15_n63# 0.103f
C6 a_15_n63# VSUBS 0.0348f
C7 a_n73_n63# VSUBS 0.0348f
C8 a_n33_n160# VSUBS 0.116f
C9 w_n211_n282# VSUBS 1.1f
.ends

.subckt sky130_fd_pr__nfet_01v8_DPSGWY a_350_n100# a_n408_n100# a_n350_n188# a_n510_n274#
X0 a_350_n100# a_n350_n188# a_n408_n100# a_n510_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3.5
C0 a_n408_n100# a_350_n100# 0.0188f
C1 a_n350_n188# a_n408_n100# 0.0439f
C2 a_n350_n188# a_350_n100# 0.0439f
C3 a_350_n100# a_n510_n274# 0.159f
C4 a_n408_n100# a_n510_n274# 0.159f
C5 a_n350_n188# a_n510_n274# 2.13f
.ends

.subckt preamp Vp Vin Vpamp Vn
XXM0 Vn Vin Vp Vpamp Vn sky130_fd_pr__pfet_01v8_MWHFPY
XXM1 Vpamp Vp Vin Vn sky130_fd_pr__nfet_01v8_DPSGWY
C0 Vpamp Vn 0.047f
C1 Vpamp Vp 0.0552f
C2 Vn Vp 0.297f
C3 Vin Vpamp 0.0777f
C4 Vin Vn 0.29f
C5 Vin Vp 0.324f
C6 Vn 0 0.193f
C7 Vpamp 0 0.444f
C8 Vp 0 1.53f
C9 Vin 0 2.21f
.ends

.subckt sky130_fd_pr__pfet_01v8_LDQF7K a_n33_n147# a_29_n50# a_n87_n50# w_n225_n269#
+ VSUBS
X0 a_29_n50# a_n33_n147# a_n87_n50# w_n225_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.29
C0 a_n33_n147# a_n87_n50# 0.00691f
C1 w_n225_n269# a_n33_n147# 0.176f
C2 a_29_n50# a_n87_n50# 0.0628f
C3 w_n225_n269# a_29_n50# 0.0186f
C4 w_n225_n269# a_n87_n50# 0.0457f
C5 a_n33_n147# a_29_n50# 0.00691f
C6 a_29_n50# VSUBS 0.0581f
C7 a_n87_n50# VSUBS 0.0403f
C8 a_n33_n147# VSUBS 0.158f
C9 w_n225_n269# VSUBS 0.854f
.ends

.subckt sky130_fd_pr__nfet_01v8_HZA4VB a_326_n230# a_n200_n130# a_200_n42# li_n360_158#
+ a_n258_n42#
X0 a_200_n42# a_n200_n130# a_n258_n42# a_326_n230# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_n258_n42# a_200_n42# 0.0134f
C1 a_n200_n130# a_n258_n42# 0.0196f
C2 a_n200_n130# a_200_n42# 0.0196f
C3 li_n360_158# a_326_n230# 0.0244f
C4 a_200_n42# a_326_n230# 0.0748f
C5 a_n258_n42# a_326_n230# 0.0746f
C6 a_n200_n130# a_326_n230# 1.15f
.ends

.subckt sky130_fd_pr__pfet_01v8_GEY2B5 w_n275_n270# a_n137_n51# a_79_n51# a_n79_n148#
+ VSUBS
X0 a_79_n51# a_n79_n148# a_n137_n51# w_n275_n270# sky130_fd_pr__pfet_01v8 ad=0.148 pd=1.6 as=0.148 ps=1.6 w=0.51 l=0.79
C0 a_n79_n148# a_n137_n51# 0.0141f
C1 w_n275_n270# a_n79_n148# 0.294f
C2 a_79_n51# a_n137_n51# 0.0345f
C3 w_n275_n270# a_79_n51# 0.0232f
C4 w_n275_n270# a_n137_n51# 0.0232f
C5 a_n79_n148# a_79_n51# 0.0141f
C6 a_79_n51# VSUBS 0.0573f
C7 a_n137_n51# VSUBS 0.0573f
C8 a_n79_n148# VSUBS 0.294f
C9 w_n275_n270# VSUBS 1.01f
.ends

.subckt sky130_fd_pr__pfet_01v8_KQKFM4 w_n526_n261# a_n330_n139# a_330_n42# a_n388_n42#
+ VSUBS
X0 a_330_n42# a_n330_n139# a_n388_n42# w_n526_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.3
C0 a_n330_n139# a_n388_n42# 0.0223f
C1 w_n526_n261# a_n330_n139# 0.911f
C2 a_330_n42# a_n388_n42# 0.00853f
C3 w_n526_n261# a_330_n42# 0.0224f
C4 w_n526_n261# a_n388_n42# 0.0224f
C5 a_n330_n139# a_330_n42# 0.0223f
C6 a_330_n42# VSUBS 0.0545f
C7 a_n388_n42# VSUBS 0.0545f
C8 a_n330_n139# VSUBS 1.02f
C9 w_n526_n261# VSUBS 1.89f
.ends

.subckt sky130_fd_pr__nfet_01v8_5NW376 a_n73_n251# a_n141_391# a_15_n251# a_n33_n339#
X0 a_15_n251# a_n33_n339# a_n73_n251# a_n141_391# sky130_fd_pr__nfet_01v8 ad=0.728 pd=5.6 as=0.728 ps=5.6 w=2.51 l=0.15
C0 a_n73_n251# a_15_n251# 0.402f
C1 a_n33_n339# a_n73_n251# 0.0337f
C2 a_n33_n339# a_15_n251# 0.0337f
C3 a_15_n251# a_n141_391# 0.241f
C4 a_n73_n251# a_n141_391# 0.241f
C5 a_n33_n339# a_n141_391# 0.327f
.ends

.subckt th15 V15 Vin m1_597_n912# Vp m1_849_n157# Vn
XXM0 Vn Vn m1_597_n912# Vp Vn sky130_fd_pr__pfet_01v8_LDQF7K
XXM1 Vn Vin m1_849_n157# Vn m1_597_n912# sky130_fd_pr__nfet_01v8_HZA4VB
XXM2 Vp Vp m1_849_n157# Vin Vn sky130_fd_pr__pfet_01v8_GEY2B5
XXM3 Vp m1_849_n157# V15 Vp Vn sky130_fd_pr__pfet_01v8_KQKFM4
XXM4 Vn Vn V15 m1_849_n157# sky130_fd_pr__nfet_01v8_5NW376
C0 m1_849_n157# V15 0.202f
C1 Vin m1_597_n912# 0.211f
C2 m1_849_n157# Vp 0.226f
C3 Vn V15 2.72e-19
C4 Vn Vp 0.0678f
C5 m1_849_n157# m1_597_n912# 0.00715f
C6 V15 Vp 0.0762f
C7 Vn m1_597_n912# 0.175f
C8 m1_597_n912# Vp 0.0557f
C9 m1_849_n157# Vin 0.0977f
C10 Vn Vin 0.38f
C11 V15 Vin 0.00573f
C12 Vin Vp 0.166f
C13 m1_849_n157# Vn 0.171f
C14 V15 0 0.332f
C15 Vn 0 0.276f
C16 m1_849_n157# 0 1.28f
C17 Vp 0 3.52f
C18 Vin 0 1.58f
C19 m1_597_n912# 0 0.19f
.ends

.subckt sky130_fd_pr__nfet_01v8_JSJ4VK a_113_n42# a_n239_n216# a_n171_n42# a_n113_n130#
X0 a_113_n42# a_n113_n130# a_n171_n42# a_n239_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.13
C0 a_n171_n42# a_113_n42# 0.0218f
C1 a_n113_n130# a_113_n42# 0.0154f
C2 a_n171_n42# a_n113_n130# 0.0154f
C3 a_113_n42# a_n239_n216# 0.0734f
C4 a_n171_n42# a_n239_n216# 0.0734f
C5 a_n113_n130# a_n239_n216# 0.746f
.ends

.subckt sky130_fd_pr__pfet_01v8_EVXEQ2 a_16_n67# a_n33_n164# a_n74_n67# w_n212_n286#
+ VSUBS
X0 a_16_n67# a_n33_n164# a_n74_n67# w_n212_n286# sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.92 as=0.194 ps=1.92 w=0.67 l=0.16
C0 a_16_n67# a_n74_n67# 0.107f
C1 a_16_n67# a_n33_n164# 0.0198f
C2 a_16_n67# w_n212_n286# 0.0544f
C3 a_n33_n164# a_n74_n67# 0.0198f
C4 w_n212_n286# a_n74_n67# 0.0184f
C5 a_n33_n164# w_n212_n286# 0.183f
C6 a_16_n67# VSUBS 0.0435f
C7 a_n74_n67# VSUBS 0.0673f
C8 a_n33_n164# VSUBS 0.147f
C9 w_n212_n286# VSUBS 0.864f
.ends

.subckt sky130_fd_pr__pfet_01v8_BBE9QE w_n244_n262# a_n106_n43# a_48_n43# a_n48_n140#
+ VSUBS
X0 a_48_n43# a_n48_n140# a_n106_n43# w_n244_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.48
C0 a_48_n43# a_n106_n43# 0.041f
C1 a_48_n43# a_n48_n140# 0.00893f
C2 a_48_n43# w_n244_n262# 0.0225f
C3 a_n48_n140# a_n106_n43# 0.00893f
C4 w_n244_n262# a_n106_n43# 0.0225f
C5 a_n48_n140# w_n244_n262# 0.218f
C6 a_48_n43# VSUBS 0.0495f
C7 a_n106_n43# VSUBS 0.0495f
C8 a_n48_n140# VSUBS 0.203f
C9 w_n244_n262# VSUBS 0.876f
.ends

.subckt sky130_fd_pr__nfet_01v8_NCP4B2 a_n73_n47# a_n141_n221# a_n33_n135# a_15_n47#
X0 a_15_n47# a_n33_n135# a_n73_n47# a_n141_n221# sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.52 as=0.136 ps=1.52 w=0.47 l=0.15
C0 a_n73_n47# a_15_n47# 0.0779f
C1 a_n33_n135# a_15_n47# 0.0213f
C2 a_n73_n47# a_n33_n135# 0.0213f
C3 a_15_n47# a_n141_n221# 0.0686f
C4 a_n73_n47# a_n141_n221# 0.0686f
C5 a_n33_n135# a_n141_n221# 0.317f
.ends

.subckt th08 Vin V08 m1_477_n803# Vp Vn
XXM0 Vn Vn m1_477_n803# Vin sky130_fd_pr__nfet_01v8_JSJ4VK
XXM1 Vp Vin m1_477_n803# Vp Vn sky130_fd_pr__pfet_01v8_EVXEQ2
XXM2 Vp Vp V08 m1_477_n803# Vn sky130_fd_pr__pfet_01v8_BBE9QE
XXM3 Vn Vn m1_477_n803# V08 sky130_fd_pr__nfet_01v8_NCP4B2
C0 Vin m1_477_n803# 0.356f
C1 V08 m1_477_n803# 0.108f
C2 Vin V08 0.00163f
C3 Vp m1_477_n803# 0.154f
C4 Vin Vp 0.0933f
C5 V08 Vp 0.0461f
C6 m1_477_n803# Vn 0.656f
C7 Vin Vn 1.02f
C8 V08 Vn 0.271f
C9 Vp Vn 1.66f
.ends

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X a_208_47# a_75_199#
+ a_544_297# a_315_47# a_201_297#
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_208_47# X 1.91e-19
C1 X A1 1.2e-19
C2 a_201_297# A1 0.011f
C3 VGND a_208_47# 0.00302f
C4 VGND A1 0.0113f
C5 X a_544_297# 2.35e-19
C6 VPWR a_208_47# 8.35e-19
C7 A3 A2 0.0747f
C8 a_201_297# a_544_297# 0.00702f
C9 VPWR A1 0.0151f
C10 B1 a_75_199# 0.102f
C11 X A2 3.01e-19
C12 VGND a_544_297# 0.00256f
C13 a_201_297# A2 0.0112f
C14 VPWR a_544_297# 0.0105f
C15 VGND A2 0.0119f
C16 a_75_199# A3 0.163f
C17 VPB A1 0.0306f
C18 VPWR A2 0.0174f
C19 X a_75_199# 0.0959f
C20 a_201_297# a_75_199# 0.16f
C21 VGND a_75_199# 0.362f
C22 VPWR a_75_199# 0.109f
C23 VPB A2 0.0376f
C24 VGND a_315_47# 0.00427f
C25 VPWR a_315_47# 0.00154f
C26 VPB a_75_199# 0.0486f
C27 a_208_47# A2 0.00102f
C28 A1 A2 0.0689f
C29 B1 C1 0.066f
C30 a_208_47# a_75_199# 0.0159f
C31 A1 a_75_199# 0.0696f
C32 C1 X 5.14e-20
C33 A1 a_315_47# 0.00313f
C34 a_75_199# a_544_297# 0.0176f
C35 a_201_297# C1 0.00243f
C36 a_75_199# A2 0.0621f
C37 VGND C1 0.0181f
C38 VPWR C1 0.0146f
C39 a_315_47# A2 0.00335f
C40 B1 X 7.79e-20
C41 a_201_297# B1 0.00594f
C42 VPB C1 0.0394f
C43 VGND B1 0.0171f
C44 a_75_199# a_315_47# 0.0202f
C45 B1 VPWR 0.0125f
C46 X A3 0.00317f
C47 a_201_297# A3 0.00642f
C48 a_201_297# X 0.0131f
C49 VGND A3 0.0161f
C50 C1 A1 3.21e-19
C51 VGND X 0.0609f
C52 VPWR A3 0.0181f
C53 B1 VPB 0.0292f
C54 VGND a_201_297# 0.00403f
C55 VPWR X 0.0676f
C56 a_201_297# VPWR 0.211f
C57 VGND VPWR 0.0735f
C58 VPB A3 0.0268f
C59 B1 A1 0.0716f
C60 VPB X 0.0107f
C61 a_201_297# VPB 0.00186f
C62 VGND VPB 0.00772f
C63 C1 a_75_199# 0.0628f
C64 B1 a_544_297# 1.13e-19
C65 a_208_47# A3 3.65e-19
C66 VPWR VPB 0.0749f
C67 VGND VNB 0.437f
C68 VPWR VNB 0.365f
C69 X VNB 0.0906f
C70 C1 VNB 0.148f
C71 B1 VNB 0.0947f
C72 A1 VNB 0.101f
C73 A2 VNB 0.11f
C74 A3 VNB 0.0908f
C75 VPB VNB 0.782f
C76 a_201_297# VNB 0.00345f
C77 a_75_199# VNB 0.205f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_181_47# a_109_47# a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_181_47# a_27_47# 0.00401f
C1 VPWR X 0.0766f
C2 B X 0.00111f
C3 VPWR a_109_47# 3.29e-19
C4 A a_27_47# 0.157f
C5 a_181_47# VGND 0.00261f
C6 C VPB 0.0347f
C7 VPB a_27_47# 0.0501f
C8 VPWR C 0.00464f
C9 VPWR a_27_47# 0.145f
C10 VGND A 0.0154f
C11 B C 0.0746f
C12 B a_27_47# 0.0625f
C13 VPB VGND 0.00604f
C14 VPWR VGND 0.0475f
C15 B VGND 0.00714f
C16 C X 0.0149f
C17 X a_27_47# 0.087f
C18 a_109_47# a_27_47# 0.00517f
C19 X VGND 0.0708f
C20 a_109_47# VGND 0.00123f
C21 C a_27_47# 0.186f
C22 C VGND 0.0703f
C23 VGND a_27_47# 0.134f
C24 VPWR a_181_47# 3.97e-19
C25 VPB A 0.0426f
C26 VPWR A 0.0185f
C27 VPWR VPB 0.0795f
C28 B A 0.0869f
C29 B VPB 0.0836f
C30 VPWR B 0.128f
C31 X VPB 0.0121f
C32 a_109_47# A 6.45e-19
C33 a_181_47# C 0.00151f
C34 VGND VNB 0.3f
C35 X VNB 0.0923f
C36 C VNB 0.12f
C37 A VNB 0.174f
C38 VPWR VNB 0.274f
C39 B VNB 0.102f
C40 VPB VNB 0.516f
C41 a_27_47# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
C0 VPWR VGND 0.353f
C1 VPB VGND 0.0797f
C2 VPWR VPB 0.0625f
C3 VPWR VNB 0.47f
C4 VGND VNB 0.427f
C5 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VPWR VGND 0.546f
C1 VPB VGND 0.116f
C2 VPWR VPB 0.0787f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_384_47# a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
C0 VGND X 0.0512f
C1 VPB A2 0.0373f
C2 A1 A2 0.0921f
C3 a_81_21# A2 7.47e-19
C4 VGND a_384_47# 0.00366f
C5 VGND B1 0.0181f
C6 a_299_297# VPWR 0.202f
C7 a_299_297# VPB 0.0111f
C8 a_299_297# A1 0.0585f
C9 a_81_21# a_299_297# 0.0821f
C10 VPWR VPB 0.068f
C11 VPWR A1 0.0209f
C12 a_81_21# VPWR 0.146f
C13 VPWR X 0.0847f
C14 VPB A1 0.0264f
C15 a_299_297# a_384_47# 1.48e-19
C16 a_81_21# VPB 0.0593f
C17 a_81_21# A1 0.0568f
C18 VPB X 0.0108f
C19 VPWR a_384_47# 4.08e-19
C20 a_299_297# B1 0.00863f
C21 a_81_21# X 0.112f
C22 VPWR B1 0.0196f
C23 a_384_47# A1 0.00884f
C24 a_81_21# a_384_47# 0.00138f
C25 A1 B1 0.0817f
C26 VPB B1 0.0387f
C27 VGND A2 0.0495f
C28 a_81_21# B1 0.148f
C29 B1 X 3.04e-20
C30 VGND a_299_297# 0.00772f
C31 VGND VPWR 0.0579f
C32 a_299_297# A2 0.0468f
C33 VGND VPB 0.00713f
C34 VGND A1 0.0786f
C35 VPWR A2 0.0201f
C36 VGND a_81_21# 0.173f
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15 M=2
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15 M=2
C0 Y VPB 0.0061f
C1 VGND VPB 0.00649f
C2 A VPWR 0.0631f
C3 VPWR Y 0.209f
C4 VGND VPWR 0.0423f
C5 A Y 0.0894f
C6 A VGND 0.0638f
C7 VPWR VPB 0.0521f
C8 VGND Y 0.155f
C9 A VPB 0.0742f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X a_29_53# a_183_297# a_111_297#
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 a_183_297# a_29_53# 0.00868f
C1 B X 6.52e-19
C2 VPWR X 0.0885f
C3 A C 0.0343f
C4 C a_29_53# 0.0857f
C5 VPWR a_111_297# 5.94e-19
C6 a_183_297# VGND 5.75e-19
C7 A VPB 0.0377f
C8 VPB a_29_53# 0.0491f
C9 B A 0.0787f
C10 B a_29_53# 0.121f
C11 VGND C 0.0161f
C12 VPWR A 0.00936f
C13 VPWR a_29_53# 0.0833f
C14 VPB VGND 0.00724f
C15 B VGND 0.0152f
C16 VPWR VGND 0.0459f
C17 A X 0.00127f
C18 X a_29_53# 0.0991f
C19 A a_111_297# 0.00223f
C20 a_111_297# a_29_53# 0.005f
C21 X VGND 0.036f
C22 a_111_297# VGND 3.96e-19
C23 A a_29_53# 0.242f
C24 A VGND 0.0187f
C25 VGND a_29_53# 0.217f
C26 a_183_297# VPWR 8.13e-19
C27 VPB C 0.0396f
C28 B C 0.0802f
C29 B VPB 0.0962f
C30 VPWR C 0.00457f
C31 VPWR VPB 0.0649f
C32 B VPWR 0.147f
C33 X VPB 0.0109f
C34 a_183_297# A 0.00239f
C35 VGND VNB 0.306f
C36 X VNB 0.0882f
C37 A VNB 0.117f
C38 C VNB 0.16f
C39 B VNB 0.117f
C40 VPWR VNB 0.253f
C41 VPB VNB 0.516f
C42 a_29_53# VNB 0.18f
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
C0 VPWR VGND 0.903f
C1 VPB VGND 0.161f
C2 VPWR VPB 0.0858f
C3 VPWR VNB 0.867f
C4 VGND VNB 0.761f
C5 VPB VNB 0.605f
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 A VGND 0.0486f
C1 VPWR VGND 0.0314f
C2 a_109_297# VGND 0.00128f
C3 B A 0.0584f
C4 B VPWR 0.0148f
C5 VPB VGND 0.00456f
C6 B VPB 0.0367f
C7 Y VGND 0.154f
C8 B Y 0.0877f
C9 A VPWR 0.0528f
C10 a_109_297# VPWR 0.00638f
C11 VPB A 0.0415f
C12 VPB VPWR 0.0449f
C13 A Y 0.0471f
C14 VPWR Y 0.0995f
C15 a_109_297# Y 0.0113f
C16 VPB Y 0.0139f
C17 B VGND 0.0451f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X a_193_297# a_465_47#
+ a_205_47# a_109_297# a_27_47#
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
C0 a_193_297# a_27_47# 0.144f
C1 VPB B1 0.0321f
C2 VPWR C1 0.0139f
C3 VGND C1 0.0196f
C4 VPB a_109_297# 0.00421f
C5 a_465_47# VPWR 5.05e-19
C6 a_465_47# VGND 0.00257f
C7 B2 C1 0.0726f
C8 C1 a_27_47# 0.0792f
C9 A2 VPWR 0.0209f
C10 A2 VGND 0.0168f
C11 a_193_297# A1 0.0109f
C12 a_465_47# a_27_47# 0.013f
C13 VPB VPWR 0.0799f
C14 VPB VGND 0.00844f
C15 A2 a_27_47# 0.153f
C16 a_193_297# X 0.00367f
C17 VPB B2 0.0256f
C18 VPB a_27_47# 0.0512f
C19 A1 C1 1.77e-20
C20 a_465_47# A1 7.06e-19
C21 A2 A1 0.0692f
C22 B1 a_109_297# 0.00736f
C23 X C1 5.03e-20
C24 VPB A1 0.0343f
C25 a_465_47# X 1.56e-19
C26 A2 X 0.00157f
C27 B1 VPWR 0.00982f
C28 B1 VGND 0.0133f
C29 VPB X 0.0113f
C30 B2 B1 0.0784f
C31 B1 a_27_47# 0.112f
C32 a_109_297# VPWR 0.15f
C33 a_109_297# VGND 0.00284f
C34 B2 a_109_297# 0.0133f
C35 a_109_297# a_27_47# 0.0961f
C36 VPWR VGND 0.0722f
C37 B1 A1 0.0609f
C38 B2 VPWR 0.00842f
C39 B2 VGND 0.0174f
C40 VPWR a_27_47# 0.099f
C41 VGND a_27_47# 0.395f
C42 a_109_297# A1 1.05e-19
C43 B2 a_27_47# 0.0959f
C44 B1 X 9.58e-20
C45 a_109_297# X 3.99e-19
C46 A1 VPWR 0.0161f
C47 A1 VGND 0.0126f
C48 A1 a_27_47# 0.0984f
C49 VPWR X 0.0897f
C50 VGND X 0.061f
C51 B2 X 6.77e-20
C52 X a_27_47# 0.0921f
C53 A2 a_193_297# 0.00683f
C54 VPB a_193_297# 0.00774f
C55 A1 X 2.77e-19
C56 A2 C1 9.03e-21
C57 VPB C1 0.0367f
C58 VPB A2 0.027f
C59 a_205_47# VPWR 1.62e-19
C60 a_205_47# VGND 0.00156f
C61 a_193_297# B1 0.00869f
C62 a_205_47# a_27_47# 0.00762f
C63 a_193_297# a_109_297# 0.0927f
C64 B1 C1 6.46e-19
C65 a_193_297# VPWR 0.169f
C66 a_193_297# VGND 0.00438f
C67 a_109_297# C1 0.00739f
C68 a_193_297# B2 0.00126f
C69 VGND VNB 0.437f
C70 X VNB 0.0919f
C71 VPWR VNB 0.364f
C72 A2 VNB 0.0896f
C73 A1 VNB 0.106f
C74 B1 VNB 0.108f
C75 B2 VNB 0.0887f
C76 C1 VNB 0.139f
C77 VPB VNB 0.782f
C78 a_193_297# VNB 0.0011f
C79 a_109_297# VNB 7.11e-19
C80 a_27_47# VNB 0.216f
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X a_256_47# a_584_47#
+ a_93_21# a_250_297# a_346_47#
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
C0 B1 A2 1.44e-20
C1 VGND a_250_297# 0.0072f
C2 X A1 6.03e-20
C3 a_346_47# A1 0.00465f
C4 VPWR a_250_297# 0.313f
C5 VPB A3 0.0291f
C6 VGND A1 0.0133f
C7 X VPB 0.0108f
C8 a_93_21# A3 0.124f
C9 A3 A2 0.0788f
C10 VPWR A1 0.016f
C11 B1 a_256_47# 2.07e-20
C12 a_93_21# X 0.0841f
C13 X A2 1.19e-19
C14 a_346_47# a_93_21# 0.0119f
C15 VGND VPB 0.00788f
C16 VGND a_584_47# 0.00683f
C17 a_346_47# A2 0.00252f
C18 VPWR a_584_47# 9.47e-19
C19 VPWR VPB 0.0756f
C20 VGND a_93_21# 0.251f
C21 VGND A2 0.0114f
C22 a_256_47# A3 4.42e-19
C23 VPWR a_93_21# 0.0907f
C24 VPWR A2 0.0133f
C25 a_250_297# A1 0.0129f
C26 VGND a_256_47# 0.00394f
C27 VPWR a_256_47# 9.47e-19
C28 a_250_297# a_584_47# 2.43e-19
C29 a_250_297# VPB 0.00616f
C30 a_93_21# a_250_297# 0.188f
C31 a_250_297# A2 0.0129f
C32 A1 VPB 0.0296f
C33 a_93_21# A1 0.0641f
C34 A1 A2 0.0971f
C35 B1 B2 0.0823f
C36 a_93_21# a_584_47# 0.00278f
C37 a_93_21# VPB 0.0485f
C38 VPB A2 0.0287f
C39 a_93_21# A2 0.0747f
C40 B2 A3 9.12e-20
C41 a_93_21# a_256_47# 0.0114f
C42 a_256_47# A2 0.00256f
C43 VGND B2 0.0469f
C44 VPWR B2 0.0108f
C45 B1 A3 7.88e-22
C46 B1 X 3.83e-20
C47 a_346_47# B1 5.39e-20
C48 VGND B1 0.0344f
C49 B1 VPWR 0.01f
C50 X A3 2.45e-19
C51 a_250_297# B2 0.0344f
C52 VGND A3 0.00974f
C53 B2 A1 3.14e-19
C54 VGND X 0.06f
C55 VPWR A3 0.0158f
C56 VGND a_346_47# 0.00514f
C57 VPWR X 0.0849f
C58 a_346_47# VPWR 0.00109f
C59 B2 VPB 0.0355f
C60 B1 a_250_297# 0.0125f
C61 a_93_21# B2 0.0147f
C62 VGND VPWR 0.076f
C63 B2 A2 1.46e-19
C64 B1 A1 0.0965f
C65 a_250_297# A3 0.00602f
C66 a_250_297# X 5.42e-19
C67 B1 a_584_47# 0.00143f
C68 B1 VPB 0.0276f
C69 B1 a_93_21# 0.0774f
C70 VGND VNB 0.465f
C71 VPWR VNB 0.365f
C72 X VNB 0.0937f
C73 B2 VNB 0.14f
C74 B1 VNB 0.101f
C75 A1 VNB 0.0951f
C76 A2 VNB 0.0921f
C77 A3 VNB 0.0929f
C78 VPB VNB 0.782f
C79 a_250_297# VNB 0.0278f
C80 a_93_21# VNB 0.151f
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X a_277_297# a_205_297# a_27_297#
+ a_109_297#
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 a_205_297# a_27_297# 0.00412f
C1 VPWR C 0.00723f
C2 VPB C 0.0338f
C3 VGND B 0.0159f
C4 VPWR a_109_297# 9.23e-19
C5 D B 0.00287f
C6 B a_27_297# 0.159f
C7 X VGND 0.0354f
C8 VPWR VGND 0.0546f
C9 X a_27_297# 0.0991f
C10 VPB VGND 0.00796f
C11 VPWR D 0.00503f
C12 VPWR a_27_297# 0.084f
C13 A B 0.0639f
C14 VPB D 0.0405f
C15 VPB a_27_297# 0.0517f
C16 X A 0.00133f
C17 C a_109_297# 0.00356f
C18 VPWR A 0.00769f
C19 VPB A 0.033f
C20 C VGND 0.0191f
C21 D C 0.0954f
C22 C a_27_297# 0.158f
C23 a_109_297# VGND 7.58e-19
C24 a_109_297# a_27_297# 0.00695f
C25 C A 0.028f
C26 D VGND 0.0517f
C27 VGND a_27_297# 0.235f
C28 D a_27_297# 0.054f
C29 a_277_297# B 2.29e-19
C30 A VGND 0.016f
C31 X a_277_297# 6.43e-20
C32 D A 2.13e-19
C33 VPWR a_277_297# 7.48e-19
C34 A a_27_297# 0.163f
C35 VPWR a_205_297# 5.16e-19
C36 C a_277_297# 5.54e-19
C37 X B 6.42e-19
C38 VPWR B 0.193f
C39 VPB B 0.106f
C40 VPWR X 0.0878f
C41 X VPB 0.0109f
C42 a_277_297# VGND 4.65e-19
C43 a_205_297# C 0.00261f
C44 VPWR VPB 0.075f
C45 a_277_297# a_27_297# 0.00876f
C46 C B 0.0917f
C47 a_277_297# A 2.28e-19
C48 a_205_297# VGND 3.36e-19
C49 VGND VNB 0.367f
C50 X VNB 0.0883f
C51 A VNB 0.109f
C52 C VNB 0.105f
C53 D VNB 0.175f
C54 B VNB 0.115f
C55 VPWR VNB 0.29f
C56 VPB VNB 0.605f
C57 a_27_297# VNB 0.163f
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
C0 VPWR VGND 1.57f
C1 VPB VGND 0.35f
C2 VPWR VPB 0.137f
C3 VPWR VNB 1.67f
C4 VGND VNB 1.47f
C5 VPB VNB 1.14f
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X a_369_47# a_469_47#
+ a_297_47# a_193_413# a_27_47#
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
C0 X C 0.00479f
C1 a_369_47# C 0.00448f
C2 VGND a_193_413# 0.0915f
C3 VPB A_N 0.0832f
C4 X a_469_47# 0.001f
C5 X VPB 0.0108f
C6 a_27_47# A_N 0.237f
C7 VGND C 0.0395f
C8 a_369_47# B 0.00129f
C9 VGND a_469_47# 0.00551f
C10 VGND VPB 0.0123f
C11 VGND a_27_47# 0.103f
C12 VGND B 0.037f
C13 a_193_413# C 0.0389f
C14 VGND a_297_47# 0.00183f
C15 a_193_413# a_469_47# 0.00109f
C16 a_193_413# VPB 0.0644f
C17 a_27_47# a_193_413# 0.125f
C18 a_193_413# B 0.144f
C19 C a_469_47# 0.00202f
C20 C VPB 0.0742f
C21 C B 0.164f
C22 D VPWR 0.0186f
C23 a_193_413# a_297_47# 0.00137f
C24 a_27_47# VPB 0.092f
C25 VPB B 0.089f
C26 a_27_47# B 0.0794f
C27 VPWR A_N 0.02f
C28 VPWR X 0.0586f
C29 a_369_47# VPWR 6.65e-19
C30 a_297_47# B 0.00353f
C31 VGND VPWR 0.0727f
C32 D X 0.0168f
C33 D VGND 0.0372f
C34 a_193_413# VPWR 0.281f
C35 VPWR C 0.0182f
C36 VGND A_N 0.0205f
C37 VGND X 0.0588f
C38 a_369_47# VGND 0.00505f
C39 VPWR a_469_47# 7.77e-19
C40 VPWR VPB 0.0818f
C41 D a_193_413# 0.155f
C42 a_27_47# VPWR 0.106f
C43 VPWR B 0.0186f
C44 D C 0.183f
C45 a_193_413# A_N 0.00151f
C46 a_193_413# X 0.108f
C47 D a_469_47# 0.00183f
C48 VPWR a_297_47# 2.82e-19
C49 D VPB 0.0763f
C50 a_369_47# a_193_413# 0.00181f
C51 VGND VNB 0.456f
C52 X VNB 0.0934f
C53 VPWR VNB 0.368f
C54 D VNB 0.123f
C55 C VNB 0.108f
C56 B VNB 0.12f
C57 A_N VNB 0.198f
C58 VPB VNB 0.782f
C59 a_193_413# VNB 0.136f
C60 a_27_47# VNB 0.224f
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X a_109_93# a_368_53# a_209_311#
+ a_296_53#
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
C0 a_296_53# a_109_93# 1.84e-19
C1 A_N C 7.6e-19
C2 VGND a_209_311# 0.131f
C3 VPB C 0.0339f
C4 A_N a_209_311# 0.00515f
C5 B VPWR 0.131f
C6 VPWR a_109_93# 0.0984f
C7 VPB a_209_311# 0.0515f
C8 VGND B 0.00796f
C9 VGND a_109_93# 0.0784f
C10 A_N B 2.03e-19
C11 A_N a_109_93# 0.117f
C12 X VPWR 0.0732f
C13 VPB B 0.0914f
C14 VPB a_109_93# 0.0652f
C15 VGND X 0.0647f
C16 C a_209_311# 0.19f
C17 A_N X 1.44e-19
C18 VPB X 0.0119f
C19 B C 0.0671f
C20 C a_109_93# 3.91e-20
C21 B a_209_311# 0.0609f
C22 a_209_311# a_109_93# 0.168f
C23 C X 0.0176f
C24 a_209_311# X 0.0877f
C25 B a_109_93# 0.0802f
C26 a_368_53# VPWR 4.26e-19
C27 VGND a_368_53# 0.0031f
C28 B X 0.00119f
C29 a_296_53# VPWR 1.15e-19
C30 VGND a_296_53# 6.07e-19
C31 C a_368_53# 0.00415f
C32 VGND VPWR 0.0657f
C33 A_N VPWR 0.0513f
C34 a_368_53# a_209_311# 0.0026f
C35 VPB VPWR 0.104f
C36 A_N VGND 0.045f
C37 VGND VPB 0.00909f
C38 A_N VPB 0.111f
C39 a_296_53# a_209_311# 0.0049f
C40 C VPWR 0.005f
C41 VGND C 0.0678f
C42 a_209_311# VPWR 0.155f
C43 VGND VNB 0.44f
C44 X VNB 0.0925f
C45 C VNB 0.114f
C46 B VNB 0.101f
C47 VPWR VNB 0.342f
C48 A_N VNB 0.197f
C49 VPB VNB 0.693f
C50 a_209_311# VNB 0.143f
C51 a_109_93# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15 M=4
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=4
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
C0 A VPWR 0.022f
C1 A VGND 0.0431f
C2 A a_27_47# 0.195f
C3 A VPB 0.0321f
C4 A X 0.014f
C5 VPWR VGND 0.057f
C6 a_27_47# VPWR 0.219f
C7 a_27_47# VGND 0.148f
C8 VPB VPWR 0.0632f
C9 VPB VGND 0.00583f
C10 a_27_47# VPB 0.139f
C11 VPWR X 0.317f
C12 VGND X 0.216f
C13 a_27_47# X 0.328f
C14 VPB X 0.0122f
C15 VGND VNB 0.358f
C16 X VNB 0.067f
C17 VPWR VNB 0.308f
C18 A VNB 0.148f
C19 VPB VNB 0.605f
C20 a_27_47# VNB 0.543f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
C0 VPWR X 0.111f
C1 B X 0.00276f
C2 a_59_75# X 0.109f
C3 X VGND 0.0993f
C4 VPB VPWR 0.0729f
C5 VPB B 0.0629f
C6 VPB a_59_75# 0.0563f
C7 VPB VGND 0.008f
C8 A X 1.68e-19
C9 VPB A 0.0806f
C10 a_145_75# VPWR 6.31e-19
C11 a_59_75# a_145_75# 0.00658f
C12 a_145_75# VGND 0.00468f
C13 VPWR B 0.0117f
C14 a_59_75# VPWR 0.15f
C15 a_59_75# B 0.143f
C16 VPWR VGND 0.0461f
C17 B VGND 0.0115f
C18 a_59_75# VGND 0.116f
C19 VPWR A 0.0362f
C20 B A 0.0971f
C21 a_59_75# A 0.0809f
C22 A VGND 0.0147f
C23 VPB X 0.0127f
C24 a_145_75# X 5.76e-19
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y a_297_297# a_191_297#
+ a_109_297#
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
C0 C Y 0.125f
C1 VGND a_191_297# 9.29e-19
C2 D Y 0.108f
C3 C a_191_297# 0.0195f
C4 A B 0.11f
C5 a_297_297# VPWR 0.00317f
C6 A VPB 0.041f
C7 VGND A 0.0526f
C8 VGND a_109_297# 0.00181f
C9 C A 0.00268f
C10 C a_109_297# 0.0062f
C11 VPWR B 0.0887f
C12 VPB VPWR 0.0524f
C13 VGND VPWR 0.0492f
C14 Y a_191_297# 0.00142f
C15 C VPWR 0.0509f
C16 D VPWR 0.0128f
C17 A Y 0.0175f
C18 Y a_109_297# 0.0122f
C19 Y VPWR 0.0561f
C20 a_191_297# VPWR 0.0049f
C21 A VPWR 0.0483f
C22 VPWR a_109_297# 0.00576f
C23 a_297_297# B 0.0132f
C24 VGND a_297_297# 8.1e-19
C25 VPB B 0.0304f
C26 VGND B 0.0191f
C27 VGND VPB 0.0048f
C28 C B 0.173f
C29 C VPB 0.0299f
C30 C VGND 0.0184f
C31 D VPB 0.0376f
C32 VGND D 0.0456f
C33 a_297_297# Y 1.24e-19
C34 C D 0.0523f
C35 Y B 0.0403f
C36 Y VPB 0.0127f
C37 VGND Y 0.151f
C38 a_191_297# B 0.00223f
C39 a_297_297# A 3.16e-19
C40 VGND VNB 0.322f
C41 VPWR VNB 0.276f
C42 Y VNB 0.0645f
C43 A VNB 0.174f
C44 B VNB 0.0968f
C45 C VNB 0.0911f
C46 D VNB 0.159f
C47 VPB VNB 0.516f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X a_75_212#
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 A X 8.48e-19
C1 A VGND 0.0184f
C2 A a_75_212# 0.178f
C3 A VPB 0.0525f
C4 A VPWR 0.0217f
C5 X VGND 0.0545f
C6 a_75_212# X 0.107f
C7 a_75_212# VGND 0.105f
C8 VPB X 0.0128f
C9 VPB VGND 0.00507f
C10 a_75_212# VPB 0.0571f
C11 X VPWR 0.0896f
C12 VGND VPWR 0.0289f
C13 a_75_212# VPWR 0.134f
C14 VPB VPWR 0.0355f
C15 VGND VNB 0.207f
C16 VPWR VNB 0.176f
C17 X VNB 0.0942f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_75_212# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 A VPWR 0.0215f
C1 A VGND 0.0184f
C2 A a_27_47# 0.181f
C3 A VPB 0.0524f
C4 A X 8.48e-19
C5 VPWR VGND 0.029f
C6 a_27_47# VPWR 0.135f
C7 a_27_47# VGND 0.105f
C8 VPB VPWR 0.0355f
C9 VPB VGND 0.00505f
C10 a_27_47# VPB 0.0592f
C11 VPWR X 0.0897f
C12 VGND X 0.0546f
C13 a_27_47# X 0.107f
C14 VPB X 0.0128f
C15 VGND VNB 0.207f
C16 X VNB 0.0941f
C17 VPWR VNB 0.175f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_27_47# VNB 0.208f
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X a_664_47# a_841_47#
+ a_381_47# a_62_47# a_558_47#
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VGND X 0.106f
C1 a_664_47# VPWR 0.131f
C2 VPB A 0.105f
C3 a_62_47# A 0.244f
C4 A X 0.0142f
C5 a_664_47# a_841_47# 0.134f
C6 a_664_47# VPB 0.043f
C7 VGND a_558_47# 0.0816f
C8 a_664_47# X 6.67e-19
C9 a_664_47# a_558_47# 0.314f
C10 a_381_47# VPWR 0.134f
C11 a_381_47# VPB 0.0447f
C12 a_381_47# X 0.318f
C13 VPWR a_841_47# 0.0614f
C14 VPWR VPB 0.103f
C15 a_62_47# VPWR 0.149f
C16 VPWR X 0.108f
C17 a_841_47# VPB 0.0108f
C18 a_381_47# a_558_47# 0.16f
C19 a_62_47# VPB 0.0515f
C20 VPB X 0.126f
C21 VPWR a_558_47# 0.084f
C22 a_62_47# X 0.156f
C23 a_558_47# a_841_47# 0.00368f
C24 a_558_47# VPB 0.115f
C25 a_558_47# X 0.0144f
C26 VGND A 0.0176f
C27 a_664_47# VGND 0.125f
C28 VGND a_381_47# 0.125f
C29 VGND VPWR 0.0902f
C30 a_381_47# A 5.42e-19
C31 VGND a_841_47# 0.0585f
C32 VGND VPB 0.008f
C33 VPWR A 0.0174f
C34 VGND a_62_47# 0.144f
C35 VGND VNB 0.537f
C36 VPWR VNB 0.439f
C37 X VNB 0.163f
C38 A VNB 0.198f
C39 VPB VNB 0.959f
C40 a_841_47# VNB 0.0929f
C41 a_664_47# VNB 0.13f
C42 a_558_47# VNB 0.164f
C43 a_381_47# VNB 0.11f
C44 a_62_47# VNB 0.169f
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y a_129_47# a_47_47# a_285_47#
+ a_377_297#
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 a_129_47# a_47_47# 0.00369f
C1 B Y 0.00334f
C2 VPB Y 0.00878f
C3 B a_377_297# 0.00254f
C4 VPWR A 0.0349f
C5 A a_47_47# 0.0307f
C6 a_129_47# VGND 0.00547f
C7 B VPWR 0.0408f
C8 B a_47_47# 0.356f
C9 VGND A 0.0635f
C10 VPB VPWR 0.0718f
C11 VPB a_47_47# 0.0444f
C12 Y a_377_297# 0.00188f
C13 B VGND 0.0389f
C14 VPB VGND 0.00568f
C15 VPWR Y 0.107f
C16 Y a_47_47# 0.143f
C17 VPWR a_377_297# 0.00559f
C18 a_377_297# a_47_47# 0.00899f
C19 Y VGND 0.0381f
C20 a_377_297# VGND 0.00125f
C21 VPWR a_47_47# 0.273f
C22 a_285_47# A 0.0353f
C23 VPWR VGND 0.0665f
C24 VGND a_47_47# 0.104f
C25 B a_285_47# 0.067f
C26 VPB a_285_47# 5.53e-19
C27 B a_129_47# 0.00236f
C28 Y a_285_47# 0.0439f
C29 B A 0.236f
C30 VPB A 0.0822f
C31 VPWR a_285_47# 0.00255f
C32 B VPB 0.0643f
C33 a_285_47# a_47_47# 0.0175f
C34 Y A 0.00181f
C35 a_285_47# VGND 0.211f
C36 a_129_47# VPWR 9.47e-19
C37 VGND VNB 0.4f
C38 Y VNB 0.0783f
C39 VPWR VNB 0.352f
C40 A VNB 0.217f
C41 B VNB 0.212f
C42 VPB VNB 0.693f
C43 a_285_47# VNB 0.0174f
C44 a_47_47# VNB 0.199f
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X a_472_297# a_80_21#
+ a_300_47# a_217_297#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
C0 X B1 1.18e-19
C1 VGND C1 0.0176f
C2 VPWR VPB 0.0754f
C3 A2 A1 0.0881f
C4 VGND A2 0.0191f
C5 a_80_21# A1 0.111f
C6 A1 B1 0.0834f
C7 X a_472_297# 2.6e-19
C8 a_80_21# VGND 0.293f
C9 VGND B1 0.0175f
C10 a_300_47# a_80_21# 0.00997f
C11 X VPB 0.0118f
C12 VGND a_472_297# 0.00188f
C13 a_217_297# C1 0.00262f
C14 VPB A1 0.0266f
C15 VGND VPB 0.00775f
C16 a_217_297# A2 0.0135f
C17 a_80_21# a_217_297# 0.127f
C18 a_217_297# B1 0.00651f
C19 a_80_21# C1 0.079f
C20 C1 B1 0.0846f
C21 X VPWR 0.0884f
C22 a_217_297# a_472_297# 0.00517f
C23 a_80_21# A2 0.128f
C24 a_217_297# VPB 0.00494f
C25 a_80_21# B1 0.0964f
C26 VPWR A1 0.0149f
C27 VPWR VGND 0.0665f
C28 C1 VPB 0.0379f
C29 a_300_47# VPWR 8.53e-19
C30 a_80_21# a_472_297# 0.0164f
C31 a_472_297# B1 1.87e-19
C32 A2 VPB 0.0384f
C33 X A1 3.62e-19
C34 a_80_21# VPB 0.0661f
C35 VPB B1 0.0267f
C36 X VGND 0.0654f
C37 a_300_47# X 5.31e-19
C38 VGND A1 0.0147f
C39 a_217_297# VPWR 0.197f
C40 a_300_47# A1 5.95e-19
C41 a_300_47# VGND 0.00536f
C42 VPWR C1 0.0137f
C43 VPWR A2 0.0161f
C44 X a_217_297# 0.00271f
C45 a_80_21# VPWR 0.119f
C46 VPWR B1 0.0129f
C47 X C1 7.15e-20
C48 a_217_297# A1 0.0124f
C49 a_217_297# VGND 0.00342f
C50 VPWR a_472_297# 0.00703f
C51 X A2 6.82e-19
C52 X a_80_21# 0.118f
C53 VGND VNB 0.385f
C54 VPWR VNB 0.325f
C55 X VNB 0.0899f
C56 C1 VNB 0.144f
C57 B1 VNB 0.0899f
C58 A1 VNB 0.0905f
C59 A2 VNB 0.108f
C60 VPB VNB 0.693f
C61 a_217_297# VNB 0.00117f
C62 a_80_21# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_197_47# a_27_47# 0.00167f
C1 VPB D 0.0782f
C2 VGND B 0.0453f
C3 C B 0.161f
C4 B a_27_47# 0.13f
C5 X VGND 0.0903f
C6 a_197_47# VPWR 5.24e-19
C7 A VGND 0.0151f
C8 X a_27_47# 0.0754f
C9 VPB VGND 0.00852f
C10 A a_27_47# 0.153f
C11 VPWR B 0.0231f
C12 VPB C 0.0609f
C13 VPB a_27_47# 0.082f
C14 X VPWR 0.0945f
C15 A VPWR 0.044f
C16 VPB VPWR 0.077f
C17 D VGND 0.0898f
C18 C D 0.18f
C19 D a_27_47# 0.107f
C20 a_109_47# VGND 0.00223f
C21 C a_109_47# 1.72e-20
C22 a_109_47# a_27_47# 0.00578f
C23 D VPWR 0.0207f
C24 C VGND 0.0408f
C25 VGND a_27_47# 0.132f
C26 a_109_47# VPWR 4.66e-19
C27 C a_27_47# 0.0516f
C28 VPWR VGND 0.0662f
C29 C VPWR 0.021f
C30 VPWR a_27_47# 0.326f
C31 a_197_47# B 0.00623f
C32 D a_303_47# 0.00119f
C33 A B 0.0839f
C34 VPB B 0.0643f
C35 X VPB 0.0111f
C36 a_303_47# VGND 0.00381f
C37 C a_303_47# 0.00527f
C38 A VPB 0.0907f
C39 a_303_47# a_27_47# 0.00119f
C40 a_303_47# VPWR 4.83e-19
C41 a_197_47# VGND 0.00387f
C42 X D 0.00746f
C43 a_109_47# B 0.00153f
C44 a_197_47# C 0.00123f
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X a_489_413# a_226_47#
+ a_556_47# a_226_297# a_76_199#
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPWR B1 0.0188f
C1 A2_N X 2.55e-19
C2 VGND a_226_47# 0.149f
C3 a_556_47# B2 0.00291f
C4 VPB B2 0.0645f
C5 A2_N VPB 0.0327f
C6 a_76_199# B2 0.0626f
C7 B2 B1 0.182f
C8 VGND X 0.0627f
C9 VPWR a_489_413# 0.143f
C10 a_76_199# A2_N 0.0125f
C11 a_226_297# a_76_199# 0.00354f
C12 VGND a_556_47# 0.00639f
C13 VGND VPB 0.0128f
C14 a_489_413# B2 0.0541f
C15 VGND a_76_199# 0.108f
C16 VGND B1 0.0471f
C17 a_226_47# X 0.0108f
C18 VGND a_489_413# 0.0058f
C19 a_226_47# VPB 0.111f
C20 a_76_199# a_226_47# 0.188f
C21 X VPB 0.0113f
C22 a_76_199# X 0.0995f
C23 VPWR A1_N 0.00672f
C24 a_226_47# a_489_413# 0.00579f
C25 a_76_199# a_556_47# 0.0017f
C26 a_76_199# VPB 0.0817f
C27 VPB B1 0.0803f
C28 a_76_199# B1 0.00185f
C29 A1_N A2_N 0.11f
C30 a_489_413# VPB 0.015f
C31 a_226_297# A1_N 0.00184f
C32 a_76_199# a_489_413# 0.0473f
C33 a_489_413# B1 0.0382f
C34 VGND A1_N 0.0261f
C35 VPWR B2 0.0161f
C36 VPWR A2_N 0.00449f
C37 a_226_297# VPWR 8.54e-19
C38 VPWR VGND 0.0743f
C39 a_226_47# A1_N 0.0209f
C40 A1_N X 0.00211f
C41 VGND B2 0.0335f
C42 VGND A2_N 0.0174f
C43 a_226_297# VGND 5.63e-19
C44 A1_N VPB 0.0339f
C45 VPWR a_226_47# 0.0187f
C46 a_76_199# A1_N 0.119f
C47 VPWR X 0.0589f
C48 a_226_47# B2 0.0975f
C49 a_226_47# A2_N 0.141f
C50 VPWR a_556_47# 7.24e-19
C51 VPWR VPB 0.0951f
C52 a_226_297# a_226_47# 0.00128f
C53 VPWR a_76_199# 0.2f
C54 VGND VNB 0.462f
C55 A2_N VNB 0.103f
C56 A1_N VNB 0.111f
C57 VPWR VNB 0.369f
C58 X VNB 0.0975f
C59 B1 VNB 0.206f
C60 B2 VNB 0.106f
C61 VPB VNB 0.782f
C62 a_489_413# VNB 0.0254f
C63 a_226_47# VNB 0.162f
C64 a_76_199# VNB 0.141f
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X a_515_93# a_223_47#
+ a_615_93# a_343_93# a_429_93# a_27_47#
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
C0 a_343_93# a_27_47# 0.0406f
C1 a_515_93# a_223_47# 0.00482f
C2 D a_223_47# 4.03e-19
C3 VPWR VPB 0.106f
C4 VGND VPB 0.0167f
C5 a_515_93# VPWR 7.86e-19
C6 a_515_93# VGND 0.00408f
C7 A_N VPB 0.0848f
C8 VPB a_27_47# 0.154f
C9 D VPWR 0.0143f
C10 D VGND 0.0414f
C11 a_343_93# C 0.0397f
C12 a_615_93# VPWR 8.49e-19
C13 a_615_93# VGND 0.0044f
C14 a_343_93# X 0.126f
C15 C VPB 0.0686f
C16 a_515_93# C 0.00389f
C17 D C 0.163f
C18 B_N a_223_47# 0.0431f
C19 X VPB 0.0103f
C20 D X 0.0193f
C21 a_615_93# C 0.00407f
C22 B_N VPWR 0.0168f
C23 B_N VGND 0.0427f
C24 A_N B_N 0.117f
C25 B_N a_27_47# 0.138f
C26 a_223_47# VPWR 0.114f
C27 a_223_47# VGND 0.199f
C28 A_N a_223_47# 0.00833f
C29 a_223_47# a_27_47# 0.267f
C30 VPWR VGND 0.0906f
C31 a_343_93# a_429_93# 0.00484f
C32 B_N C 9.56e-20
C33 A_N VPWR 0.0318f
C34 A_N VGND 0.0146f
C35 VPWR a_27_47# 0.0897f
C36 VGND a_27_47# 0.0715f
C37 a_223_47# C 0.151f
C38 A_N a_27_47# 0.0906f
C39 B_N X 4.64e-20
C40 C VPWR 0.012f
C41 C VGND 0.025f
C42 VPWR X 0.0582f
C43 VGND X 0.0609f
C44 a_343_93# VPB 0.0857f
C45 a_343_93# a_515_93# 0.00115f
C46 D a_343_93# 0.114f
C47 a_343_93# a_615_93# 0.00103f
C48 D VPB 0.081f
C49 a_429_93# a_223_47# 0.00492f
C50 D a_615_93# 0.00564f
C51 a_429_93# VPWR 5.19e-19
C52 a_429_93# VGND 0.00122f
C53 a_343_93# B_N 0.00112f
C54 a_343_93# a_223_47# 0.269f
C55 B_N VPB 0.0646f
C56 a_343_93# VPWR 0.255f
C57 a_343_93# VGND 0.0548f
C58 D B_N 6.67e-20
C59 a_223_47# VPB 0.0799f
C60 VGND VNB 0.553f
C61 X VNB 0.0908f
C62 VPWR VNB 0.453f
C63 D VNB 0.124f
C64 C VNB 0.107f
C65 B_N VNB 0.134f
C66 A_N VNB 0.144f
C67 VPB VNB 0.959f
C68 a_343_93# VNB 0.172f
C69 a_223_47# VNB 0.141f
C70 a_27_47# VNB 0.259f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VGND VPWR 0.0643f
C1 a_285_47# X 0.00206f
C2 B A 0.221f
C3 a_35_297# A 0.0633f
C4 A VPWR 0.0348f
C5 a_285_47# B 3.98e-19
C6 VGND a_285_297# 0.00394f
C7 a_285_47# a_35_297# 0.00723f
C8 a_285_47# VPWR 8.6e-19
C9 VGND VPB 0.00696f
C10 a_285_297# A 0.00749f
C11 a_117_297# X 2.25e-19
C12 VPB A 0.051f
C13 a_117_297# B 0.00777f
C14 a_35_297# a_117_297# 0.00641f
C15 a_117_297# VPWR 0.00852f
C16 X B 0.0149f
C17 a_35_297# X 0.166f
C18 X VPWR 0.0537f
C19 a_35_297# B 0.203f
C20 B VPWR 0.0703f
C21 X a_285_297# 0.0712f
C22 a_35_297# VPWR 0.096f
C23 X VPB 0.0154f
C24 a_285_297# B 0.0553f
C25 a_35_297# a_285_297# 0.025f
C26 a_285_297# VPWR 0.246f
C27 B VPB 0.0697f
C28 VGND A 0.0325f
C29 a_35_297# VPB 0.0699f
C30 VPB VPWR 0.0689f
C31 a_285_47# VGND 0.00552f
C32 a_285_297# VPB 0.0133f
C33 VGND a_117_297# 0.00177f
C34 VGND X 0.173f
C35 VGND B 0.0304f
C36 X A 0.00166f
C37 VGND a_35_297# 0.177f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X a_465_297# a_297_297#
+ a_215_297# a_392_297# a_109_53#
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 a_297_297# a_215_297# 0.00659f
C1 VPB D_N 0.0461f
C2 a_392_297# VGND 3.44e-19
C3 A a_109_53# 1.19e-19
C4 X VPWR 0.0885f
C5 VPB a_109_53# 0.0547f
C6 B VPWR 0.255f
C7 VPWR a_215_297# 0.0871f
C8 A X 0.00127f
C9 a_297_297# C 0.00375f
C10 a_465_297# a_215_297# 0.00827f
C11 A B 0.0666f
C12 VPB X 0.011f
C13 A a_215_297# 0.157f
C14 a_297_297# VGND 6.5e-19
C15 VPB B 0.116f
C16 VPB a_215_297# 0.0508f
C17 C VPWR 0.00753f
C18 a_465_297# C 6.89e-19
C19 A C 0.0281f
C20 D_N a_109_53# 0.0889f
C21 VGND VPWR 0.075f
C22 VPB C 0.0337f
C23 a_465_297# VGND 5.02e-19
C24 A VGND 0.0158f
C25 VPB VGND 0.0115f
C26 D_N a_215_297# 3.19e-19
C27 B a_109_53# 0.0246f
C28 a_109_53# a_215_297# 0.0807f
C29 B X 6.65e-19
C30 X a_215_297# 0.0991f
C31 a_109_53# C 0.0984f
C32 B a_215_297# 0.159f
C33 D_N VGND 0.0531f
C34 a_392_297# VPWR 5.29e-19
C35 a_109_53# VGND 0.118f
C36 B C 0.0893f
C37 C a_215_297# 0.161f
C38 X VGND 0.0359f
C39 a_297_297# VPWR 8.59e-19
C40 B VGND 0.0161f
C41 VGND a_215_297# 0.237f
C42 C VGND 0.0202f
C43 a_465_297# VPWR 7.08e-19
C44 A VPWR 0.0073f
C45 A a_465_297# 5.42e-19
C46 VPB VPWR 0.122f
C47 VPB A 0.0325f
C48 a_392_297# a_215_297# 0.00419f
C49 a_297_297# a_109_53# 7.06e-21
C50 D_N VPWR 0.0412f
C51 a_392_297# C 0.00267f
C52 a_109_53# VPWR 0.0418f
C53 VGND VNB 0.469f
C54 X VNB 0.0884f
C55 A VNB 0.108f
C56 C VNB 0.101f
C57 D_N VNB 0.185f
C58 B VNB 0.101f
C59 VPWR VNB 0.399f
C60 VPB VNB 0.782f
C61 a_109_53# VNB 0.159f
C62 a_215_297# VNB 0.142f
.ends

.subckt therm b[0] b[2] b[3] p[0] p[10] p[11] p[12] p[13] p[14] p[1] p[2] p[3] p[4]
+ p[5] p[6] p[7] p[8] p[9] input3/a_27_47# _30_/a_297_297# _43_/a_369_47# net7 _35_/a_556_47#
+ input13/a_27_47# _43_/a_469_47# _42_/a_368_53# _25_ _30_/a_215_297# _40_/a_191_297#
+ output19/a_27_47# net19 net4 _24_ input10/a_27_47# _18_ _10_ _52_/a_93_21# _31_/a_35_297#
+ _07_ input7/a_27_47# _04_ output16/a_27_47# input9/a_75_212# _30_/a_109_53# _40_/a_109_297#
+ b[1] _42_/a_209_311# _44_/a_584_47# _27_/a_27_297# input1/a_75_212# _41_/a_59_75#
+ input5/a_62_47# _27_/a_277_297# net2 input14/a_27_47# net3 _42_/a_296_53# input5/a_841_47#
+ _31_/a_285_297# _47_/a_81_21# _35_/a_76_199# input1/A net14 _55_/a_217_297# input5/a_381_47#
+ _27_/a_205_297# _13_ _34_/a_47_47# net15 _37_/a_109_47# _19_ input11/a_27_47# _23_
+ net12 _34_/a_285_47# net18 _49_/a_75_199# _47_/a_384_47# net8 net6 net11 _17_ input8/a_27_47#
+ _33_/a_209_311# _09_ output17/a_27_47# _01_ _37_/a_27_47# _38_/a_109_47# _48_/a_109_47#
+ _47_/a_299_297# _44_/a_250_297# _44_/a_93_21# _48_/a_181_47# _44_/a_346_47# _37_/a_197_47#
+ net13 _42_/a_109_93# _02_ input15/a_27_47# _43_/a_27_47# _43_/a_193_413# _37_/a_303_47#
+ _55_/a_80_21# _50_/a_515_93# input2/a_27_47# _33_/a_109_93# _38_/a_197_47# input5/a_558_47#
+ _15_ _21_ _50_/a_615_93# _14_ input12/a_27_47# _20_ net1 _38_/a_303_47# _38_/a_27_47#
+ _40_/a_297_297# _34_/a_129_47# _03_ _06_ _53_/a_29_53# _49_/a_315_47# net16 net10
+ output18/a_27_47# _08_ input5/a_664_47# _16_ _11_ _27_/a_109_297# _12_ net9 _00_
+ _44_/a_256_47# _05_ _48_/a_27_47# input6/a_27_47# net17 _31_/a_117_297# _50_/a_343_93#
+ net5 VPWR VGND _29_/a_29_53#
X_49_ net7 _02_ _19_ _20_ _21_ VGND VGND VPWR VPWR net17 _49_/a_208_47# _49_/a_75_199#
+ _49_/a_544_297# _49_/a_315_47# _49_/a_201_297# sky130_fd_sc_hd__a311o_1
X_48_ net11 _02_ _07_ VGND VGND VPWR VPWR _21_ _48_/a_181_47# _48_/a_109_47# _48_/a_27_47#
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ net5 _12_ _17_ VGND VGND VPWR VPWR _20_ _47_/a_384_47# _47_/a_81_21# _47_/a_299_297#
+ sky130_fd_sc_hd__a21o_1
X_46_ _04_ VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__inv_2
X_29_ net11 net13 net12 VGND VGND VPWR VPWR _03_ _29_/a_29_53# _29_/a_183_297# _29_/a_111_297#
+ sky130_fd_sc_hd__or3_1
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28_ _00_ _01_ VGND VGND VPWR VPWR _02_ _28_/a_109_297# sky130_fd_sc_hd__nor2_1
X_45_ _02_ _09_ _12_ _13_ _18_ VGND VGND VPWR VPWR net16 _45_/a_193_297# _45_/a_465_47#
+ _45_/a_205_47# _45_/a_109_297# _45_/a_27_47# sky130_fd_sc_hd__a221o_1
X_44_ net14 _14_ _15_ _17_ net2 VGND VGND VPWR VPWR _18_ _44_/a_256_47# _44_/a_584_47#
+ _44_/a_93_21# _44_/a_250_297# _44_/a_346_47# sky130_fd_sc_hd__a32o_1
X_27_ net14 net15 net3 net2 VGND VGND VPWR VPWR _01_ _27_/a_277_297# _27_/a_205_297#
+ _27_/a_27_297# _27_/a_109_297# sky130_fd_sc_hd__or4_1
XFILLER_0_7_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_26_ net5 net4 net6 VGND VGND VPWR VPWR _00_ _26_/a_29_53# _26_/a_183_297# _26_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_43_ _00_ _06_ _10_ _16_ VGND VGND VPWR VPWR _17_ _43_/a_369_47# _43_/a_469_47# _43_/a_297_47#
+ _43_/a_193_413# _43_/a_27_47# sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_42_ net3 net15 net14 VGND VGND VPWR VPWR _16_ _42_/a_109_93# _42_/a_368_53# _42_/a_209_311#
+ _42_/a_296_53# sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_3_Left_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND VPWR VPWR b[0] output16/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_41_ _06_ _10_ VGND VGND VPWR VPWR _15_ _41_/a_145_75# _41_/a_59_75# sky130_fd_sc_hd__and2_1
Xoutput17 net17 VGND VGND VPWR VPWR b[1] output17/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_40_ net15 net3 net2 _00_ VGND VGND VPWR VPWR _14_ _40_/a_297_297# _40_/a_191_297#
+ _40_/a_109_297# sky130_fd_sc_hd__nor4_1
Xoutput18 net18 VGND VGND VPWR VPWR b[2] output18/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR b[3] output19/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_7_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 input1/A VGND VGND VPWR VPWR net1 input1/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput2 p[10] VGND VGND VPWR VPWR net2 input2/a_27_47# sky130_fd_sc_hd__buf_1
Xinput3 p[11] VGND VGND VPWR VPWR net3 input3/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 p[12] VGND VGND VPWR VPWR net4 input4/a_75_212# sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 p[13] VGND VGND VPWR VPWR net5 input5/a_664_47# input5/a_841_47# input5/a_381_47#
+ input5/a_62_47# input5/a_558_47# sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_1_Left_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 p[14] VGND VGND VPWR VPWR net6 input6/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 p[1] VGND VGND VPWR VPWR net7 input7/a_27_47# sky130_fd_sc_hd__buf_1
Xinput10 p[4] VGND VGND VPWR VPWR net10 input10/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 p[2] VGND VGND VPWR VPWR net8 input8/a_27_47# sky130_fd_sc_hd__buf_1
Xinput11 p[5] VGND VGND VPWR VPWR net11 input11/a_27_47# sky130_fd_sc_hd__buf_1
X_39_ net5 net6 VGND VGND VPWR VPWR _13_ _39_/a_129_47# _39_/a_47_47# _39_/a_285_47#
+ _39_/a_377_297# sky130_fd_sc_hd__xnor2_1
Xinput9 p[3] VGND VGND VPWR VPWR net9 input9/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput12 p[6] VGND VGND VPWR VPWR net12 input12/a_27_47# sky130_fd_sc_hd__buf_1
X_55_ _14_ _15_ _20_ _22_ VGND VGND VPWR VPWR net19 _55_/a_472_297# _55_/a_80_21#
+ _55_/a_300_47# _55_/a_217_297# sky130_fd_sc_hd__a211o_1
X_38_ net4 _06_ _10_ _11_ VGND VGND VPWR VPWR _12_ _38_/a_109_47# _38_/a_197_47# _38_/a_303_47#
+ _38_/a_27_47# sky130_fd_sc_hd__and4_1
X_54_ _25_ VGND VGND VPWR VPWR net18 _54_/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput13 p[7] VGND VGND VPWR VPWR net13 input13/a_27_47# sky130_fd_sc_hd__buf_1
X_37_ net14 net15 net3 net2 VGND VGND VPWR VPWR _11_ _37_/a_109_47# _37_/a_197_47#
+ _37_/a_303_47# _37_/a_27_47# sky130_fd_sc_hd__and4_1
X_53_ _21_ _22_ _24_ VGND VGND VPWR VPWR _25_ _53_/a_29_53# _53_/a_183_297# _53_/a_111_297#
+ sky130_fd_sc_hd__or3_1
Xinput14 p[8] VGND VGND VPWR VPWR net14 input14/a_27_47# sky130_fd_sc_hd__buf_1
X_36_ net11 net10 net13 net12 VGND VGND VPWR VPWR _10_ _36_/a_109_47# _36_/a_197_47#
+ _36_/a_303_47# _36_/a_27_47# sky130_fd_sc_hd__and4_1
X_52_ _02_ _06_ _23_ _12_ net5 VGND VGND VPWR VPWR _24_ _52_/a_256_47# _52_/a_584_47#
+ _52_/a_93_21# _52_/a_250_297# _52_/a_346_47# sky130_fd_sc_hd__a32o_1
X_35_ _04_ _05_ _07_ _08_ VGND VGND VPWR VPWR _09_ _35_/a_489_413# _35_/a_226_47#
+ _35_/a_556_47# _35_/a_226_297# _35_/a_76_199# sky130_fd_sc_hd__a2bb2o_1
Xinput15 p[9] VGND VGND VPWR VPWR net15 input15/a_27_47# sky130_fd_sc_hd__buf_1
X_51_ _03_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__inv_2
X_34_ net11 net12 VGND VGND VPWR VPWR _08_ _34_/a_129_47# _34_/a_47_47# _34_/a_285_47#
+ _34_/a_377_297# sky130_fd_sc_hd__xnor2_1
X_33_ net13 _06_ net10 VGND VGND VPWR VPWR _07_ _33_/a_109_93# _33_/a_368_53# _33_/a_209_311#
+ _33_/a_296_53# sky130_fd_sc_hd__and3b_1
X_50_ net5 net6 _15_ _11_ VGND VGND VPWR VPWR _22_ _50_/a_515_93# _50_/a_223_47# _50_/a_615_93#
+ _50_/a_343_93# _50_/a_429_93# _50_/a_27_47# sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ net7 net1 net9 net8 VGND VGND VPWR VPWR _06_ _32_/a_109_47# _32_/a_197_47# _32_/a_303_47#
+ _32_/a_27_47# sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_5_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31_ net7 net8 VGND VGND VPWR VPWR _05_ _31_/a_117_297# _31_/a_285_297# _31_/a_285_47#
+ _31_/a_35_297# sky130_fd_sc_hd__xor2_1
X_30_ net9 net10 _03_ net1 VGND VGND VPWR VPWR _04_ _30_/a_465_297# _30_/a_297_297#
+ _30_/a_215_297# _30_/a_392_297# _30_/a_109_53# sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
C0 p[6] net10 0.00236f
C1 _20_ _16_ 0.00271f
C2 p[2] VPWR 0.113f
C3 _02_ _00_ 0.0269f
C4 _47_/a_81_21# _11_ 0.0454f
C5 b[1] _31_/a_285_47# 8.76e-19
C6 _31_/a_285_297# net8 0.0215f
C7 net17 _49_/a_75_199# 0.00127f
C8 b[1] _27_/a_27_297# 0.00644f
C9 _06_ _45_/a_193_297# 0.00201f
C10 VPWR b[3] 0.144f
C11 input11/a_27_47# p[4] 0.0646f
C12 _36_/a_27_47# net13 0.0488f
C13 input4/a_75_212# _10_ 0.00372f
C14 b[1] net18 0.00134f
C15 net6 _43_/a_27_47# 9.07e-20
C16 _52_/a_584_47# _02_ 0.00389f
C17 _17_ _50_/a_223_47# 5.24e-20
C18 b[3] _41_/a_59_75# 9.66e-22
C19 p[2] _31_/a_285_297# 0.00175f
C20 p[12] net15 2.99e-19
C21 p[11] p[13] 0.0137f
C22 _04_ net7 0.0602f
C23 _07_ _24_ 5.67e-19
C24 _35_/a_76_199# _05_ 0.00238f
C25 input2/a_27_47# net8 0.0207f
C26 net5 _32_/a_197_47# 5.61e-21
C27 net15 p[9] 0.00295f
C28 p[7] _35_/a_76_199# 1.78e-19
C29 net11 _45_/a_27_47# 3.64e-20
C30 p[13] input5/a_381_47# 0.00146f
C31 _36_/a_27_47# _21_ 0.0276f
C32 _23_ _11_ 2e-20
C33 net7 net14 2.23e-19
C34 _02_ _27_/a_27_297# 0.00179f
C35 _34_/a_47_47# b[1] 0.0197f
C36 _33_/a_368_53# _05_ 9.2e-19
C37 p[3] _10_ 1.37e-20
C38 _04_ _49_/a_544_297# 0.00204f
C39 _53_/a_29_53# _25_ 0.00146f
C40 _08_ _35_/a_489_413# 5.56e-19
C41 _04_ _49_/a_75_199# 0.0782f
C42 _43_/a_193_413# p[9] 1.09e-19
C43 _02_ net18 8.53e-20
C44 output19/a_27_47# net14 0.00142f
C45 _04_ _44_/a_93_21# 4.47e-21
C46 _42_/a_296_53# net14 2.18e-19
C47 _42_/a_209_311# _01_ 1.58e-19
C48 _14_ _43_/a_369_47# 0.00135f
C49 b[1] _10_ 2.37e-20
C50 net19 net5 0.00124f
C51 net6 net2 0.00139f
C52 net5 _30_/a_109_53# 5.84e-22
C53 input5/a_664_47# b[1] 0.00195f
C54 net12 _35_/a_489_413# 3.97e-20
C55 p[4] net10 0.00268f
C56 _42_/a_209_311# _22_ 1.72e-19
C57 net13 _35_/a_226_297# 6.88e-19
C58 net6 _37_/a_27_47# 4.3e-20
C59 net14 _49_/a_75_199# 3.67e-19
C60 p[13] net2 0.0246f
C61 _03_ _26_/a_29_53# 7.93e-21
C62 _39_/a_47_47# _11_ 3.9e-19
C63 _32_/a_27_47# net5 0.0961f
C64 net13 _33_/a_109_93# 0.0254f
C65 VPWR _40_/a_109_297# -4.23e-19
C66 net14 _44_/a_93_21# 0.0646f
C67 _14_ _26_/a_183_297# 6.98e-22
C68 _22_ _26_/a_29_53# 0.09f
C69 _03_ _24_ 9.46e-20
C70 _31_/a_35_297# _19_ 1.47e-19
C71 net13 _09_ 0.0379f
C72 _34_/a_47_47# _02_ 1.09e-19
C73 _20_ _42_/a_209_311# 1.66e-20
C74 b[1] _30_/a_465_297# 4.8e-19
C75 _00_ _30_/a_109_53# 3.67e-20
C76 _40_/a_191_297# _06_ 5.84e-19
C77 _22_ _24_ 0.0846f
C78 net3 _37_/a_109_47# 0.00212f
C79 net15 _37_/a_303_47# 0.00118f
C80 _32_/a_27_47# _00_ 0.00228f
C81 _21_ _33_/a_109_93# 1.62e-20
C82 _50_/a_343_93# net8 7.25e-19
C83 _20_ _26_/a_29_53# 0.00447f
C84 _02_ _10_ 0.0537f
C85 input8/a_27_47# p[3] 0.0023f
C86 input5/a_664_47# _02_ 0.00187f
C87 _18_ _36_/a_27_47# 5.46e-20
C88 net13 _06_ 0.0758f
C89 _14_ _47_/a_81_21# 6.24e-20
C90 input8/a_27_47# b[1] 0.00172f
C91 _36_/a_27_47# VPWR -0.00832f
C92 _21_ _09_ 0.263f
C93 b[1] _35_/a_226_47# 0.00334f
C94 p[11] net15 3.03e-20
C95 _54_/a_75_212# net18 0.0143f
C96 p[5] net18 1.98e-19
C97 net5 _01_ 0.0779f
C98 p[13] net9 1.72e-19
C99 _36_/a_109_47# _06_ 0.00168f
C100 net5 _03_ 1.04e-19
C101 net7 _49_/a_208_47# 0.00312f
C102 _34_/a_47_47# input12/a_27_47# 2.17e-19
C103 net1 _49_/a_201_297# 0.00304f
C104 net19 _27_/a_27_297# 1.98e-19
C105 _17_ _02_ 0.00482f
C106 net5 _22_ 0.405f
C107 input6/a_27_47# p[12] 2.78e-19
C108 input5/a_381_47# net15 7.15e-19
C109 _21_ _06_ 0.143f
C110 _28_/a_109_297# _10_ 4.34e-19
C111 net4 _39_/a_377_297# 8.88e-19
C112 _29_/a_29_53# net3 1.68e-20
C113 _23_ net10 0.00216f
C114 net16 _24_ 6.93e-19
C115 _19_ net8 0.0322f
C116 _03_ _00_ 2.31e-20
C117 input6/a_27_47# p[9] 0.0756f
C118 input8/a_27_47# _02_ 5.08e-20
C119 _01_ _00_ 0.00124f
C120 net3 net17 3.72e-19
C121 _35_/a_556_47# _09_ 0.00122f
C122 _20_ net5 0.0651f
C123 net1 input1/a_75_212# 0.00208f
C124 net7 b[1] 0.0783f
C125 _15_ _44_/a_250_297# 0.00517f
C126 _50_/a_615_93# _10_ 8.82e-19
C127 _12_ _52_/a_93_21# 0.0157f
C128 _02_ _35_/a_226_47# 2.21e-19
C129 _22_ _00_ 0.477f
C130 _33_/a_209_311# _09_ 3.79e-20
C131 _04_ _52_/a_93_21# 2.35e-19
C132 input7/a_27_47# net17 4.99e-20
C133 _17_ _37_/a_197_47# 9.19e-21
C134 p[2] _19_ 1.08e-19
C135 input11/a_27_47# net11 0.00318f
C136 p[10] net3 3.61e-19
C137 VPWR _35_/a_226_297# -8.54e-19
C138 net2 net15 0.324f
C139 _42_/a_296_53# b[1] 2.38e-20
C140 _04_ _49_/a_315_47# 7.71e-19
C141 VPWR _33_/a_109_93# -0.00817f
C142 p[11] _16_ 4e-20
C143 p[3] input13/a_27_47# 0.00101f
C144 _49_/a_75_199# p[3] 1.79e-20
C145 _39_/a_47_47# net10 4.72e-22
C146 _42_/a_209_311# p[9] 5.51e-21
C147 _16_ _43_/a_27_47# 2.47e-19
C148 net15 _37_/a_27_47# 0.0541f
C149 output18/a_27_47# _25_ 0.072f
C150 _34_/a_285_47# _08_ 0.00414f
C151 _04_ _27_/a_109_297# 7.2e-20
C152 _52_/a_584_47# _22_ 6.24e-19
C153 net10 _52_/a_250_297# 2.86e-21
C154 _34_/a_47_47# _07_ 0.011f
C155 net12 net8 0.00458f
C156 _20_ _00_ 0.271f
C157 _18_ _09_ 7.01e-21
C158 _39_/a_47_47# b[0] 2.04e-19
C159 b[1] input13/a_27_47# 0.00624f
C160 _04_ _34_/a_377_297# 1.7e-20
C161 b[1] _49_/a_75_199# 0.00805f
C162 net1 _31_/a_35_297# 0.0111f
C163 VPWR _09_ 0.297f
C164 b[1] _49_/a_544_297# 8.23e-19
C165 _33_/a_209_311# _06_ 0.0187f
C166 net2 _43_/a_193_413# 1.52e-19
C167 net16 net5 0.00476f
C168 net19 _10_ 0.00224f
C169 _03_ _31_/a_285_47# 8.54e-19
C170 net19 input5/a_664_47# 1.38e-21
C171 _01_ _31_/a_285_47# 3.36e-19
C172 _55_/a_80_21# net14 4.7e-19
C173 _07_ _10_ 2.19e-19
C174 net12 _34_/a_285_47# 8.07e-20
C175 _03_ _27_/a_27_297# 2.68e-19
C176 net7 _02_ 0.445f
C177 net3 _12_ 3.09e-20
C178 _43_/a_193_413# _37_/a_27_47# 0.0102f
C179 _32_/a_27_47# _10_ 0.00217f
C180 _35_/a_489_413# _45_/a_27_47# 3.89e-21
C181 input5/a_62_47# _44_/a_250_297# 2.45e-20
C182 _04_ net3 0.113f
C183 net14 _27_/a_109_297# 1.32e-19
C184 _01_ _27_/a_27_297# 8.04e-19
C185 _15_ net8 1.79e-19
C186 _55_/a_217_297# _14_ 0.0116f
C187 _55_/a_472_297# _15_ 0.00626f
C188 p[14] net14 6.11e-20
C189 net10 _34_/a_129_47# 0.003f
C190 input5/a_558_47# net2 5.99e-21
C191 _18_ _06_ 0.54f
C192 net18 _03_ 2.07e-21
C193 VPWR _06_ 1.4f
C194 net2 _16_ 0.00654f
C195 _22_ net18 1.68e-19
C196 net15 net9 8.49e-20
C197 VPWR _31_/a_117_297# 5.04e-19
C198 _41_/a_59_75# _06_ 0.0429f
C199 _02_ _49_/a_75_199# 0.0354f
C200 net10 net11 0.592f
C201 net14 net3 0.689f
C202 _16_ _37_/a_27_47# 2.07e-19
C203 _17_ net19 0.0269f
C204 _20_ _27_/a_27_297# 3.14e-20
C205 input9/a_75_212# net10 0.00699f
C206 p[1] net15 1.81e-19
C207 input7/a_27_47# net14 3.48e-19
C208 _36_/a_303_47# net11 7.63e-20
C209 net5 p[12] 4.99e-20
C210 net14 input14/a_27_47# 0.0232f
C211 _53_/a_29_53# _24_ 0.0835f
C212 b[3] _15_ 1.89e-19
C213 _31_/a_285_297# _06_ 1.01e-20
C214 _34_/a_47_47# _03_ 4.5e-20
C215 _48_/a_109_47# _06_ 9.47e-19
C216 input10/a_27_47# _25_ 2.03e-20
C217 VPWR _44_/a_256_47# -7.56e-19
C218 input5/a_62_47# net8 2.05e-19
C219 net1 net8 0.381f
C220 _34_/a_47_47# _22_ 3.9e-21
C221 _35_/a_226_47# _07_ 8.96e-19
C222 net6 _35_/a_76_199# 4.6e-21
C223 _01_ _10_ 2.22e-19
C224 _03_ _10_ 0.00244f
C225 input5/a_558_47# net9 4.42e-19
C226 net11 _50_/a_27_47# 6.05e-21
C227 _13_ _09_ 0.0927f
C228 p[11] _42_/a_209_311# 2.58e-19
C229 VPWR _47_/a_299_297# 0.0643f
C230 _38_/a_197_47# _12_ 0.00173f
C231 _22_ _10_ 0.0904f
C232 input5/a_558_47# p[1] 1.61e-21
C233 p[2] net1 0.0274f
C234 VPWR _39_/a_129_47# -9.47e-19
C235 net16 net18 0.00585f
C236 VPWR _52_/a_346_47# -0.00109f
C237 _41_/a_59_75# _47_/a_299_297# 0.00146f
C238 b[2] _09_ 4.28e-20
C239 _42_/a_209_311# input5/a_381_47# 3.88e-19
C240 _38_/a_109_47# _10_ 5.44e-19
C241 _39_/a_285_47# _06_ 1.23e-20
C242 net9 _30_/a_392_297# 9.92e-19
C243 _03_ _30_/a_465_297# 7.72e-19
C244 _55_/a_300_47# VPWR -4.61e-19
C245 _20_ _10_ 0.179f
C246 _13_ _06_ 0.00188f
C247 input6/a_27_47# net2 0.0047f
C248 _17_ _01_ 1.46e-20
C249 net19 output19/a_27_47# 0.0273f
C250 input6/a_27_47# _37_/a_27_47# 9.35e-19
C251 b[1] _52_/a_93_21# 2.82e-19
C252 p[5] input13/a_27_47# 3.09e-19
C253 net19 _42_/a_296_53# 2.71e-19
C254 _32_/a_27_47# net7 0.00559f
C255 _36_/a_27_47# net4 0.0103f
C256 _17_ _22_ 0.00334f
C257 net6 net15 0.0664f
C258 VPWR _45_/a_193_297# -0.00859f
C259 _55_/a_80_21# b[1] 6.03e-19
C260 _00_ _05_ 5.03e-22
C261 p[6] _48_/a_27_47# 4.48e-19
C262 b[2] _06_ 0.0116f
C263 input1/A output17/a_27_47# 0.00805f
C264 b[1] _49_/a_315_47# 5.66e-19
C265 input8/a_27_47# _01_ 1.43e-19
C266 _42_/a_209_311# net2 5.1e-19
C267 p[13] net15 1.46e-19
C268 b[1] _27_/a_109_297# 8.35e-20
C269 _03_ _35_/a_226_47# 0.028f
C270 net16 _10_ 0.0338f
C271 _49_/a_75_199# _07_ 4.05e-21
C272 _42_/a_209_311# _37_/a_27_47# 1.59e-20
C273 b[1] _34_/a_377_297# 0.00115f
C274 _36_/a_109_47# net13 0.00126f
C275 _36_/a_27_47# net12 0.0185f
C276 _17_ _20_ 0.102f
C277 net19 _44_/a_93_21# 0.0074f
C278 _22_ _35_/a_226_47# 1.39e-20
C279 VPWR p[8] 0.148f
C280 net6 _43_/a_193_413# 2.41e-20
C281 _21_ net13 0.13f
C282 _50_/a_343_93# _06_ 0.0376f
C283 net3 b[1] 0.00334f
C284 net5 _32_/a_303_47# 7.18e-21
C285 _02_ _52_/a_93_21# 0.0962f
C286 _20_ _35_/a_226_47# 5.19e-20
C287 b[3] input15/a_27_47# 0.00109f
C288 input7/a_27_47# b[1] 0.00663f
C289 VPWR output17/a_27_47# 0.0268f
C290 _02_ _49_/a_315_47# 0.00134f
C291 net11 _45_/a_109_297# 7.46e-20
C292 _55_/a_80_21# _02_ 0.164f
C293 _31_/a_285_47# _05_ 5.61e-19
C294 p[13] input5/a_558_47# 0.00156f
C295 net5 input5/a_381_47# 0.0546f
C296 net7 _03_ 0.078f
C297 net6 _16_ 1.62e-20
C298 net7 _01_ 0.233f
C299 net14 _43_/a_369_47# 6.79e-21
C300 input3/a_27_47# _44_/a_250_297# 2.07e-19
C301 net7 _22_ 2.73e-20
C302 _19_ _09_ 4.8e-21
C303 _00_ _43_/a_27_47# 0.0431f
C304 _53_/a_29_53# net18 0.0118f
C305 b[3] _44_/a_584_47# 1.26e-19
C306 p[12] _10_ 0.0994f
C307 _42_/a_368_53# net14 7.39e-19
C308 _14_ _43_/a_469_47# 0.00259f
C309 net4 _09_ 0.00262f
C310 input5/a_841_47# b[1] 7.07e-19
C311 _10_ p[9] 0.00225f
C312 net9 _26_/a_29_53# 0.00343f
C313 _49_/a_75_199# _03_ 0.0849f
C314 net3 _02_ 9.52e-20
C315 _08_ _09_ 0.106f
C316 net12 _33_/a_109_93# 0.0435f
C317 _01_ _49_/a_75_199# 0.009f
C318 net13 _33_/a_209_311# 0.0227f
C319 _03_ _49_/a_544_297# 0.00568f
C320 _39_/a_377_297# _11_ 2.57e-20
C321 net5 net2 0.0616f
C322 _36_/a_27_47# net1 6.99e-20
C323 _01_ _49_/a_544_297# 0.00109f
C324 _20_ net7 0.0257f
C325 net10 _35_/a_489_413# 0.00225f
C326 _22_ _49_/a_75_199# 9.85e-21
C327 net5 _37_/a_27_47# 1.13e-20
C328 VPWR _40_/a_191_297# -6.82e-19
C329 _22_ _26_/a_111_297# 0.00137f
C330 _47_/a_81_21# _12_ 0.00158f
C331 _53_/a_29_53# _34_/a_47_47# 5.88e-22
C332 _55_/a_80_21# _28_/a_109_297# 2.05e-20
C333 net12 _09_ 0.0374f
C334 net4 _06_ 0.281f
C335 _34_/a_47_47# _05_ 1.26e-20
C336 net8 _11_ 1.81e-20
C337 _14_ _49_/a_201_297# 4.76e-21
C338 _40_/a_297_297# _06_ 1.64e-19
C339 _18_ net13 1.06e-20
C340 input2/a_27_47# output17/a_27_47# 0.107f
C341 _08_ _06_ 0.0343f
C342 _21_ _35_/a_556_47# 2.69e-19
C343 VPWR net13 0.599f
C344 net3 _37_/a_197_47# 0.0028f
C345 net2 _00_ 0.00732f
C346 _53_/a_29_53# _10_ 0.00779f
C347 _20_ _49_/a_75_199# 0.0233f
C348 _17_ p[9] 1.03e-20
C349 _10_ _05_ 9.25e-21
C350 input5/a_841_47# _02_ 0.00591f
C351 _00_ _37_/a_27_47# 6.15e-20
C352 p[6] b[1] 0.0043f
C353 net6 input6/a_27_47# 0.00208f
C354 _36_/a_109_47# VPWR -4.66e-19
C355 net12 _06_ 0.284f
C356 input5/a_381_47# _27_/a_27_297# 1.47e-19
C357 _31_/a_285_297# net13 3.85e-20
C358 net19 _55_/a_80_21# 0.00423f
C359 net5 net9 0.0368f
C360 net15 _43_/a_193_413# 0.00169f
C361 VPWR _21_ 0.869f
C362 _23_ _12_ 0.00743f
C363 input3/a_27_47# b[3] 1.4e-19
C364 _36_/a_197_47# _06_ 6.18e-19
C365 _31_/a_35_297# net10 3.95e-20
C366 net19 p[14] 0.101f
C367 _15_ _06_ 0.22f
C368 net6 _42_/a_209_311# 1.32e-20
C369 input5/a_558_47# net15 0.00672f
C370 net4 _47_/a_299_297# 3.28e-19
C371 net2 _27_/a_27_297# 0.0131f
C372 _34_/a_377_297# _07_ 5.8e-19
C373 _29_/a_29_53# net11 0.00514f
C374 net6 _26_/a_29_53# 0.0032f
C375 net1 _09_ 5.26e-20
C376 net9 _00_ 0.00501f
C377 _39_/a_47_47# _12_ 0.0317f
C378 input9/a_75_212# _29_/a_29_53# 9.7e-21
C379 _16_ net15 0.214f
C380 input8/a_27_47# _05_ 1.58e-19
C381 net17 net11 3.19e-20
C382 _43_/a_27_47# _10_ 0.0279f
C383 net19 net3 0.611f
C384 output19/a_27_47# p[12] 1.78e-19
C385 input1/A VPWR 0.0833f
C386 _14_ _44_/a_250_297# 4.82e-19
C387 _12_ _52_/a_250_297# 0.0139f
C388 net6 _24_ 0.00121f
C389 _04_ _52_/a_250_297# 3.98e-21
C390 _35_/a_226_47# _05_ 0.0134f
C391 net11 _30_/a_215_297# 1.04e-19
C392 VPWR _35_/a_556_47# -7.24e-19
C393 net19 input14/a_27_47# 3.63e-19
C394 _17_ _37_/a_303_47# 1.23e-20
C395 _13_ net13 4e-21
C396 output19/a_27_47# p[9] 0.0832f
C397 _42_/a_368_53# b[1] 5.32e-20
C398 input9/a_75_212# _30_/a_215_297# 6.24e-21
C399 VPWR _33_/a_209_311# -0.0131f
C400 net1 _06_ 0.0115f
C401 _35_/a_226_47# p[7] 3.42e-19
C402 _42_/a_109_93# _44_/a_250_297# 6.38e-19
C403 _16_ _43_/a_193_413# 0.0261f
C404 output18/a_27_47# net18 0.0106f
C405 _29_/a_183_297# _10_ 6.24e-20
C406 net4 _45_/a_193_297# 7.41e-19
C407 _04_ _27_/a_205_297# 6.42e-19
C408 p[4] b[1] 0.00675f
C409 net10 _52_/a_256_47# 8.13e-20
C410 _03_ _52_/a_93_21# 0.00985f
C411 _15_ _47_/a_299_297# 0.0103f
C412 _40_/a_109_297# _11_ 0.00522f
C413 _18_ VPWR 0.0721f
C414 net10 net8 2.05e-21
C415 p[6] input12/a_27_47# 0.0176f
C416 _03_ _49_/a_315_47# 9.22e-19
C417 _55_/a_217_297# net14 2.1e-19
C418 _55_/a_80_21# _01_ 0.0121f
C419 _17_ _43_/a_27_47# 0.00131f
C420 _22_ _52_/a_93_21# 0.0347f
C421 _30_/a_297_297# _10_ 1.25e-20
C422 _01_ _49_/a_315_47# 1.82e-19
C423 net14 _27_/a_205_297# 3.63e-19
C424 _03_ _27_/a_109_297# 1.97e-20
C425 net7 _05_ 0.0129f
C426 net2 _10_ 3.15e-19
C427 net11 _12_ 0.00799f
C428 _13_ _21_ 1.69e-19
C429 _14_ net8 4.23e-19
C430 _04_ net11 0.078f
C431 _55_/a_80_21# _22_ 0.00926f
C432 _55_/a_300_47# _15_ 1.42e-20
C433 _55_/a_472_297# _14_ 0.00192f
C434 net6 net5 0.725f
C435 p[1] _27_/a_27_297# 4.83e-19
C436 _03_ _34_/a_377_297# 3.13e-20
C437 net10 _34_/a_285_47# 0.0454f
C438 input5/a_664_47# net2 8.11e-20
C439 VPWR _41_/a_59_75# 0.0292f
C440 _04_ input9/a_75_212# 7.69e-22
C441 output17/a_27_47# _19_ 7.69e-19
C442 p[13] net5 0.00689f
C443 _09_ _45_/a_27_47# 0.00823f
C444 input6/a_27_47# net15 0.00115f
C445 p[6] p[5] 0.0388f
C446 _21_ b[2] 2.14e-19
C447 _01_ net3 1.16e-19
C448 VPWR _31_/a_285_297# 0.013f
C449 net3 _03_ 4.27e-20
C450 _55_/a_80_21# _20_ 0.0291f
C451 net14 net11 9.95e-19
C452 input13/a_27_47# _05_ 3.93e-19
C453 _48_/a_27_47# net11 0.0179f
C454 net6 _00_ 0.00178f
C455 net3 _22_ 9.39e-20
C456 _17_ net2 0.181f
C457 _34_/a_47_47# net9 1.41e-20
C458 input13/a_27_47# p[7] 0.0205f
C459 input10/a_27_47# net18 4.16e-20
C460 _06_ input15/a_27_47# 4.73e-19
C461 input4/a_75_212# _39_/a_47_47# 3.1e-19
C462 _48_/a_181_47# _06_ 6.4e-19
C463 p[6] _07_ 2.01e-19
C464 VPWR _44_/a_346_47# -8.74e-19
C465 _17_ _37_/a_27_47# 0.00277f
C466 _06_ _45_/a_27_47# 0.0021f
C467 _42_/a_209_311# net15 0.0157f
C468 input2/a_27_47# VPWR 0.00832f
C469 net9 _10_ 0.0438f
C470 _38_/a_27_47# net11 1.68e-20
C471 _20_ net3 4.07e-19
C472 net7 _43_/a_27_47# 6.31e-19
C473 _02_ _47_/a_81_21# 1.59e-20
C474 input5/a_664_47# net9 5.29e-19
C475 net15 _26_/a_29_53# 9.06e-21
C476 _23_ b[1] 7.65e-19
C477 p[4] input12/a_27_47# 8.26e-19
C478 VPWR _47_/a_384_47# -1.45e-19
C479 _18_ _13_ 0.019f
C480 _38_/a_303_47# _12_ 0.00153f
C481 VPWR _39_/a_285_47# -9.53e-19
C482 input5/a_664_47# p[1] 1.21e-20
C483 input5/a_381_47# net7 4.91e-19
C484 net13 _19_ 4.45e-20
C485 _13_ VPWR 0.0804f
C486 net5 _35_/a_76_199# 3.38e-19
C487 net4 net13 2.48e-19
C488 _42_/a_209_311# input5/a_558_47# 7.85e-20
C489 net9 _30_/a_465_297# 0.00138f
C490 net13 _08_ 1.82e-19
C491 input5/a_62_47# p[8] 1.22e-19
C492 _17_ net9 2.89e-23
C493 p[4] p[5] 0.235f
C494 _09_ _45_/a_465_47# 2.77e-19
C495 VPWR b[2] 0.262f
C496 _42_/a_209_311# _16_ 0.00129f
C497 net5 _25_ 6.42e-19
C498 net2 net7 0.00234f
C499 net19 _42_/a_368_53# 5.12e-19
C500 VPWR _45_/a_205_47# -1.62e-19
C501 _23_ _02_ 0.0648f
C502 _09_ _11_ 0.0665f
C503 net13 net12 0.363f
C504 _14_ _40_/a_109_297# -1.78e-33
C505 output19/a_27_47# net2 0.00168f
C506 p[14] p[12] 0.00101f
C507 input8/a_27_47# net9 3.71e-20
C508 input5/a_62_47# output17/a_27_47# 1.02e-19
C509 net4 _21_ 0.00535f
C510 net1 output17/a_27_47# 8.12e-19
C511 net9 _35_/a_226_47# 1.22e-20
C512 b[1] _27_/a_205_297# 1.41e-19
C513 input8/a_27_47# p[1] 5.13e-20
C514 _21_ _08_ 0.00139f
C515 net5 net15 0.0226f
C516 _18_ _50_/a_343_93# 0.0276f
C517 _36_/a_197_47# net13 1.06e-19
C518 VPWR _50_/a_343_93# -0.0126f
C519 p[14] p[9] 0.355f
C520 b[1] _34_/a_129_47# 3.51e-19
C521 net6 _43_/a_297_47# 8.23e-22
C522 _11_ _06_ 0.493f
C523 _36_/a_27_47# net10 0.0366f
C524 _21_ net12 0.23f
C525 net2 _44_/a_93_21# 0.0273f
C526 _41_/a_59_75# _50_/a_343_93# 6.13e-22
C527 _39_/a_47_47# _02_ 0.0127f
C528 net6 _10_ 0.0965f
C529 _50_/a_429_93# _06_ 0.00169f
C530 net5 _43_/a_193_413# 1.39e-20
C531 _53_/a_29_53# _52_/a_93_21# 0.00116f
C532 input9/a_75_212# p[3] 0.0158f
C533 net15 _00_ 0.00147f
C534 _02_ _52_/a_250_297# 0.0128f
C535 _13_ _39_/a_285_47# 0.00451f
C536 b[1] net11 0.0777f
C537 _52_/a_93_21# _05_ 1.12e-20
C538 _37_/a_27_47# _44_/a_93_21# 3.19e-19
C539 net3 p[9] 1.63e-19
C540 input9/a_75_212# b[1] 0.00598f
C541 _55_/a_217_297# _02_ 6.01e-19
C542 p[13] input5/a_664_47# 7.57e-19
C543 net7 net9 0.00233f
C544 net5 input5/a_558_47# 0.0597f
C545 input14/a_27_47# p[9] 8.53e-21
C546 _21_ _15_ 1.13e-21
C547 _38_/a_197_47# net16 5.89e-19
C548 _32_/a_27_47# _47_/a_81_21# 5.06e-21
C549 _08_ _35_/a_556_47# 7.71e-19
C550 net14 _43_/a_469_47# 1.44e-20
C551 p[1] net7 0.00514f
C552 _00_ _43_/a_193_413# 0.00721f
C553 _08_ _33_/a_209_311# 0.0122f
C554 _36_/a_27_47# _50_/a_27_47# 6.08e-19
C555 net5 _16_ 1.99e-20
C556 _53_/a_111_297# _09_ 3.4e-19
C557 _04_ _49_/a_201_297# 0.0253f
C558 net1 net13 3.51e-19
C559 _17_ net6 3.12e-19
C560 VPWR _19_ 0.0335f
C561 _31_/a_35_297# net17 0.0514f
C562 _13_ _45_/a_205_47# 7.51e-20
C563 _18_ net4 0.023f
C564 net9 input13/a_27_47# 2.42e-19
C565 _49_/a_75_199# net9 0.00382f
C566 _47_/a_299_297# _11_ 0.00738f
C567 net12 _33_/a_209_311# 0.0769f
C568 _02_ net11 0.0327f
C569 _25_ net18 0.0594f
C570 net4 VPWR 1.08f
C571 _31_/a_35_297# _30_/a_215_297# 6.37e-19
C572 net10 _35_/a_226_297# 2.48e-19
C573 p[10] _31_/a_35_297# 2.39e-19
C574 net15 _27_/a_27_297# 0.00888f
C575 VPWR _08_ -0.0171f
C576 VPWR _40_/a_297_297# -5.42e-19
C577 _16_ _00_ 0.00613f
C578 _22_ _26_/a_183_297# 0.00184f
C579 _53_/a_111_297# _06_ 3.82e-19
C580 net14 _49_/a_201_297# 1.52e-19
C581 net10 _33_/a_109_93# 0.0336f
C582 net4 _41_/a_59_75# 1.76e-19
C583 _31_/a_285_297# _19_ 1.34e-19
C584 _23_ _07_ 1.27e-19
C585 _13_ _50_/a_343_93# 5.63e-20
C586 net1 _21_ 0.0252f
C587 _18_ net12 2.25e-21
C588 _35_/a_76_199# _10_ 7.19e-20
C589 _55_/a_80_21# p[11] 6.43e-20
C590 _55_/a_80_21# _43_/a_27_47# 1.56e-19
C591 _32_/a_109_47# net8 0.0011f
C592 net10 _09_ 0.037f
C593 VPWR net12 0.82f
C594 net3 _37_/a_303_47# 0.00133f
C595 _01_ _47_/a_81_21# 6.05e-21
C596 _34_/a_47_47# _25_ 1.08e-19
C597 _11_ _45_/a_193_297# 0.0292f
C598 _18_ _15_ 0.042f
C599 _04_ _31_/a_35_297# 1.89e-20
C600 _36_/a_197_47# VPWR -5.24e-19
C601 _22_ _47_/a_81_21# 7.25e-19
C602 input12/a_27_47# net11 0.00246f
C603 input5/a_558_47# _27_/a_27_297# 1.57e-19
C604 input2/a_27_47# _19_ 5.26e-20
C605 VPWR _15_ 0.929f
C606 net10 _06_ 0.184f
C607 _26_/a_29_53# _24_ 2.11e-20
C608 _25_ _10_ 0.0109f
C609 input5/a_62_47# input1/A 1.39e-19
C610 input1/A net1 0.00473f
C611 p[11] net3 0.00296f
C612 net17 net8 0.18f
C613 _36_/a_303_47# _06_ 5.3e-19
C614 _41_/a_59_75# _15_ 0.0139f
C615 _04_ _44_/a_250_297# 5.57e-21
C616 _16_ _27_/a_27_297# 3.74e-22
C617 p[8] _11_ 5.85e-20
C618 _14_ _06_ 0.0556f
C619 _09_ _50_/a_27_47# 1.3e-19
C620 net6 output19/a_27_47# 0.00112f
C621 p[11] input14/a_27_47# 3.98e-20
C622 input3/a_27_47# p[8] 6.2e-19
C623 _20_ _47_/a_81_21# 0.0457f
C624 net8 _30_/a_215_297# 8.14e-21
C625 p[13] net7 1.91e-19
C626 net15 _10_ 0.0101f
C627 p[10] net8 0.00463f
C628 _54_/a_75_212# net11 0.00956f
C629 input5/a_381_47# net3 0.0299f
C630 input5/a_664_47# net15 0.0216f
C631 p[5] net11 0.0599f
C632 net4 _39_/a_285_47# 9.71e-19
C633 net2 _27_/a_109_297# 7.24e-20
C634 _29_/a_183_297# net3 7.38e-21
C635 _29_/a_111_297# net11 8.27e-19
C636 _42_/a_109_93# _06_ 5.53e-20
C637 _23_ _03_ 0.0564f
C638 _13_ net4 0.212f
C639 p[14] net2 1.38e-19
C640 _42_/a_209_311# net5 3.27e-21
C641 _35_/a_226_47# _35_/a_76_199# -2.84e-32
C642 net6 _26_/a_111_297# 1.12e-19
C643 net14 _44_/a_250_297# 4.24e-20
C644 _39_/a_377_297# _12_ 6.77e-19
C645 p[14] _37_/a_27_47# 1.37e-19
C646 input3/a_27_47# output17/a_27_47# 3.15e-19
C647 _43_/a_193_413# _10_ 0.0174f
C648 _23_ _22_ 0.0187f
C649 _21_ _45_/a_27_47# 1.18e-20
C650 _06_ _50_/a_27_47# 0.00972f
C651 input5/a_62_47# VPWR 0.0601f
C652 _14_ _44_/a_256_47# 0.00124f
C653 net1 VPWR 1.17f
C654 net6 _44_/a_93_21# 1.08e-20
C655 p[6] p[7] 0.0545f
C656 net5 _26_/a_29_53# 0.0237f
C657 net11 _07_ 0.0206f
C658 net2 net3 0.519f
C659 _04_ net8 0.02f
C660 input2/a_27_47# _15_ 3.18e-20
C661 _17_ net15 0.195f
C662 net3 _37_/a_27_47# 0.094f
C663 _39_/a_47_47# _03_ 1.47e-19
C664 net5 _24_ 5.83e-20
C665 input7/a_27_47# net2 3.24e-19
C666 _04_ _27_/a_277_297# 0.00113f
C667 net2 input14/a_27_47# 0.0235f
C668 _15_ _47_/a_384_47# 0.00112f
C669 net1 _31_/a_285_297# 5.85e-19
C670 net7 _35_/a_76_199# 1.79e-20
C671 _16_ _10_ 0.00486f
C672 _00_ _26_/a_29_53# 0.0466f
C673 _39_/a_129_47# b[0] 2.6e-20
C674 _13_ _15_ 3.69e-20
C675 b[1] _35_/a_489_413# 0.00104f
C676 _40_/a_191_297# _11_ 0.00207f
C677 _17_ _43_/a_193_413# 0.0503f
C678 _22_ _52_/a_250_297# 0.0996f
C679 _04_ p[2] 3.32e-20
C680 b[1] _49_/a_201_297# 0.0025f
C681 net14 net8 0.0516f
C682 _55_/a_217_297# _01_ 0.00112f
C683 net4 _50_/a_343_93# 0.00124f
C684 _03_ _27_/a_205_297# 1.46e-20
C685 net14 _27_/a_277_297# 5.1e-19
C686 _55_/a_300_47# _14_ 8.09e-19
C687 _52_/a_584_47# _26_/a_29_53# 7.45e-20
C688 _20_ _39_/a_47_47# 2.3e-20
C689 p[1] _27_/a_109_297# 8.88e-21
C690 _17_ input5/a_558_47# 2.13e-21
C691 VPWR _41_/a_145_75# 3.84e-19
C692 _48_/a_27_47# _34_/a_285_47# 6.66e-20
C693 net1 input2/a_27_47# 4.81e-19
C694 input5/a_841_47# _37_/a_27_47# 4.64e-20
C695 _18_ input15/a_27_47# 8.27e-21
C696 net3 net9 5.09e-20
C697 input1/a_75_212# b[1] 0.0074f
C698 _42_/a_209_311# _27_/a_27_297# 4.7e-20
C699 _17_ _16_ 0.242f
C700 _18_ _45_/a_27_47# 0.00347f
C701 _03_ net11 0.0952f
C702 _55_/a_217_297# _20_ 0.0013f
C703 VPWR input15/a_27_47# 0.0198f
C704 _01_ net11 3.82e-20
C705 VPWR _48_/a_181_47# -3.35e-19
C706 VPWR _45_/a_27_47# -0.00418f
C707 b[3] net14 9.2e-19
C708 p[1] net3 0.00192f
C709 input9/a_75_212# _03_ 9.32e-20
C710 net7 net15 2.91e-19
C711 _02_ _35_/a_489_413# 3.86e-19
C712 p[4] p[7] 7.8e-20
C713 _22_ net11 6.82e-21
C714 _41_/a_59_75# input15/a_27_47# 3.96e-20
C715 _15_ _50_/a_343_93# 0.0098f
C716 net16 _39_/a_47_47# 7.7e-20
C717 output19/a_27_47# net15 6.88e-19
C718 input7/a_27_47# p[1] 0.0164f
C719 VPWR _44_/a_584_47# -2.28e-19
C720 net5 _00_ 0.00954f
C721 _06_ _45_/a_109_297# 0.0023f
C722 _21_ _11_ 9.98e-20
C723 net18 _26_/a_29_53# 2.57e-21
C724 _31_/a_35_297# b[1] 0.0176f
C725 _36_/a_27_47# _29_/a_29_53# 6.92e-20
C726 input6/a_27_47# _10_ 4.57e-20
C727 _20_ net11 0.00128f
C728 net7 _43_/a_193_413# 3.49e-19
C729 output17/a_27_47# net10 1.31e-20
C730 net15 _49_/a_75_199# 5.13e-20
C731 net18 _24_ 5.57e-21
C732 input5/a_841_47# net9 2.7e-19
C733 _52_/a_584_47# net5 0.0022f
C734 net6 _52_/a_93_21# 2.33e-19
C735 input5/a_558_47# net7 0.00358f
C736 net15 _44_/a_93_21# 0.00573f
C737 _36_/a_27_47# _30_/a_215_297# 7.13e-20
C738 net6 p[14] 0.00245f
C739 net8 _49_/a_208_47# 1.4e-19
C740 _42_/a_109_93# output17/a_27_47# 8.6e-21
C741 _42_/a_209_311# input5/a_664_47# 0.0124f
C742 net4 net12 2.57e-20
C743 p[12] _39_/a_47_47# 3.32e-19
C744 net7 _16_ 7.5e-20
C745 _31_/a_35_297# _02_ 0.00316f
C746 net12 _08_ 0.0269f
C747 net16 net11 4.43e-22
C748 _15_ _19_ 1.46e-20
C749 _17_ input6/a_27_47# 7.13e-22
C750 _43_/a_193_413# _44_/a_93_21# 0.0161f
C751 net5 _27_/a_27_297# 3.48e-19
C752 _34_/a_47_47# _24_ 6.84e-21
C753 _26_/a_29_53# _10_ 0.0265f
C754 p[12] _52_/a_250_297# 1.84e-20
C755 p[2] _49_/a_208_47# 3.83e-20
C756 p[3] net8 0.0015f
C757 b[1] _52_/a_256_47# 8.49e-20
C758 net6 net3 0.00152f
C759 _13_ _45_/a_27_47# 0.0703f
C760 net4 _15_ 0.00427f
C761 _53_/a_111_297# _21_ 4.38e-19
C762 input5/a_558_47# _44_/a_93_21# 2.71e-19
C763 _14_ _40_/a_191_297# 2.4e-19
C764 VPWR _45_/a_465_47# -5.05e-19
C765 _24_ _10_ 0.00484f
C766 _36_/a_27_47# _12_ 0.00178f
C767 _18_ _11_ 0.484f
C768 b[1] net8 0.0729f
C769 _04_ _36_/a_27_47# 0.00169f
C770 VPWR _11_ 0.352f
C771 p[13] net3 3.64e-19
C772 b[1] _27_/a_277_297# 1.24e-19
C773 net13 net10 0.375f
C774 input3/a_27_47# VPWR 0.0688f
C775 _17_ _42_/a_209_311# 1.22e-19
C776 _16_ _44_/a_93_21# 0.00354f
C777 p[2] p[3] 0.0394f
C778 _36_/a_197_47# net12 4.67e-20
C779 _36_/a_303_47# net13 5.5e-20
C780 VPWR _50_/a_429_93# -3.61e-19
C781 b[1] _34_/a_285_47# 0.00368f
C782 p[13] input14/a_27_47# 3.88e-19
C783 _41_/a_59_75# _11_ 8.7e-19
C784 _35_/a_489_413# _07_ 0.00429f
C785 _35_/a_76_199# _52_/a_93_21# 6.83e-21
C786 _29_/a_29_53# _09_ 0.00488f
C787 p[2] b[1] 0.0022f
C788 p[6] input10/a_27_47# 0.00214f
C789 input5/a_62_47# _19_ 0.00159f
C790 net1 _19_ 2.86e-19
C791 _33_/a_109_93# _30_/a_215_297# 0.00104f
C792 _50_/a_515_93# _06_ 0.00244f
C793 _52_/a_250_297# _05_ 8.86e-22
C794 _02_ _52_/a_256_47# 0.00344f
C795 _21_ net10 0.0275f
C796 net13 _50_/a_27_47# 7.27e-21
C797 _55_/a_472_297# _02_ 1.25e-19
C798 net5 _10_ 0.199f
C799 p[13] input5/a_841_47# 1.59e-19
C800 _02_ net8 0.334f
C801 net5 input5/a_664_47# 0.0536f
C802 _29_/a_29_53# _06_ 0.00111f
C803 _38_/a_303_47# net16 6.47e-19
C804 net2 _47_/a_81_21# 4.95e-19
C805 output19/a_27_47# input6/a_27_47# 0.107f
C806 input11/a_27_47# VPWR 0.0375f
C807 _00_ _43_/a_297_47# 1.26e-19
C808 _36_/a_27_47# _50_/a_223_47# 1.27e-20
C809 _35_/a_226_297# _12_ 3.35e-20
C810 _02_ _34_/a_285_47# 7.14e-19
C811 _53_/a_183_297# _09_ 4.18e-19
C812 net1 net12 1.17e-19
C813 _33_/a_109_93# _12_ 9.75e-20
C814 _04_ _35_/a_226_297# 4.51e-19
C815 p[2] _02_ 8.19e-19
C816 _04_ _33_/a_109_93# 0.0299f
C817 _00_ _10_ 0.301f
C818 _06_ _30_/a_215_297# 2.03e-20
C819 _31_/a_117_297# net17 0.00149f
C820 _53_/a_29_53# net11 8.31e-19
C821 _21_ _50_/a_27_47# 3.38e-21
C822 VPWR _53_/a_111_297# 1.11e-34
C823 _13_ _45_/a_465_47# 0.00134f
C824 _55_/a_80_21# net15 0.00759f
C825 _47_/a_384_47# _11_ 7.23e-20
C826 _31_/a_35_297# _30_/a_109_53# 2.89e-20
C827 net11 _05_ 2.76e-19
C828 _04_ _09_ 0.0904f
C829 _17_ net5 0.00408f
C830 _09_ _12_ 0.00526f
C831 input6/a_27_47# _44_/a_93_21# 8.53e-19
C832 _32_/a_27_47# _31_/a_35_297# 9.17e-20
C833 _03_ _35_/a_489_413# 0.0205f
C834 net10 _35_/a_556_47# 5.59e-19
C835 _13_ _11_ 0.164f
C836 p[14] net15 0.00137f
C837 input9/a_75_212# _05_ 1.24e-21
C838 net10 _33_/a_209_311# 0.0426f
C839 _03_ _49_/a_201_297# 0.00842f
C840 _53_/a_183_297# _06_ 0.00146f
C841 _01_ _49_/a_201_297# 0.0105f
C842 net19 _44_/a_250_297# 0.00592f
C843 input9/a_75_212# p[7] 0.00102f
C844 _22_ _49_/a_201_297# 2.45e-20
C845 _55_/a_80_21# _43_/a_193_413# 2.54e-19
C846 _55_/a_217_297# _43_/a_27_47# 2.18e-19
C847 _32_/a_197_47# net8 3.39e-20
C848 _17_ _00_ 0.0851f
C849 _06_ _12_ 0.136f
C850 input10/a_27_47# p[4] 0.0215f
C851 _04_ _06_ 0.0132f
C852 _48_/a_27_47# _09_ 0.00541f
C853 _42_/a_209_311# _44_/a_93_21# 2.21e-19
C854 _47_/a_81_21# net9 3.49e-19
C855 _18_ net10 1.47e-21
C856 net15 net3 0.394f
C857 net4 _45_/a_27_47# 0.024f
C858 VPWR net10 0.375f
C859 input7/a_27_47# net15 1.88e-19
C860 _20_ _49_/a_201_297# 5.24e-21
C861 _18_ _14_ 0.243f
C862 _36_/a_303_47# VPWR -4.83e-19
C863 VPWR b[0] 0.142f
C864 input5/a_664_47# _27_/a_27_297# 0.0116f
C865 VPWR _14_ 0.186f
C866 input5/a_62_47# net1 7.59e-20
C867 net14 _06_ 1.94e-19
C868 _55_/a_80_21# _16_ 0.0143f
C869 net3 _43_/a_193_413# 5.65e-20
C870 _38_/a_27_47# _09_ 0.00195f
C871 net19 net8 1.15e-19
C872 _48_/a_27_47# _06_ 0.0251f
C873 net6 _43_/a_369_47# 3.62e-21
C874 _50_/a_343_93# _11_ 0.0384f
C875 _31_/a_35_297# _03_ 0.00749f
C876 _31_/a_285_297# net10 1.68e-19
C877 VPWR _42_/a_109_93# -0.00118f
C878 _31_/a_35_297# _01_ 4.27e-19
C879 _18_ _50_/a_27_47# 0.0665f
C880 net8 _30_/a_109_53# 1.76e-20
C881 _36_/a_27_47# b[1] 7.95e-19
C882 net5 net7 0.195f
C883 input5/a_558_47# net3 0.0137f
C884 input5/a_841_47# net15 0.00585f
C885 _32_/a_27_47# net8 0.0275f
C886 VPWR _50_/a_27_47# -0.00335f
C887 _15_ input15/a_27_47# 2.15e-20
C888 input7/a_27_47# input5/a_558_47# 1.22e-20
C889 _17_ _27_/a_27_297# 6.78e-22
C890 _29_/a_183_297# net11 3.64e-19
C891 _23_ net9 1.21e-19
C892 _34_/a_285_47# _07_ 0.00975f
C893 _38_/a_27_47# _06_ 0.0172f
C894 _47_/a_299_297# _12_ 0.00805f
C895 _41_/a_59_75# _50_/a_27_47# 9.59e-22
C896 net14 _44_/a_256_47# 0.00379f
C897 _16_ net3 1.77e-19
C898 _39_/a_129_47# _12_ 0.00175f
C899 _06_ _50_/a_223_47# 0.0481f
C900 _43_/a_297_47# _10_ 0.00118f
C901 net7 _00_ 8.12e-21
C902 _14_ _44_/a_346_47# 3.76e-19
C903 _12_ _52_/a_346_47# 3.8e-19
C904 net19 b[3] 0.054f
C905 input2/a_27_47# net10 1.17e-20
C906 _20_ _31_/a_35_297# 1.69e-19
C907 net5 _44_/a_93_21# 3.61e-20
C908 _36_/a_27_47# _02_ 9.37e-20
C909 net6 _47_/a_81_21# 2.14e-19
C910 _13_ net10 4.52e-21
C911 _09_ _49_/a_208_47# 5.43e-21
C912 _39_/a_285_47# b[0] 1.88e-19
C913 _00_ _26_/a_111_297# 3.7e-19
C914 _13_ b[0] 0.00299f
C915 net4 _11_ 0.0858f
C916 input4/a_75_212# _06_ 0.00205f
C917 _13_ _14_ 1.47e-20
C918 input5/a_841_47# _16_ 8.62e-19
C919 _45_/a_193_297# _12_ 0.0103f
C920 output17/a_27_47# net17 0.0149f
C921 b[1] _35_/a_226_297# 1.03e-19
C922 output18/a_27_47# net11 6.84e-20
C923 _03_ net8 0.0287f
C924 _17_ _43_/a_297_47# 5.72e-20
C925 _40_/a_297_297# _11_ 9.94e-19
C926 p[14] input6/a_27_47# 0.0157f
C927 b[1] _33_/a_109_93# 0.00411f
C928 _55_/a_472_297# _01_ 6.28e-19
C929 _01_ net8 0.0802f
C930 _00_ _44_/a_93_21# 4.54e-20
C931 net4 _50_/a_429_93# 4.16e-19
C932 _03_ _27_/a_277_297# 2.1e-20
C933 p[10] output17/a_27_47# 0.117f
C934 net7 _31_/a_285_47# 0.00132f
C935 _22_ net8 3.3e-20
C936 _17_ _10_ 0.0233f
C937 p[1] _27_/a_205_297# 3.18e-20
C938 net7 _27_/a_27_297# 1.22e-19
C939 net12 _11_ 3.82e-21
C940 _47_/a_299_297# _50_/a_223_47# 2.74e-20
C941 b[2] b[0] 0.183f
C942 b[1] _09_ 0.00408f
C943 _13_ _50_/a_27_47# 0.00169f
C944 p[2] _01_ 0.00164f
C945 _33_/a_296_53# _06_ 1.11e-20
C946 _55_/a_80_21# _42_/a_209_311# 0.0175f
C947 input6/a_27_47# net3 2.52e-19
C948 _20_ net8 5.07e-19
C949 _55_/a_472_297# _20_ 0.00212f
C950 p[14] _42_/a_209_311# 3.45e-22
C951 p[3] _06_ 1.59e-20
C952 net9 net11 0.136f
C953 _35_/a_226_47# _10_ 1.25e-19
C954 net6 _23_ 2.13e-19
C955 _15_ _11_ 0.113f
C956 VPWR _45_/a_109_297# -0.011f
C957 input9/a_75_212# net9 0.0245f
C958 input3/a_27_47# _15_ 7.53e-19
C959 _24_ _52_/a_93_21# 0.0211f
C960 b[1] _06_ 0.0885f
C961 _04_ output17/a_27_47# 0.027f
C962 _49_/a_75_199# _27_/a_27_297# 0.011f
C963 _29_/a_29_53# net13 0.00104f
C964 _02_ _33_/a_109_93# 1.54e-21
C965 net14 p[8] 0.00965f
C966 _15_ _50_/a_429_93# 6.82e-19
C967 _14_ _50_/a_343_93# 9.76e-19
C968 _42_/a_209_311# net3 0.029f
C969 _31_/a_117_297# b[1] 0.00281f
C970 net13 net17 5.21e-20
C971 net4 _53_/a_111_297# 2.09e-19
C972 _02_ _09_ 0.297f
C973 net13 _30_/a_215_297# 0.0246f
C974 net6 _39_/a_47_47# 0.0249f
C975 input10/a_27_47# net11 0.112f
C976 net3 _26_/a_29_53# 2.83e-21
C977 _43_/a_369_47# _43_/a_193_413# -1.25e-19
C978 net6 _52_/a_250_297# 0.00133f
C979 net7 _10_ 6.22e-20
C980 _29_/a_29_53# _21_ 0.0775f
C981 input5/a_664_47# net7 0.00199f
C982 output19/a_27_47# _10_ 3.23e-20
C983 input5/a_62_47# input3/a_27_47# 0.00179f
C984 _32_/a_27_47# _36_/a_27_47# 0.011f
C985 net5 _52_/a_93_21# 0.0124f
C986 _02_ _06_ 0.85f
C987 _21_ _30_/a_215_297# 1.48e-19
C988 _55_/a_80_21# net5 2.78e-19
C989 _31_/a_35_297# _05_ 0.00649f
C990 net4 net10 8.28e-22
C991 _14_ _19_ 2.71e-21
C992 net13 _12_ 0.00632f
C993 _26_/a_111_297# _10_ 7.13e-20
C994 VPWR _37_/a_109_47# -4.38e-19
C995 net15 _47_/a_81_21# 0.00106f
C996 _04_ net13 0.569f
C997 net10 _08_ 0.194f
C998 input1/a_75_212# p[0] 0.00122f
C999 b[1] _52_/a_346_47# 6.37e-20
C1000 net4 _14_ 1.54e-20
C1001 _44_/a_93_21# _10_ 2.48e-19
C1002 net4 b[0] 0.0024f
C1003 _42_/a_109_93# _19_ 1.14e-21
C1004 input5/a_664_47# _44_/a_93_21# 1.88e-20
C1005 _14_ _40_/a_297_297# 1.58e-19
C1006 net6 net11 1.08e-19
C1007 _55_/a_300_47# b[1] 1.1e-19
C1008 _04_ _36_/a_109_47# 2.39e-19
C1009 _55_/a_80_21# _00_ 5.5e-19
C1010 _17_ output19/a_27_47# 0.00122f
C1011 net13 net14 2.21e-21
C1012 net12 net10 0.539f
C1013 net5 net3 0.0365f
C1014 input8/a_27_47# net7 1.47e-19
C1015 VPWR _32_/a_109_47# 0.00124f
C1016 p[10] input1/A 6.79e-20
C1017 input12/a_27_47# _06_ 5.3e-22
C1018 net7 _35_/a_226_47# 2.93e-20
C1019 _36_/a_303_47# net12 1.37e-19
C1020 _04_ _21_ 0.39f
C1021 _23_ _25_ 0.00465f
C1022 VPWR _50_/a_515_93# -5.03e-19
C1023 _21_ _12_ 7.99e-20
C1024 net17 _33_/a_209_311# 7.03e-21
C1025 _29_/a_111_297# _09_ 5.79e-20
C1026 _35_/a_76_199# _52_/a_250_297# 3.4e-21
C1027 _20_ _40_/a_109_297# 2.35e-20
C1028 net4 _50_/a_27_47# 0.0239f
C1029 _33_/a_109_93# _07_ 3.2e-19
C1030 p[12] b[3] 7.54e-20
C1031 _33_/a_209_311# _30_/a_215_297# 1.56e-19
C1032 _17_ _44_/a_93_21# 0.0646f
C1033 _50_/a_615_93# _06_ 0.00264f
C1034 VPWR _29_/a_29_53# 0.0299f
C1035 _02_ _52_/a_346_47# 0.00526f
C1036 net3 _00_ 2.12e-19
C1037 _11_ input15/a_27_47# 4.4e-19
C1038 _36_/a_27_47# _22_ 2.82e-20
C1039 _54_/a_75_212# _06_ 0.00727f
C1040 _15_ _14_ 0.148f
C1041 _11_ _45_/a_27_47# 0.0703f
C1042 input8/a_27_47# _49_/a_75_199# 1.99e-20
C1043 _21_ net14 7.17e-21
C1044 _09_ _07_ 0.0416f
C1045 b[3] p[9] 0.107f
C1046 _55_/a_300_47# _02_ 0.00371f
C1047 VPWR net17 0.037f
C1048 _49_/a_75_199# _35_/a_226_47# 8.73e-20
C1049 net12 _50_/a_27_47# 7.99e-21
C1050 _21_ _48_/a_27_47# 0.0121f
C1051 net8 _05_ 0.0146f
C1052 _29_/a_111_297# _06_ 6.74e-20
C1053 _35_/a_226_47# input13/a_27_47# 3.94e-20
C1054 net5 input5/a_841_47# 0.0221f
C1055 VPWR _30_/a_215_297# -0.00548f
C1056 net18 _52_/a_93_21# 8.21e-21
C1057 _42_/a_109_93# _15_ 0.00367f
C1058 p[10] VPWR 0.234f
C1059 _36_/a_27_47# _20_ 0.00148f
C1060 net19 _06_ 0.00522f
C1061 _34_/a_285_47# _05_ 7.85e-21
C1062 _27_/a_27_297# _27_/a_109_297# -3.68e-20
C1063 _39_/a_47_47# net15 9.44e-22
C1064 _33_/a_209_311# _12_ 2.88e-20
C1065 net11 _35_/a_76_199# 4e-19
C1066 _15_ _50_/a_27_47# 5.65e-19
C1067 _02_ _45_/a_193_297# 0.00988f
C1068 p[2] _05_ 4.53e-19
C1069 _06_ _30_/a_109_53# 1.96e-19
C1070 _04_ _33_/a_209_311# 0.00133f
C1071 _06_ _07_ 0.185f
C1072 _38_/a_27_47# _21_ 3.87e-19
C1073 output17/a_27_47# b[1] 0.0373f
C1074 _32_/a_27_47# _06_ 0.00663f
C1075 net1 net10 0.00388f
C1076 _21_ _50_/a_223_47# 2.91e-21
C1077 p[2] p[7] 0.00131f
C1078 _55_/a_217_297# net15 7.79e-19
C1079 _03_ _35_/a_226_297# 0.00101f
C1080 net2 _31_/a_35_297# 0.0635f
C1081 net7 _49_/a_75_199# 0.09f
C1082 net3 _27_/a_27_297# 0.0166f
C1083 _18_ _12_ 0.0115f
C1084 _18_ _04_ 1.94e-21
C1085 net7 _49_/a_544_297# 2.72e-19
C1086 _03_ _33_/a_109_93# 2.78e-19
C1087 VPWR _12_ 0.28f
C1088 input7/a_27_47# _27_/a_27_297# 0.00119f
C1089 _04_ VPWR 0.456f
C1090 _25_ net11 0.0262f
C1091 _22_ _33_/a_109_93# 1.34e-22
C1092 input2/a_27_47# net17 0.0398f
C1093 _32_/a_303_47# net8 2.22e-34
C1094 net2 _44_/a_250_297# 0.0188f
C1095 _41_/a_59_75# _12_ 0.00101f
C1096 _03_ _09_ 0.326f
C1097 _10_ _52_/a_93_21# 0.00534f
C1098 output19/a_27_47# _44_/a_93_21# 7.25e-20
C1099 _01_ _09_ 4.69e-21
C1100 net13 _33_/a_296_53# 3.71e-20
C1101 _18_ net14 0.0147f
C1102 input2/a_27_47# _30_/a_215_297# 3.51e-20
C1103 _55_/a_80_21# _10_ 5.49e-19
C1104 net4 _45_/a_109_297# 6.43e-20
C1105 _22_ _09_ 0.0279f
C1106 p[10] input2/a_27_47# 0.00905f
C1107 input5/a_381_47# net8 7.48e-19
C1108 VPWR net14 0.182f
C1109 net13 p[3] 9.49e-19
C1110 VPWR _48_/a_27_47# 0.0158f
C1111 p[14] _10_ 1.53e-19
C1112 input1/a_75_212# p[1] 0.0023f
C1113 _01_ _06_ 0.00157f
C1114 net13 b[1] 0.0495f
C1115 _03_ _06_ 0.00635f
C1116 _55_/a_217_297# _16_ 0.0017f
C1117 _20_ _09_ 7.11e-19
C1118 net6 _43_/a_469_47# 4.85e-21
C1119 _31_/a_117_297# _03_ 5.32e-19
C1120 _22_ _06_ 0.124f
C1121 net8 _30_/a_297_297# 2.42e-21
C1122 net3 _10_ 3.89e-19
C1123 _18_ _50_/a_223_47# 0.0367f
C1124 _38_/a_27_47# VPWR -0.0142f
C1125 input5/a_664_47# net3 0.00215f
C1126 net2 net8 0.0525f
C1127 _04_ input2/a_27_47# 4.5e-21
C1128 _21_ p[3] 3.79e-20
C1129 _17_ _55_/a_80_21# 7.64e-21
C1130 VPWR _50_/a_223_47# -0.00601f
C1131 _14_ input15/a_27_47# 9.48e-21
C1132 input7/a_27_47# input5/a_664_47# 1.08e-21
C1133 net8 _37_/a_27_47# 6.66e-21
C1134 _17_ p[14] 5.46e-21
C1135 _21_ b[1] 0.00892f
C1136 net14 _44_/a_346_47# 0.00464f
C1137 _20_ _06_ 0.133f
C1138 _47_/a_384_47# _12_ 9.51e-20
C1139 _39_/a_285_47# _12_ 0.0221f
C1140 _35_/a_226_47# _52_/a_93_21# 4.89e-20
C1141 _13_ _12_ 0.462f
C1142 _04_ _13_ 1.17e-21
C1143 net16 _09_ 0.00707f
C1144 net13 _02_ 0.00154f
C1145 VPWR output16/a_27_47# 0.122f
C1146 input2/a_27_47# net14 0.0102f
C1147 net19 p[8] 1.25e-19
C1148 input4/a_75_212# _18_ 4.36e-19
C1149 _17_ net3 0.0698f
C1150 _50_/a_27_47# _45_/a_27_47# 0.109f
C1151 net2 b[3] 0.00395f
C1152 input4/a_75_212# VPWR 0.0739f
C1153 _36_/a_27_47# _05_ 3.67e-21
C1154 b[2] _12_ 3.89e-20
C1155 net16 _06_ 0.0511f
C1156 input1/A b[1] 0.00126f
C1157 input4/a_75_212# _41_/a_59_75# 0.00153f
C1158 _00_ _26_/a_183_297# 4.53e-19
C1159 _45_/a_205_47# _12_ 7.46e-19
C1160 b[1] _35_/a_556_47# 3.23e-19
C1161 _21_ _02_ 0.397f
C1162 input8/a_27_47# input7/a_27_47# 3.2e-20
C1163 _55_/a_300_47# _01_ 0.00113f
C1164 VPWR _49_/a_208_47# -5.93e-19
C1165 net9 net8 0.0605f
C1166 net5 _47_/a_81_21# 4.59e-19
C1167 b[1] _33_/a_209_311# 0.0129f
C1168 p[13] input1/a_75_212# 4.16e-19
C1169 _23_ _24_ 0.012f
C1170 p[6] _34_/a_47_47# 0.00102f
C1171 _55_/a_80_21# net7 0.00163f
C1172 _38_/a_197_47# _10_ 6.29e-19
C1173 VPWR _33_/a_296_53# -1.15e-19
C1174 net7 _49_/a_315_47# 0.00706f
C1175 _55_/a_300_47# _22_ 2.08e-19
C1176 _20_ _47_/a_299_297# 0.002f
C1177 p[1] _27_/a_277_297# 1.57e-20
C1178 _20_ _39_/a_129_47# 1.71e-20
C1179 _50_/a_343_93# _12_ 5.63e-20
C1180 _38_/a_27_47# _13_ 4.58e-19
C1181 _03_ _45_/a_193_297# 2.57e-20
C1182 VPWR p[3] 0.0975f
C1183 p[2] net9 1.4e-20
C1184 net17 _19_ 0.0211f
C1185 _13_ _50_/a_223_47# 8.2e-20
C1186 _47_/a_81_21# _00_ 0.0258f
C1187 p[14] output19/a_27_47# 0.0943f
C1188 VPWR b[1] 1.05f
C1189 _22_ _45_/a_193_297# 0.0234f
C1190 p[2] p[1] 0.0414f
C1191 p[10] _19_ 9.65e-20
C1192 p[12] _06_ 0.0535f
C1193 p[5] net13 1.05e-19
C1194 net14 _50_/a_343_93# 1.07e-20
C1195 _14_ _11_ 0.0415f
C1196 net7 net3 7.45e-20
C1197 _21_ input12/a_27_47# 2.32e-19
C1198 _24_ _52_/a_250_297# 3.03e-19
C1199 _13_ output16/a_27_47# 4.58e-19
C1200 _29_/a_29_53# net12 0.0132f
C1201 net15 _43_/a_469_47# 7.41e-19
C1202 input7/a_27_47# net7 0.00318f
C1203 _33_/a_109_93# _05_ 0.0206f
C1204 net5 _23_ 0.0052f
C1205 net2 _40_/a_109_297# 0.0011f
C1206 _15_ _50_/a_515_93# 0.00147f
C1207 output19/a_27_47# net3 0.00348f
C1208 _06_ p[9] 0.00205f
C1209 _35_/a_226_297# p[7] 1.48e-20
C1210 p[13] _44_/a_250_297# 4.09e-20
C1211 p[14] _44_/a_93_21# 2.82e-20
C1212 net12 net17 2.11e-21
C1213 _31_/a_285_297# b[1] 0.0101f
C1214 _42_/a_296_53# net3 1.81e-19
C1215 input3/a_27_47# _42_/a_109_93# 0.00249f
C1216 _53_/a_29_53# _09_ 0.00642f
C1217 _33_/a_109_93# p[7] 4.69e-19
C1218 output19/a_27_47# input14/a_27_47# 0.0101f
C1219 _48_/a_109_47# b[1] 9.32e-20
C1220 _09_ _05_ 0.0683f
C1221 net13 _07_ 0.00686f
C1222 net6 _39_/a_377_297# 0.00143f
C1223 _11_ _50_/a_27_47# 0.0592f
C1224 output17/a_27_47# _03_ 1.94e-19
C1225 net13 _30_/a_109_53# 1.05e-19
C1226 net12 _30_/a_215_297# 0.00676f
C1227 _18_ _02_ 2.96e-20
C1228 net3 _49_/a_75_199# 2.01e-19
C1229 net11 _26_/a_29_53# 1.08e-20
C1230 _04_ _19_ 0.356f
C1231 VPWR _02_ 0.332f
C1232 _09_ p[7] 6.7e-20
C1233 net3 _44_/a_93_21# 0.0102f
C1234 _43_/a_369_47# _10_ 0.00199f
C1235 net5 _39_/a_47_47# 0.0389f
C1236 net4 _12_ 0.105f
C1237 net15 _49_/a_201_297# 1.41e-19
C1238 input5/a_841_47# net7 0.00193f
C1239 _53_/a_29_53# _06_ 0.0709f
C1240 net16 _45_/a_193_297# 0.00187f
C1241 input2/a_27_47# b[1] 0.014f
C1242 _04_ _08_ 5.99e-19
C1243 net5 _52_/a_250_297# 0.018f
C1244 net14 _19_ 0.0512f
C1245 _06_ _05_ 0.00724f
C1246 p[12] _47_/a_299_297# 8.13e-21
C1247 _21_ _07_ 0.133f
C1248 _55_/a_217_297# net5 8.84e-20
C1249 _21_ _30_/a_109_53# 3.31e-20
C1250 _31_/a_285_297# _02_ 5.86e-20
C1251 p[13] net8 0.00353f
C1252 _06_ p[7] 0.00864f
C1253 _32_/a_27_47# _21_ 8.95e-19
C1254 net12 _12_ 7.94e-21
C1255 VPWR _37_/a_197_47# -3.27e-19
C1256 _26_/a_183_297# _10_ 5.74e-19
C1257 _04_ net12 0.267f
C1258 net4 net14 2.21e-21
C1259 _39_/a_47_47# _00_ 1.85e-20
C1260 net1 _29_/a_29_53# 9.76e-19
C1261 _48_/a_27_47# _08_ 2.58e-19
C1262 _17_ _43_/a_369_47# 5.87e-19
C1263 VPWR _28_/a_109_297# -1.71e-19
C1264 net6 b[3] 0.00152f
C1265 VPWR input12/a_27_47# 0.0646f
C1266 _15_ _12_ 0.00833f
C1267 net1 net17 2.89e-19
C1268 net13 _03_ 0.271f
C1269 _04_ _15_ 3.61e-20
C1270 b[2] b[1] 5.48e-19
C1271 net13 _01_ 0.00228f
C1272 net5 net11 0.0129f
C1273 _38_/a_27_47# net4 0.0119f
C1274 net1 _30_/a_215_297# 0.00375f
C1275 net12 _48_/a_27_47# 0.0126f
C1276 _23_ net18 -4.05e-24
C1277 VPWR _32_/a_197_47# 0.00146f
C1278 VPWR _50_/a_615_93# -5.34e-19
C1279 p[10] net1 1.22e-19
C1280 net13 _22_ 4.63e-20
C1281 _47_/a_81_21# _10_ 0.0061f
C1282 _35_/a_556_47# _07_ 0.00128f
C1283 _29_/a_183_297# _09_ 4.51e-20
C1284 _20_ _40_/a_191_297# 2.07e-20
C1285 net4 _50_/a_223_47# 0.0107f
C1286 _36_/a_27_47# net9 0.00493f
C1287 _54_/a_75_212# VPWR 0.0475f
C1288 _43_/a_27_47# _06_ 0.0329f
C1289 _39_/a_285_47# _02_ 0.0019f
C1290 _33_/a_209_311# _07_ 0.00859f
C1291 VPWR p[5] 0.0962f
C1292 VPWR _29_/a_111_297# -5.85e-19
C1293 net14 _15_ 0.225f
C1294 _13_ _02_ 0.0676f
C1295 p[6] input13/a_27_47# 1.07e-19
C1296 net15 _44_/a_250_297# 8.86e-20
C1297 _21_ _03_ 0.0818f
C1298 _18_ net19 4.89e-20
C1299 _11_ _45_/a_109_297# 0.00168f
C1300 _21_ _01_ 7.94e-19
C1301 input5/a_381_47# _06_ 1.6e-19
C1302 _20_ net13 5.95e-19
C1303 net4 output16/a_27_47# 0.00706f
C1304 net19 VPWR 0.189f
C1305 p[8] p[9] 0.00275f
C1306 _21_ _22_ 0.00314f
C1307 _04_ input5/a_62_47# 0.00345f
C1308 _18_ _32_/a_27_47# 1.18e-20
C1309 VPWR _07_ 0.0728f
C1310 _04_ net1 0.018f
C1311 _42_/a_109_93# _14_ 0.00141f
C1312 b[2] _02_ 2.81e-19
C1313 input4/a_75_212# net4 0.0189f
C1314 VPWR _30_/a_109_53# 9.49e-19
C1315 net10 _50_/a_27_47# 3.78e-21
C1316 _17_ _47_/a_81_21# 0.0456f
C1317 net19 _41_/a_59_75# 3.1e-20
C1318 _32_/a_27_47# VPWR 0.0395f
C1319 _19_ _49_/a_208_47# 7.12e-20
C1320 _23_ _10_ 0.00192f
C1321 _45_/a_193_297# _05_ 4.84e-22
C1322 _15_ _50_/a_223_47# 0.00698f
C1323 _20_ _21_ 0.191f
C1324 net2 _06_ 0.0108f
C1325 net6 _40_/a_109_297# 2.53e-20
C1326 input5/a_62_47# net14 5.28e-20
C1327 net1 net14 6.64e-20
C1328 net15 net8 0.2f
C1329 _06_ _37_/a_27_47# 2.5e-20
C1330 _55_/a_80_21# net3 2.35e-19
C1331 _02_ _50_/a_343_93# 6.94e-19
C1332 net15 _27_/a_277_297# 1.93e-19
C1333 net11 _27_/a_27_297# 1.58e-20
C1334 _48_/a_109_47# _07_ 3.01e-19
C1335 net3 _27_/a_109_297# 5.45e-19
C1336 _16_ _44_/a_250_297# 3.25e-19
C1337 p[14] net3 0.00446f
C1338 net9 _33_/a_109_93# 0.00211f
C1339 _03_ _33_/a_209_311# 8.38e-19
C1340 net19 _44_/a_346_47# 0.00124f
C1341 b[1] _19_ 0.00967f
C1342 output18/a_27_47# _06_ 0.0114f
C1343 _39_/a_47_47# _10_ 0.00824f
C1344 net18 net11 0.00221f
C1345 _10_ _52_/a_250_297# 0.00368f
C1346 net19 input2/a_27_47# 2.9e-23
C1347 net9 _09_ 2.62e-19
C1348 _43_/a_193_413# net8 1.62e-20
C1349 net16 _21_ 1.89e-19
C1350 _18_ _03_ 7.25e-23
C1351 net6 _36_/a_27_47# 5.1e-19
C1352 _18_ _01_ 6.1e-20
C1353 net12 _33_/a_296_53# 1.23e-20
C1354 p[4] input13/a_27_47# 7.37e-20
C1355 b[1] _08_ 0.0127f
C1356 _55_/a_217_297# _10_ 1.43e-19
C1357 input2/a_27_47# _30_/a_109_53# 1.54e-20
C1358 output17/a_27_47# _05_ 1.12e-19
C1359 VPWR _03_ 0.835f
C1360 b[3] net15 0.00302f
C1361 input5/a_558_47# net8 0.00357f
C1362 VPWR _01_ 0.521f
C1363 _18_ _22_ 0.0211f
C1364 net3 input14/a_27_47# 9.36e-19
C1365 _45_/a_27_47# _12_ 0.0867f
C1366 _23_ _35_/a_226_47# 4.21e-19
C1367 VPWR _22_ 1.4f
C1368 net9 _06_ 0.0505f
C1369 net12 b[1] 0.12f
C1370 _13_ _07_ 3.22e-23
C1371 net2 _47_/a_299_297# 1.18e-19
C1372 _16_ net8 0.00624f
C1373 _34_/a_47_47# net11 0.0309f
C1374 _17_ _39_/a_47_47# 1.47e-20
C1375 _55_/a_472_297# _16_ 3.71e-19
C1376 _02_ _19_ 0.213f
C1377 _41_/a_59_75# _22_ 6.24e-22
C1378 _18_ _20_ 0.0151f
C1379 _31_/a_285_297# _03_ 0.00677f
C1380 _31_/a_285_297# _01_ 1.92e-19
C1381 p[11] p[8] 0.0027f
C1382 _38_/a_109_47# VPWR -4.66e-19
C1383 _20_ VPWR 0.34f
C1384 net11 _10_ 0.0109f
C1385 net4 _02_ 0.00376f
C1386 output17/a_27_47# p[0] 2.47e-19
C1387 _15_ b[1] 1.19e-19
C1388 input9/a_75_212# _10_ 5.49e-21
C1389 _02_ _08_ 2.26e-20
C1390 _20_ _41_/a_59_75# 1.78e-20
C1391 _35_/a_226_47# _52_/a_250_297# 2.63e-20
C1392 net14 _44_/a_584_47# 7.2e-19
C1393 net12 _02_ 2.28e-19
C1394 input2/a_27_47# _03_ 2.71e-19
C1395 net13 _05_ 0.192f
C1396 _36_/a_27_47# _35_/a_76_199# 3.22e-19
C1397 _18_ net16 8.17e-21
C1398 p[6] _34_/a_377_297# 6.2e-19
C1399 net16 VPWR 0.518f
C1400 net13 p[7] 0.0137f
C1401 input5/a_381_47# output17/a_27_47# 6.6e-20
C1402 net1 p[3] 0.00629f
C1403 _32_/a_27_47# _50_/a_343_93# 6.48e-20
C1404 net15 _40_/a_109_297# 0.0016f
C1405 net6 _09_ 5.43e-20
C1406 net2 p[8] 0.027f
C1407 _15_ _02_ 0.101f
C1408 _13_ _03_ 1.74e-20
C1409 input5/a_62_47# b[1] 0.0024f
C1410 net1 b[1] 0.0593f
C1411 p[8] _37_/a_27_47# 9.82e-21
C1412 _53_/a_29_53# _21_ 0.00959f
C1413 _13_ _22_ 0.00309f
C1414 _45_/a_465_47# _12_ 0.00211f
C1415 _21_ _05_ 0.0104f
C1416 input8/a_27_47# input9/a_75_212# 3.09e-20
C1417 net11 _35_/a_226_47# 3.21e-19
C1418 _36_/a_27_47# _25_ 2.34e-20
C1419 _11_ _12_ 0.195f
C1420 input4/a_75_212# input15/a_27_47# 1.1e-21
C1421 net6 _06_ 0.308f
C1422 _21_ p[7] 2.29e-21
C1423 net2 output17/a_27_47# 0.0285f
C1424 _04_ input3/a_27_47# 3.55e-19
C1425 _55_/a_217_297# net7 1.04e-19
C1426 _38_/a_303_47# _10_ 7.36e-19
C1427 input4/a_75_212# _45_/a_27_47# 2.18e-20
C1428 net12 input12/a_27_47# 0.0297f
C1429 _20_ _47_/a_384_47# 1.72e-19
C1430 _13_ _20_ 7.38e-21
C1431 _15_ _37_/a_197_47# 3.02e-19
C1432 _18_ p[12] 4.76e-21
C1433 b[2] _22_ 0.0043f
C1434 p[12] VPWR 0.0417f
C1435 _42_/a_209_311# net8 7.7e-21
C1436 _28_/a_109_297# _15_ 0.00346f
C1437 net14 _11_ 5e-19
C1438 input6/a_27_47# b[3] 0.00217f
C1439 p[12] _41_/a_59_75# 0.0547f
C1440 net5 _31_/a_35_297# 2.04e-21
C1441 input3/a_27_47# net14 3.47e-19
C1442 net1 _02_ 0.00251f
C1443 _33_/a_109_93# _35_/a_76_199# 3.08e-19
C1444 net19 net4 2.65e-20
C1445 VPWR p[9] 0.358f
C1446 p[5] net12 0.00294f
C1447 net14 _50_/a_429_93# 6.04e-21
C1448 _01_ _50_/a_343_93# 0.0131f
C1449 _29_/a_111_297# net12 1.21e-19
C1450 net7 net11 1.77e-19
C1451 _41_/a_59_75# p[9] 1.02e-19
C1452 _09_ _35_/a_76_199# 0.047f
C1453 _08_ _07_ 0.348f
C1454 _15_ _50_/a_615_93# 0.00183f
C1455 _22_ _50_/a_343_93# 0.0597f
C1456 net16 _39_/a_285_47# 1.29e-19
C1457 net5 _44_/a_250_297# 3.11e-20
C1458 _33_/a_209_311# _05_ 0.0311f
C1459 net2 _40_/a_191_297# 0.00143f
C1460 _13_ net16 0.0198f
C1461 _42_/a_368_53# net3 3.82e-19
C1462 _29_/a_29_53# net10 1.77e-19
C1463 _38_/a_27_47# _11_ 0.071f
C1464 _33_/a_209_311# p[7] 2.26e-19
C1465 net6 _47_/a_299_297# 3.63e-19
C1466 _48_/a_181_47# b[1] 3.46e-19
C1467 net12 _07_ 0.18f
C1468 net6 _39_/a_129_47# 6.91e-19
C1469 _11_ _50_/a_223_47# 0.0329f
C1470 net17 net10 8.67e-21
C1471 net12 _30_/a_109_53# 4.25e-20
C1472 net13 _30_/a_297_297# 3.27e-20
C1473 _20_ _50_/a_343_93# 0.00826f
C1474 VPWR _53_/a_29_53# 0.00821f
C1475 input1/A p[0] 0.0277f
C1476 _49_/a_75_199# net11 4.49e-19
C1477 _32_/a_27_47# net12 1.52e-19
C1478 net10 _30_/a_215_297# 0.0512f
C1479 _06_ _35_/a_76_199# 0.00425f
C1480 VPWR _05_ 0.118f
C1481 _25_ _09_ 1.49e-19
C1482 p[1] output17/a_27_47# 0.00138f
C1483 net1 input12/a_27_47# 7.44e-20
C1484 input9/a_75_212# input13/a_27_47# 0.00732f
C1485 _43_/a_469_47# _10_ 0.00124f
C1486 _14_ net17 2.4e-20
C1487 _00_ _44_/a_250_297# 6.39e-20
C1488 net5 _39_/a_377_297# 0.00234f
C1489 net19 _15_ 0.166f
C1490 VPWR p[7] 0.0286f
C1491 _19_ _03_ 0.0019f
C1492 _32_/a_27_47# _15_ 1.19e-19
C1493 _42_/a_109_93# net17 3.1e-21
C1494 _01_ _19_ 0.031f
C1495 net1 _32_/a_197_47# 0.00142f
C1496 _29_/a_29_53# _50_/a_27_47# 1.44e-20
C1497 net5 net8 0.48f
C1498 _33_/a_368_53# _06_ 1.7e-19
C1499 _31_/a_285_297# _05_ 6.12e-19
C1500 net3 _47_/a_81_21# 6.66e-19
C1501 VPWR _37_/a_303_47# -3.13e-19
C1502 net6 _45_/a_193_297# 9.84e-20
C1503 _02_ _45_/a_27_47# 0.00449f
C1504 p[10] _42_/a_109_93# 1.82e-21
C1505 _48_/a_181_47# _02_ 3.9e-19
C1506 _23_ _52_/a_93_21# 0.0166f
C1507 _25_ _06_ 0.144f
C1508 VPWR p[0] 0.00739f
C1509 _03_ _08_ 0.0144f
C1510 _35_/a_489_413# _10_ 3.41e-19
C1511 net4 _22_ 0.0866f
C1512 net10 _12_ 7.82e-20
C1513 _04_ net10 0.121f
C1514 _17_ _43_/a_469_47# 0.00177f
C1515 b[0] _12_ 2.61e-20
C1516 net15 _06_ 0.033f
C1517 _20_ _19_ 0.00734f
C1518 _14_ _12_ 1.98e-20
C1519 _00_ net8 3.23e-19
C1520 output18/a_27_47# _21_ 0.00103f
C1521 _18_ _43_/a_27_47# 0.0201f
C1522 net13 net9 0.0311f
C1523 net12 _03_ 0.0268f
C1524 _04_ _14_ 2.04e-21
C1525 p[11] VPWR 0.197f
C1526 net1 _07_ 6.08e-22
C1527 net12 _01_ 1.67e-21
C1528 VPWR _32_/a_303_47# 6.03e-19
C1529 VPWR _43_/a_27_47# 0.0186f
C1530 _38_/a_109_47# net4 7.32e-19
C1531 input2/a_27_47# _05_ 1.83e-19
C1532 net1 _30_/a_109_53# 0.0297f
C1533 _20_ net4 3.01e-20
C1534 _32_/a_27_47# net1 0.0211f
C1535 net12 _22_ 5.73e-20
C1536 p[13] p[8] 0.00272f
C1537 _20_ _40_/a_297_297# 9.18e-21
C1538 _39_/a_47_47# _52_/a_93_21# 1.44e-20
C1539 _04_ _42_/a_109_93# 5.77e-22
C1540 _48_/a_27_47# net10 0.00377f
C1541 input5/a_381_47# VPWR 8.33e-19
C1542 _52_/a_93_21# _52_/a_250_297# -6.97e-22
C1543 _43_/a_193_413# _06_ 0.0138f
C1544 _13_ _53_/a_29_53# 9.05e-19
C1545 p[6] p[4] 0.00747f
C1546 _01_ _15_ 0.007f
C1547 _15_ _03_ 7.39e-20
C1548 net14 _14_ 0.184f
C1549 _50_/a_27_47# _12_ 0.00354f
C1550 input3/a_27_47# b[1] 2.97e-19
C1551 VPWR _29_/a_183_297# -8.13e-19
C1552 _04_ _50_/a_27_47# 2.07e-21
C1553 _13_ _05_ 2.57e-20
C1554 _20_ net12 0.00437f
C1555 _21_ net9 0.0282f
C1556 _15_ _22_ 0.0236f
C1557 input5/a_558_47# _06_ 3.55e-19
C1558 _31_/a_285_47# net8 0.00129f
C1559 p[13] output17/a_27_47# 0.00118f
C1560 _42_/a_109_93# net14 0.00351f
C1561 _55_/a_80_21# _55_/a_217_297# 1.42e-32
C1562 net4 net16 0.155f
C1563 input8/a_27_47# _49_/a_201_297# 2.46e-21
C1564 _18_ net2 0.00181f
C1565 _53_/a_29_53# b[2] 6.22e-19
C1566 VPWR _30_/a_297_297# -5.22e-19
C1567 net8 _27_/a_27_297# 0.0108f
C1568 _35_/a_226_47# _49_/a_201_297# 1.66e-20
C1569 net2 VPWR 0.955f
C1570 _16_ _06_ 0.00162f
C1571 _18_ _37_/a_27_47# 3.31e-20
C1572 net15 _47_/a_299_297# 1.44e-20
C1573 _39_/a_47_47# net3 1.66e-20
C1574 _20_ _15_ 0.691f
C1575 _36_/a_27_47# _26_/a_29_53# 1.6e-19
C1576 VPWR _37_/a_27_47# -0.0178f
C1577 p[2] _31_/a_285_47# 4.11e-20
C1578 net11 _52_/a_93_21# 2.8e-19
C1579 net6 _40_/a_191_297# 1.16e-20
C1580 net1 _03_ 0.298f
C1581 _02_ _11_ 0.0621f
C1582 net19 input15/a_27_47# 0.00236f
C1583 net1 _01_ 0.0509f
C1584 _55_/a_300_47# net15 1.09e-19
C1585 _55_/a_217_297# net3 5.78e-20
C1586 input11/a_27_47# b[1] 0.00688f
C1587 VPWR output18/a_27_47# 0.0689f
C1588 input1/A p[1] 0.0336f
C1589 net3 _27_/a_205_297# 4.37e-19
C1590 net1 _22_ 0.0129f
C1591 _48_/a_181_47# _07_ 5.93e-19
C1592 _38_/a_27_47# _50_/a_27_47# 2.37e-20
C1593 _07_ _45_/a_27_47# 1.02e-20
C1594 output16/a_27_47# b[0] 0.014f
C1595 net9 _33_/a_209_311# 4.33e-20
C1596 _13_ _43_/a_27_47# 1.66e-20
C1597 _50_/a_27_47# _50_/a_223_47# 2.84e-32
C1598 net6 net13 0.00188f
C1599 _39_/a_377_297# _10_ 7.42e-19
C1600 net4 p[12] 0.00758f
C1601 net7 _49_/a_201_297# 0.00419f
C1602 _10_ _52_/a_256_47# 1.65e-19
C1603 input8/a_27_47# _31_/a_35_297# 0.00955f
C1604 _20_ net1 0.363f
C1605 net2 _44_/a_346_47# 1.64e-19
C1606 _17_ _44_/a_250_297# 0.0336f
C1607 _18_ net9 1.51e-19
C1608 _55_/a_472_297# _10_ 7.35e-21
C1609 net8 _10_ 5.86e-19
C1610 net2 input2/a_27_47# 0.024f
C1611 VPWR net9 0.465f
C1612 _28_/a_109_297# _11_ 6.29e-19
C1613 _33_/a_296_53# net10 8.22e-20
C1614 input5/a_664_47# net8 0.0116f
C1615 input1/a_75_212# net7 3.77e-19
C1616 VPWR p[1] 0.0919f
C1617 net15 p[8] 1.73e-20
C1618 net6 _21_ 2.92e-20
C1619 _36_/a_27_47# net5 0.0163f
C1620 _45_/a_109_297# _12_ 0.00587f
C1621 input6/a_27_47# _06_ 2.85e-19
C1622 net10 p[3] 0.00107f
C1623 b[1] net10 0.117f
C1624 _53_/a_111_297# _02_ 9.57e-20
C1625 p[12] _15_ 0.0163f
C1626 net4 _53_/a_29_53# 3.26e-19
C1627 _54_/a_75_212# _11_ 3.22e-20
C1628 _03_ _45_/a_27_47# 2.06e-20
C1629 input10/a_27_47# VPWR 0.00986f
C1630 b[3] _10_ 6.63e-21
C1631 _14_ b[1] 1.1e-19
C1632 _31_/a_35_297# net7 0.0384f
C1633 _17_ net8 4.52e-20
C1634 _42_/a_209_311# _06_ 1.66e-19
C1635 _09_ _24_ 0.0202f
C1636 _15_ p[9] 2.06e-19
C1637 _08_ _05_ 0.00897f
C1638 net13 _35_/a_76_199# 0.0337f
C1639 _22_ _45_/a_27_47# 0.0131f
C1640 _42_/a_109_93# b[1] 2.38e-19
C1641 net19 _11_ 2.19e-19
C1642 input8/a_27_47# net8 0.0181f
C1643 net19 input3/a_27_47# 0.00105f
C1644 _06_ _26_/a_29_53# 0.0135f
C1645 p[13] input1/A 1.88e-19
C1646 net12 _05_ 0.0414f
C1647 _32_/a_27_47# _11_ 1.65e-20
C1648 _31_/a_35_297# _49_/a_75_199# 6.24e-19
C1649 output18/a_27_47# b[2] 0.0141f
C1650 output19/a_27_47# _44_/a_250_297# 6.42e-20
C1651 input2/a_27_47# p[1] 0.0125f
C1652 _02_ net10 6.74e-19
C1653 _06_ _24_ 0.113f
C1654 net13 _33_/a_368_53# 2.1e-20
C1655 net12 p[7] 0.042f
C1656 net15 _40_/a_191_297# 8.41e-19
C1657 _17_ b[3] 7.54e-20
C1658 _21_ _35_/a_76_199# 0.0175f
C1659 net2 _50_/a_343_93# 1.25e-20
C1660 input8/a_27_47# p[2] 0.016f
C1661 net13 _25_ 0.00297f
C1662 _14_ _02_ 0.0316f
C1663 _18_ net6 0.166f
C1664 p[6] net11 0.01f
C1665 input11/a_27_47# p[5] 0.0433f
C1666 _29_/a_29_53# _30_/a_215_297# 1.72e-19
C1667 net5 _09_ 5.18e-19
C1668 net6 VPWR 1f
C1669 net13 net15 8.84e-19
C1670 _44_/a_93_21# _44_/a_250_297# -6.97e-22
C1671 p[13] VPWR 0.197f
C1672 _36_/a_109_47# _25_ 3.76e-21
C1673 net6 _41_/a_59_75# 0.0373f
C1674 net17 _30_/a_215_297# 4.69e-20
C1675 net14 _37_/a_109_47# 1.71e-19
C1676 net16 _45_/a_27_47# 8.68e-19
C1677 p[10] net17 0.179f
C1678 net7 net8 0.295f
C1679 _02_ _50_/a_27_47# 2.09e-19
C1680 _21_ _25_ 0.00164f
C1681 net10 input12/a_27_47# 0.00182f
C1682 _00_ _09_ 9.35e-21
C1683 net5 _06_ 0.41f
C1684 p[2] net7 0.0139f
C1685 _28_/a_109_297# _14_ 5.66e-19
C1686 p[12] _41_/a_145_75# 0.00339f
C1687 _33_/a_209_311# _35_/a_76_199# 9.95e-21
C1688 net2 _19_ 0.101f
C1689 net1 _05_ 0.151f
C1690 _04_ _29_/a_29_53# 0.0408f
C1691 _49_/a_75_199# net8 0.00214f
C1692 net14 _50_/a_515_93# 1.39e-20
C1693 net9 _50_/a_343_93# 6.64e-19
C1694 _22_ _11_ 0.15f
C1695 input3/a_27_47# _22_ 5.13e-20
C1696 p[11] _15_ 0.00178f
C1697 net1 p[7] 7.5e-20
C1698 _54_/a_75_212# net10 7.43e-19
C1699 _04_ net17 0.0218f
C1700 _15_ _43_/a_27_47# 8.96e-20
C1701 _00_ _06_ 0.1f
C1702 p[5] net10 0.00544f
C1703 p[12] input15/a_27_47# 5.48e-19
C1704 _36_/a_27_47# _10_ 0.00109f
C1705 net2 _40_/a_297_297# 0.00101f
C1706 _17_ _40_/a_109_297# 9.67e-19
C1707 _18_ _35_/a_76_199# 6.82e-21
C1708 output19/a_27_47# b[3] 0.028f
C1709 _29_/a_29_53# net14 1.61e-20
C1710 _04_ _30_/a_215_297# 0.00225f
C1711 p[2] _49_/a_75_199# 1.72e-19
C1712 _04_ p[10] 8.48e-21
C1713 VPWR _35_/a_76_199# -0.00947f
C1714 _20_ _11_ 0.268f
C1715 input15/a_27_47# p[9] 0.0192f
C1716 net13 _30_/a_392_297# 6.64e-20
C1717 net12 _30_/a_297_297# 7.14e-21
C1718 _52_/a_584_47# _06_ 0.00218f
C1719 net6 _39_/a_285_47# 1.53e-19
C1720 p[4] net11 0.0557f
C1721 net14 net17 5.43e-19
C1722 net6 _13_ 0.0106f
C1723 net10 _07_ 0.0605f
C1724 net10 _30_/a_109_53# 5.6e-20
C1725 net5 _47_/a_299_297# 0.00198f
C1726 net5 _39_/a_129_47# 0.00344f
C1727 net19 _14_ 0.00714f
C1728 _32_/a_27_47# net10 2.76e-20
C1729 net18 _09_ 1.97e-21
C1730 b[3] _44_/a_93_21# 7.01e-20
C1731 p[10] net14 1.59e-20
C1732 VPWR _33_/a_368_53# -4.26e-19
C1733 input5/a_62_47# p[11] 0.00153f
C1734 net5 _52_/a_346_47# 7.03e-19
C1735 net1 _32_/a_303_47# 1.45e-19
C1736 _04_ _12_ 1.42e-19
C1737 _29_/a_29_53# _50_/a_223_47# 1.45e-20
C1738 net2 _15_ 9.8e-19
C1739 VPWR _25_ 0.0829f
C1740 net16 _11_ 0.172f
C1741 net19 _42_/a_109_93# 0.0448f
C1742 _15_ _37_/a_27_47# 1.11e-19
C1743 p[1] _19_ 1.05e-19
C1744 _55_/a_80_21# _31_/a_35_297# 5.9e-21
C1745 net4 net9 1.99e-22
C1746 _47_/a_299_297# _00_ 7.59e-21
C1747 _18_ net15 0.0382f
C1748 _39_/a_47_47# _23_ 5.24e-21
C1749 input5/a_381_47# net1 1.27e-19
C1750 _39_/a_129_47# _00_ 1.63e-20
C1751 _53_/a_111_297# _22_ 4.7e-20
C1752 _02_ _45_/a_109_297# 8.44e-19
C1753 net6 _45_/a_205_47# 2.59e-20
C1754 net9 _08_ 7.71e-21
C1755 _23_ _52_/a_250_297# 3.17e-19
C1756 _45_/a_27_47# _05_ 9.34e-23
C1757 net18 _06_ 0.0211f
C1758 VPWR net15 0.62f
C1759 input7/a_27_47# input1/a_75_212# 3.2e-20
C1760 net5 _45_/a_193_297# 0.00935f
C1761 _04_ net14 0.0863f
C1762 _41_/a_59_75# net15 1.16e-20
C1763 net6 _50_/a_343_93# 0.00214f
C1764 _18_ _43_/a_193_413# 0.0413f
C1765 net12 net9 0.0596f
C1766 VPWR _43_/a_193_413# 0.0063f
C1767 _09_ _10_ 0.0222f
C1768 net1 _30_/a_297_297# 7.34e-20
C1769 net2 net1 1.64e-19
C1770 net10 _03_ 0.321f
C1771 input5/a_62_47# net2 0.0197f
C1772 _13_ _35_/a_76_199# 3.01e-21
C1773 _34_/a_47_47# _06_ 0.0391f
C1774 p[12] _11_ 4.25e-21
C1775 _00_ _45_/a_193_297# 4.38e-20
C1776 _38_/a_27_47# _12_ 0.0527f
C1777 input5/a_558_47# VPWR 0.0083f
C1778 _15_ net9 0.00113f
C1779 _43_/a_297_47# _06_ 4.81e-20
C1780 _52_/a_93_21# _52_/a_256_47# -6.6e-20
C1781 _01_ _14_ 0.0193f
C1782 _50_/a_223_47# _12_ 0.00327f
C1783 _23_ net11 0.0461f
C1784 net3 _44_/a_250_297# 0.0088f
C1785 _04_ _50_/a_223_47# 7.89e-22
C1786 _11_ p[9] 1.01e-19
C1787 _18_ _16_ 0.144f
C1788 _14_ _22_ 0.00449f
C1789 _06_ _10_ 1.14f
C1790 input10/a_27_47# net12 0.00115f
C1791 input5/a_664_47# _06_ 3.21e-19
C1792 VPWR _16_ 0.126f
C1793 net5 output17/a_27_47# 5.01e-20
C1794 net13 _26_/a_29_53# 2.23e-20
C1795 input14/a_27_47# _44_/a_250_297# 8.25e-21
C1796 input2/a_27_47# net15 1.61e-19
C1797 _29_/a_29_53# p[3] 3.9e-19
C1798 _55_/a_80_21# net8 1.84e-21
C1799 _20_ net10 3.23e-19
C1800 _42_/a_109_93# _22_ 1.21e-19
C1801 _29_/a_29_53# b[1] 0.0026f
C1802 _33_/a_109_93# _35_/a_226_47# 4.9e-19
C1803 net14 _50_/a_223_47# 5.89e-21
C1804 _20_ _14_ 0.144f
C1805 input4/a_75_212# _12_ 2.09e-20
C1806 _22_ _50_/a_27_47# 0.0276f
C1807 net6 net4 0.713f
C1808 p[3] _30_/a_215_297# 4.95e-19
C1809 _53_/a_29_53# _11_ 2.33e-20
C1810 net17 b[1] 0.0287f
C1811 p[2] _49_/a_315_47# 6.65e-20
C1812 net11 _52_/a_250_297# 1.2e-19
C1813 _35_/a_226_47# _09_ 0.0599f
C1814 net6 _40_/a_297_297# 7.47e-22
C1815 b[2] _25_ 0.0015f
C1816 net1 net9 0.47f
C1817 input5/a_62_47# net9 3.12e-19
C1818 _17_ _06_ 0.0341f
C1819 b[1] _30_/a_215_297# 0.0176f
C1820 _32_/a_109_47# _02_ 3.98e-19
C1821 net3 net8 9.23e-19
C1822 p[10] b[1] 0.103f
C1823 net1 p[1] 0.0295f
C1824 net3 _27_/a_277_297# 2.71e-19
C1825 input5/a_558_47# input2/a_27_47# 2.04e-20
C1826 net2 input15/a_27_47# 0.00296f
C1827 input7/a_27_47# net8 2.03e-21
C1828 _13_ _43_/a_193_413# 5.58e-21
C1829 _21_ _24_ 0.0388f
C1830 p[14] b[3] 0.0976f
C1831 net6 net12 0.00643f
C1832 _39_/a_129_47# _10_ 2.51e-19
C1833 net16 b[0] 0.0306f
C1834 _47_/a_299_297# _10_ 0.0134f
C1835 _34_/a_129_47# net11 0.00242f
C1836 _37_/a_27_47# input15/a_27_47# 3.27e-19
C1837 _29_/a_29_53# _02_ 6.76e-21
C1838 _35_/a_226_47# _06_ 0.00487f
C1839 net2 _44_/a_584_47# 0.0053f
C1840 net5 net13 0.127f
C1841 net6 _36_/a_197_47# 6.94e-20
C1842 _38_/a_27_47# output16/a_27_47# 9.02e-19
C1843 _04_ p[3] 2.63e-20
C1844 p[2] input7/a_27_47# 0.0023f
C1845 input6/a_27_47# VPWR 0.00642f
C1846 net6 _15_ 0.17f
C1847 net17 _02_ 0.0608f
C1848 net7 _09_ 0.00258f
C1849 b[3] net3 2.43e-20
C1850 input5/a_841_47# net8 0.025f
C1851 b[1] _12_ 3.18e-21
C1852 _04_ b[1] 0.0568f
C1853 _02_ _30_/a_215_297# 3.58e-21
C1854 _36_/a_109_47# net5 0.00144f
C1855 net16 _50_/a_27_47# 2.35e-20
C1856 input9/a_75_212# net11 1.1e-20
C1857 b[3] input14/a_27_47# 0.00296f
C1858 _33_/a_109_93# input13/a_27_47# 0.00348f
C1859 input3/a_27_47# p[11] 0.0137f
C1860 _18_ _42_/a_209_311# 3.21e-19
C1861 _17_ _39_/a_129_47# 1.38e-20
C1862 _43_/a_27_47# _11_ 4.27e-19
C1863 _45_/a_193_297# _10_ 0.0047f
C1864 net5 _21_ 0.00784f
C1865 net7 _06_ 0.00447f
C1866 _42_/a_209_311# VPWR -0.00753f
C1867 _53_/a_183_297# _02_ 4.14e-19
C1868 input13/a_27_47# _09_ 1.27e-21
C1869 net14 b[1] 0.00256f
C1870 _08_ _35_/a_76_199# 0.0061f
C1871 _49_/a_75_199# _09_ 2.93e-19
C1872 net19 _37_/a_109_47# 1.16e-20
C1873 _49_/a_544_297# _09_ 2.56e-20
C1874 _48_/a_27_47# b[1] 0.00666f
C1875 _18_ _26_/a_29_53# 5.26e-20
C1876 output19/a_27_47# _06_ 1.53e-19
C1877 _31_/a_117_297# net7 0.00472f
C1878 VPWR _26_/a_29_53# 0.0356f
C1879 _14_ p[9] 2.62e-21
C1880 net12 _35_/a_76_199# 0.0132f
C1881 _04_ _02_ 0.0541f
C1882 _22_ _45_/a_109_297# 0.0426f
C1883 _02_ _12_ 0.265f
C1884 _21_ _00_ 9.26e-20
C1885 _33_/a_368_53# _08_ 5.04e-19
C1886 _06_ _26_/a_111_297# 9e-19
C1887 VPWR _24_ 0.0129f
C1888 p[12] _50_/a_27_47# 1.34e-19
C1889 input5/a_62_47# p[13] 0.0201f
C1890 net15 _19_ 0.00628f
C1891 input13/a_27_47# _06_ 4.89e-19
C1892 p[13] net1 2.13e-19
C1893 p[6] _34_/a_285_47# 3e-19
C1894 _53_/a_29_53# net10 7.88e-22
C1895 net2 _11_ 0.234f
C1896 input3/a_27_47# net2 0.0229f
C1897 net10 _05_ 0.457f
C1898 net14 _02_ 0.00952f
C1899 net4 net15 8.68e-19
C1900 net12 _33_/a_368_53# 2.63e-19
C1901 _48_/a_27_47# _02_ 0.00435f
C1902 net15 _40_/a_297_297# 4.08e-19
C1903 _11_ _37_/a_27_47# 0.0018f
C1904 net3 _40_/a_109_297# 3.14e-19
C1905 net12 _25_ 4.46e-20
C1906 net10 p[7] 5.72e-19
C1907 _35_/a_226_47# _45_/a_193_297# 8.15e-21
C1908 _19_ _43_/a_193_413# 4.85e-21
C1909 _42_/a_209_311# input2/a_27_47# 1e-22
C1910 _29_/a_29_53# _07_ 1.19e-20
C1911 _29_/a_29_53# _30_/a_109_53# 0.0103f
C1912 net19 net17 8.84e-23
C1913 _18_ net5 0.0426f
C1914 _36_/a_197_47# _25_ 2.37e-21
C1915 _44_/a_93_21# _44_/a_256_47# -6.6e-20
C1916 _38_/a_27_47# _02_ 0.00103f
C1917 net5 VPWR 0.613f
C1918 net16 _45_/a_109_297# 5.1e-20
C1919 net17 _30_/a_109_53# 4.18e-20
C1920 net14 _37_/a_197_47# 7e-19
C1921 net19 p[10] 1.26e-21
C1922 _02_ _50_/a_223_47# 2.51e-20
C1923 _21_ net18 0.00215f
C1924 net5 _41_/a_59_75# 2.41e-19
C1925 net13 _34_/a_47_47# 1.68e-19
C1926 net15 _15_ 0.156f
C1927 net6 input15/a_27_47# 0.146f
C1928 b[1] _49_/a_208_47# 2.93e-19
C1929 _18_ _00_ 0.157f
C1930 net6 _45_/a_27_47# 0.021f
C1931 net9 _11_ 5.39e-19
C1932 net4 _16_ 2.73e-20
C1933 _04_ _29_/a_111_297# 9.25e-19
C1934 net13 _10_ 0.00151f
C1935 VPWR _00_ 0.416f
C1936 b[1] _33_/a_296_53# 2.69e-20
C1937 _32_/a_109_47# _01_ 0.00129f
C1938 _13_ _24_ 2.47e-19
C1939 p[11] _14_ 5.39e-21
C1940 _33_/a_109_93# _52_/a_93_21# 2.89e-21
C1941 net14 _50_/a_615_93# 1.69e-20
C1942 _41_/a_59_75# _00_ 2.43e-20
C1943 _14_ _43_/a_27_47# 0.00938f
C1944 _15_ _43_/a_193_413# 4.86e-19
C1945 _04_ net19 2.07e-20
C1946 b[1] p[3] 0.0042f
C1947 _21_ _34_/a_47_47# 8.93e-19
C1948 _07_ _12_ 2.94e-23
C1949 _04_ _07_ 9.74e-20
C1950 _29_/a_29_53# _03_ 0.0414f
C1951 _17_ _40_/a_191_297# 4.35e-19
C1952 _52_/a_584_47# VPWR -9.47e-19
C1953 _09_ _52_/a_93_21# 0.0227f
C1954 _04_ _30_/a_109_53# 9.19e-21
C1955 _29_/a_29_53# _01_ 8.33e-20
C1956 p[11] _42_/a_109_93# 1.48e-19
C1957 _04_ _32_/a_27_47# 1.43e-19
C1958 input5/a_558_47# _15_ 0.00166f
C1959 input5/a_381_47# _14_ 5.68e-20
C1960 b[2] _24_ 1.85e-19
C1961 output19/a_27_47# p[8] 0.00805f
C1962 _29_/a_29_53# _22_ 2.24e-21
C1963 _09_ _49_/a_315_47# 1.11e-20
C1964 _21_ _10_ 0.00421f
C1965 net12 _30_/a_392_297# 2.19e-20
C1966 net13 _30_/a_465_297# 6.36e-20
C1967 net1 net15 7.44e-20
C1968 net17 _03_ 5.1e-19
C1969 _02_ _49_/a_208_47# 0.00193f
C1970 net19 net14 0.148f
C1971 _01_ net17 0.0988f
C1972 input5/a_664_47# _21_ 9.42e-22
C1973 _47_/a_81_21# net8 2.08e-21
C1974 VPWR _31_/a_285_47# -2.91e-19
C1975 input5/a_381_47# _42_/a_109_93# 0.00763f
C1976 _16_ _15_ 0.0607f
C1977 _50_/a_343_93# _26_/a_29_53# 2.61e-19
C1978 _38_/a_27_47# _54_/a_75_212# 2.67e-19
C1979 net7 output17/a_27_47# 0.0018f
C1980 net10 _30_/a_297_297# 1.68e-19
C1981 _03_ _30_/a_215_297# 0.0393f
C1982 net5 _39_/a_285_47# 0.05f
C1983 net5 _47_/a_384_47# 0.00129f
C1984 net2 net10 2.05e-20
C1985 p[10] _03_ 8.74e-20
C1986 VPWR _27_/a_27_297# 0.0329f
C1987 net11 _49_/a_201_297# 1.42e-19
C1988 _48_/a_27_47# _07_ 0.0524f
C1989 _13_ net5 0.0381f
C1990 _06_ _52_/a_93_21# 0.0584f
C1991 _20_ _29_/a_29_53# 0.0111f
C1992 _22_ _30_/a_215_297# 2.46e-21
C1993 _45_/a_27_47# _35_/a_76_199# 2.04e-21
C1994 net2 _14_ 0.0104f
C1995 _55_/a_80_21# _06_ 5.15e-19
C1996 VPWR net18 0.104f
C1997 net13 _35_/a_226_47# 0.00709f
C1998 _20_ net17 4e-20
C1999 b[1] _02_ 0.00718f
C2000 _34_/a_47_47# _33_/a_209_311# 0.017f
C2001 _14_ _37_/a_27_47# 0.00137f
C2002 p[14] _06_ 1.04e-19
C2003 _47_/a_384_47# _00_ 5.15e-20
C2004 net6 _45_/a_465_47# 6.06e-20
C2005 _34_/a_377_297# _06_ 0.00427f
C2006 input5/a_558_47# net1 1.1e-19
C2007 _45_/a_109_297# _05_ 2.79e-22
C2008 net2 _42_/a_109_93# 0.00507f
C2009 _39_/a_285_47# _00_ 1.47e-21
C2010 _53_/a_183_297# _22_ 3.71e-20
C2011 net5 b[2] 7.33e-20
C2012 _20_ _30_/a_215_297# 6.08e-19
C2013 _23_ _52_/a_256_47# 6.66e-19
C2014 _13_ _00_ 3.77e-20
C2015 input11/a_27_47# input10/a_27_47# 5.3e-19
C2016 _42_/a_109_93# _37_/a_27_47# 2.55e-20
C2017 _03_ _12_ 2.76e-20
C2018 net6 _11_ 0.0257f
C2019 _04_ _03_ 0.586f
C2020 net5 _45_/a_205_47# 8.28e-20
C2021 _04_ _01_ 0.119f
C2022 net6 _50_/a_429_93# 6.18e-19
C2023 net3 _06_ 0.0072f
C2024 _22_ _12_ 0.196f
C2025 input3/a_27_47# p[13] 0.00527f
C2026 _04_ _22_ 1.76e-20
C2027 VPWR _34_/a_47_47# 0.0372f
C2028 _21_ _35_/a_226_47# 9.87e-19
C2029 VPWR _43_/a_297_47# -2.11e-19
C2030 net5 _50_/a_343_93# 0.00124f
C2031 _18_ _10_ 0.133f
C2032 net10 net9 0.111f
C2033 net7 net13 1.72e-19
C2034 net15 input15/a_27_47# 0.00325f
C2035 input2/a_27_47# _27_/a_27_297# 1.16e-19
C2036 _18_ input5/a_664_47# 1.09e-20
C2037 net14 _01_ 8.29e-19
C2038 net14 _03_ 1.5e-19
C2039 net4 _26_/a_29_53# 0.00412f
C2040 _38_/a_109_47# _12_ 0.00179f
C2041 VPWR _10_ 0.58f
C2042 b[1] input12/a_27_47# 0.00658f
C2043 input6/a_27_47# _15_ 5.75e-19
C2044 _20_ _12_ 3.9e-19
C2045 input5/a_664_47# VPWR 0.00488f
C2046 _04_ _20_ 0.0677f
C2047 _52_/a_93_21# _52_/a_346_47# -5.12e-20
C2048 net14 _22_ 2.23e-19
C2049 p[12] _50_/a_515_93# 3.12e-21
C2050 _41_/a_59_75# _10_ 0.0172f
C2051 net3 _44_/a_256_47# 0.00101f
C2052 net4 _24_ 8.65e-20
C2053 _43_/a_193_413# input15/a_27_47# 1.62e-20
C2054 input5/a_841_47# _06_ 1.66e-19
C2055 _00_ _50_/a_343_93# 0.102f
C2056 net13 input13/a_27_47# 0.00139f
C2057 net13 _49_/a_75_199# 3.2e-19
C2058 net12 _26_/a_29_53# 6.55e-19
C2059 _54_/a_75_212# b[1] 0.0023f
C2060 net7 _21_ 3e-19
C2061 net13 _49_/a_544_297# 3.43e-19
C2062 p[5] b[1] 0.00724f
C2063 input10/a_27_47# net10 0.00321f
C2064 _20_ net14 8.01e-20
C2065 _42_/a_209_311# _15_ 0.0521f
C2066 _17_ _18_ 0.271f
C2067 _03_ _50_/a_223_47# 1.41e-21
C2068 VPWR _30_/a_465_297# -4.57e-19
C2069 _33_/a_209_311# _35_/a_226_47# 1.31e-19
C2070 _45_/a_193_297# _52_/a_93_21# 6.01e-19
C2071 _38_/a_27_47# _22_ 2.86e-19
C2072 _11_ _35_/a_76_199# 6.99e-22
C2073 _17_ VPWR 0.306f
C2074 net3 _47_/a_299_297# 2.55e-19
C2075 net16 _12_ 0.131f
C2076 net5 _19_ 6.41e-21
C2077 _02_ input12/a_27_47# 1.88e-19
C2078 _44_/a_346_47# _10_ 9.13e-21
C2079 _15_ _26_/a_29_53# 0.00192f
C2080 _22_ _50_/a_223_47# 0.031f
C2081 net19 b[1] 1e-19
C2082 p[3] _30_/a_109_53# 7.23e-19
C2083 _16_ input15/a_27_47# 7.13e-19
C2084 _17_ _41_/a_59_75# 0.00149f
C2085 _38_/a_197_47# _06_ 4.32e-19
C2086 b[2] net18 0.0131f
C2087 input8/a_27_47# VPWR 0.0863f
C2088 _21_ _49_/a_75_199# 6.64e-19
C2089 b[1] _07_ 0.0417f
C2090 b[1] _30_/a_109_53# 0.00655f
C2091 _32_/a_197_47# _02_ 3.78e-19
C2092 net11 net8 1.5e-19
C2093 net4 net5 0.0447f
C2094 input1/A net7 1.36e-19
C2095 _32_/a_27_47# b[1] 6.39e-19
C2096 VPWR _35_/a_226_47# 0.00159f
C2097 input5/a_664_47# input2/a_27_47# 4.47e-21
C2098 p[6] _06_ 3.5e-19
C2099 _20_ _50_/a_223_47# 1.71e-19
C2100 _54_/a_75_212# _02_ 6.6e-20
C2101 _47_/a_384_47# _10_ 3.53e-19
C2102 _39_/a_285_47# _10_ 0.00289f
C2103 _25_ _11_ 7.05e-19
C2104 p[14] p[8] 0.00112f
C2105 _13_ _10_ 0.0621f
C2106 _29_/a_29_53# _05_ 3.79e-20
C2107 net6 net10 1.35e-20
C2108 input8/a_27_47# _31_/a_285_297# 1.04e-19
C2109 net5 net12 0.0674f
C2110 _17_ _44_/a_346_47# 7.2e-19
C2111 net4 _00_ 0.0166f
C2112 p[12] _12_ 6.43e-20
C2113 net6 _36_/a_303_47# 1.25e-19
C2114 input3/a_27_47# net15 6.19e-20
C2115 net15 _11_ 0.145f
C2116 p[2] input9/a_75_212# 5.13e-20
C2117 net19 _02_ 0.0474f
C2118 _01_ _49_/a_208_47# 2.13e-19
C2119 _03_ _49_/a_208_47# 3.86e-19
C2120 net6 _14_ 2.11e-19
C2121 net6 b[0] 2.52e-19
C2122 _38_/a_27_47# net16 0.114f
C2123 net17 _05_ 0.0111f
C2124 _18_ net7 2.58e-20
C2125 _02_ _07_ 0.0083f
C2126 net16 _50_/a_223_47# 4.77e-21
C2127 _02_ _30_/a_109_53# 5.03e-22
C2128 net3 p[8] 1.72e-19
C2129 _36_/a_197_47# net5 0.00254f
C2130 _33_/a_209_311# input13/a_27_47# 5.85e-20
C2131 _32_/a_27_47# _02_ 0.00247f
C2132 _30_/a_215_297# _05_ 0.0453f
C2133 VPWR net7 0.78f
C2134 net5 _15_ 0.0352f
C2135 p[10] _05_ 6e-20
C2136 _03_ p[3] 0.0038f
C2137 _17_ _47_/a_384_47# 1.1e-20
C2138 input14/a_27_47# p[8] 0.0121f
C2139 _17_ _39_/a_285_47# 7.36e-21
C2140 _43_/a_193_413# _11_ 5.45e-19
C2141 _45_/a_205_47# _10_ 6.19e-20
C2142 output19/a_27_47# VPWR 0.0356f
C2143 p[7] _30_/a_215_297# 4.7e-20
C2144 b[1] _03_ 0.0738f
C2145 _42_/a_296_53# VPWR -6.37e-20
C2146 net6 _50_/a_27_47# 0.0428f
C2147 input6/a_27_47# input15/a_27_47# 5.3e-19
C2148 _01_ b[1] 0.00233f
C2149 p[5] input12/a_27_47# 0.00359f
C2150 _36_/a_27_47# _23_ 0.00118f
C2151 _43_/a_369_47# _06_ -2.02e-19
C2152 net16 output16/a_27_47# 0.0101f
C2153 net3 output17/a_27_47# 0.00248f
C2154 _19_ _27_/a_27_297# 0.0819f
C2155 net14 p[9] 1.05e-19
C2156 _22_ b[1] 9.74e-20
C2157 _15_ _00_ 0.207f
C2158 _50_/a_343_93# _10_ 0.0284f
C2159 _31_/a_285_297# net7 0.00227f
C2160 VPWR input13/a_27_47# 0.0696f
C2161 VPWR _49_/a_75_199# 0.0154f
C2162 VPWR _49_/a_544_297# 0.00504f
C2163 _18_ _44_/a_93_21# 0.00485f
C2164 VPWR _26_/a_111_297# -5.92e-20
C2165 _53_/a_29_53# _12_ 3.46e-20
C2166 _16_ _11_ 4.42e-20
C2167 VPWR _44_/a_93_21# 0.005f
C2168 _13_ _35_/a_226_47# 5.62e-21
C2169 _12_ _05_ 2.52e-19
C2170 p[10] p[0] 6.78e-20
C2171 _20_ p[3] 0.00188f
C2172 net13 _52_/a_93_21# 7.21e-19
C2173 _04_ _05_ 0.0352f
C2174 net10 _35_/a_76_199# 0.0226f
C2175 _06_ _26_/a_183_297# 3.16e-19
C2176 input5/a_62_47# net5 0.00329f
C2177 _20_ b[1] 0.00465f
C2178 net5 net1 0.0772f
C2179 _04_ p[7] 0.00391f
C2180 p[11] p[10] 0.0074f
C2181 _02_ _03_ 0.00474f
C2182 input5/a_381_47# net17 1.37e-20
C2183 input2/a_27_47# net7 0.00213f
C2184 _53_/a_29_53# _48_/a_27_47# 3.14e-21
C2185 _01_ _02_ 0.106f
C2186 net3 _40_/a_191_297# 1.89e-19
C2187 _17_ _50_/a_343_93# 0.0015f
C2188 _31_/a_35_297# _49_/a_201_297# 5.52e-20
C2189 _22_ _02_ 0.552f
C2190 _33_/a_368_53# net10 0.00171f
C2191 _21_ _52_/a_93_21# 9.4e-19
C2192 net1 _00_ 9.43e-19
C2193 _45_/a_27_47# _24_ 4.57e-19
C2194 input4/a_75_212# p[12] 0.02f
C2195 _25_ net10 2.66e-19
C2196 _15_ _27_/a_27_297# 9.85e-20
C2197 _47_/a_81_21# _06_ 0.0388f
C2198 net13 net3 3.25e-21
C2199 _38_/a_27_47# _53_/a_29_53# 1.29e-19
C2200 _34_/a_47_47# _08_ 0.00123f
C2201 input5/a_664_47# _19_ 2.19e-21
C2202 _36_/a_303_47# _25_ 2.03e-21
C2203 _38_/a_109_47# _02_ 1.63e-19
C2204 _44_/a_93_21# _44_/a_346_47# -5.12e-20
C2205 _20_ _02_ 0.1f
C2206 net2 net17 0.261f
C2207 net14 _37_/a_303_47# 0.00112f
C2208 _43_/a_27_47# _12_ 2.33e-21
C2209 net4 _10_ 0.183f
C2210 _21_ _34_/a_377_297# 2.37e-19
C2211 _30_/a_215_297# _30_/a_297_297# -8.88e-34
C2212 _23_ _09_ 0.207f
C2213 _08_ _10_ 1.51e-19
C2214 net12 _34_/a_47_47# 0.0385f
C2215 _32_/a_27_47# _30_/a_109_53# 1.51e-19
C2216 _36_/a_27_47# net11 0.0717f
C2217 net15 _14_ 0.0538f
C2218 p[10] net2 0.0334f
C2219 net6 _45_/a_109_297# 7.82e-19
C2220 _32_/a_109_47# net9 6.44e-19
C2221 net12 _10_ 0.00257f
C2222 _04_ _29_/a_183_297# 0.0015f
C2223 _17_ _19_ 8.82e-21
C2224 p[11] net14 1.9e-19
C2225 net14 _43_/a_27_47# 4.87e-20
C2226 _32_/a_197_47# _01_ 0.00156f
C2227 _42_/a_109_93# net15 4.62e-19
C2228 net5 _45_/a_27_47# 0.0288f
C2229 net1 _27_/a_27_297# 6.05e-21
C2230 _33_/a_109_93# _52_/a_250_297# 5.17e-22
C2231 _23_ _06_ 0.218f
C2232 net16 _02_ 8.94e-19
C2233 _54_/a_75_212# _03_ 5.45e-21
C2234 _14_ _43_/a_193_413# 0.0297f
C2235 _39_/a_47_47# _09_ 7.7e-21
C2236 _17_ net4 7.52e-21
C2237 net8 _49_/a_201_297# 7.3e-19
C2238 _36_/a_197_47# _10_ 1.54e-19
C2239 input5/a_381_47# net14 0.00479f
C2240 _20_ _28_/a_109_297# 0.00221f
C2241 input3/a_27_47# _42_/a_209_311# 1.56e-19
C2242 _29_/a_29_53# net9 0.0205f
C2243 _29_/a_111_297# _03_ 7.48e-19
C2244 net2 _12_ 1.02e-20
C2245 _09_ _52_/a_250_297# 1.97e-20
C2246 _15_ _10_ 0.479f
C2247 _04_ net2 0.158f
C2248 input5/a_664_47# _15_ 9.15e-22
C2249 _18_ _52_/a_93_21# 1.97e-19
C2250 _11_ _26_/a_29_53# 1.09e-19
C2251 _00_ _45_/a_27_47# 4.84e-20
C2252 VPWR _52_/a_93_21# -0.00838f
C2253 net17 net9 1.26e-20
C2254 p[2] _49_/a_201_297# 5.28e-20
C2255 net12 _30_/a_465_297# 8.01e-20
C2256 _18_ _55_/a_80_21# 1.44e-20
C2257 net19 _01_ 4.9e-19
C2258 input5/a_841_47# _21_ 1.59e-21
C2259 _20_ _50_/a_615_93# 8.8e-19
C2260 _16_ _14_ 0.0584f
C2261 _39_/a_47_47# _06_ 1.44e-19
C2262 input7/a_27_47# input1/A 5.13e-20
C2263 _03_ _30_/a_109_53# 0.0189f
C2264 net10 _30_/a_392_297# 3.4e-19
C2265 input5/a_558_47# _42_/a_109_93# 1.75e-19
C2266 net9 _30_/a_215_297# 0.0426f
C2267 VPWR _49_/a_315_47# 3.4e-19
C2268 _03_ _07_ 0.0113f
C2269 _55_/a_80_21# VPWR 0.0289f
C2270 p[1] net17 8.02e-19
C2271 _32_/a_27_47# _03_ 1.9e-19
C2272 net19 _22_ 2.17e-19
C2273 _08_ _35_/a_226_47# 0.00117f
C2274 _33_/a_296_53# _05_ 4.53e-19
C2275 _11_ _24_ 7.29e-20
C2276 _06_ _52_/a_250_297# 0.0058f
C2277 VPWR _27_/a_109_297# -2.45e-19
C2278 _32_/a_27_47# _01_ 0.0266f
C2279 net11 _33_/a_109_93# 5.14e-19
C2280 net2 net14 0.151f
C2281 p[14] VPWR 0.0379f
C2282 _22_ _07_ 1.19e-20
C2283 _22_ _30_/a_109_53# 3.67e-21
C2284 p[10] p[1] 7.02e-19
C2285 p[3] _05_ 7.24e-20
C2286 VPWR _34_/a_377_297# -0.00192f
C2287 _32_/a_27_47# _22_ 1.76e-19
C2288 _55_/a_217_297# _06_ 3.46e-19
C2289 net14 _37_/a_27_47# 0.0584f
C2290 _53_/a_29_53# b[1] 4.99e-19
C2291 p[14] _41_/a_59_75# 5.13e-20
C2292 _17_ _15_ 0.0752f
C2293 net11 _09_ 0.0262f
C2294 net12 _35_/a_226_47# 8.29e-19
C2295 net1 _10_ 4.34e-19
C2296 net7 _19_ 0.0458f
C2297 b[1] _05_ 0.0316f
C2298 _18_ net3 7.34e-20
C2299 net19 _20_ 1.29e-19
C2300 _31_/a_35_297# net8 0.0408f
C2301 p[3] p[7] 0.0273f
C2302 _34_/a_129_47# _06_ 5.3e-19
C2303 input5/a_664_47# net1 2.41e-19
C2304 _20_ _07_ 1.28e-21
C2305 VPWR net3 0.351f
C2306 b[1] p[7] 0.00465f
C2307 _20_ _30_/a_109_53# 8.12e-19
C2308 _54_/a_75_212# net16 1.69e-21
C2309 input7/a_27_47# VPWR 0.0768f
C2310 _32_/a_27_47# _20_ 0.0069f
C2311 p[6] _21_ 0.00232f
C2312 net9 _12_ 4.39e-22
C2313 _04_ net9 0.0206f
C2314 VPWR input14/a_27_47# 0.0739f
C2315 net7 _08_ 9.54e-25
C2316 net6 _50_/a_515_93# 4.7e-19
C2317 _04_ p[1] 6.01e-20
C2318 p[2] _31_/a_35_297# 0.00272f
C2319 net11 _06_ 0.546f
C2320 net5 _11_ 0.207f
C2321 _49_/a_75_199# _19_ 0.0206f
C2322 _38_/a_27_47# output18/a_27_47# 8.6e-19
C2323 _53_/a_29_53# _02_ 0.0388f
C2324 b[1] p[0] 2.85e-19
C2325 net14 net9 7.12e-20
C2326 net7 net12 1.57e-19
C2327 _01_ _03_ 2.85e-19
C2328 net6 _29_/a_29_53# 1.4e-20
C2329 _23_ _45_/a_193_297# 4.13e-19
C2330 _02_ _05_ 0.00163f
C2331 _13_ _52_/a_93_21# 1.31e-19
C2332 input6/a_27_47# _14_ 3.75e-21
C2333 input5/a_841_47# VPWR 0.0775f
C2334 _53_/a_111_297# _24_ 9.08e-21
C2335 p[1] net14 0.0025f
C2336 _22_ _03_ 2.55e-20
C2337 _01_ _22_ 0.15f
C2338 p[11] b[1] 2.45e-20
C2339 _00_ _11_ 0.238f
C2340 _41_/a_145_75# _10_ 5.18e-19
C2341 input8/a_27_47# net1 0.0347f
C2342 net7 _15_ 8.4e-20
C2343 net3 _44_/a_346_47# 8.04e-19
C2344 b[3] _44_/a_250_297# 3.33e-19
C2345 net6 _30_/a_215_297# 3.3e-21
C2346 p[4] net13 2.34e-20
C2347 net1 _35_/a_226_47# 1.3e-20
C2348 output18/a_27_47# output16/a_27_47# 7.85e-19
C2349 net12 input13/a_27_47# 0.0163f
C2350 b[2] _52_/a_93_21# 1.63e-19
C2351 input5/a_381_47# b[1] 0.0023f
C2352 _20_ _03_ 0.0794f
C2353 _42_/a_296_53# _15_ 1.28e-19
C2354 _42_/a_209_311# _14_ 0.00142f
C2355 _39_/a_47_47# _45_/a_193_297# 1.4e-20
C2356 _10_ input15/a_27_47# 4.5e-19
C2357 input7/a_27_47# input2/a_27_47# 1.62e-19
C2358 net10 _26_/a_29_53# 3.48e-22
C2359 net8 _27_/a_277_297# 7.99e-20
C2360 net9 _50_/a_223_47# 2e-19
C2361 _20_ _01_ 0.161f
C2362 _45_/a_27_47# _10_ 0.0143f
C2363 p[13] p[10] 0.00177f
C2364 _38_/a_197_47# VPWR -5.24e-19
C2365 _20_ _22_ 0.183f
C2366 net19 p[12] 6.8e-20
C2367 _14_ _26_/a_29_53# 3.67e-19
C2368 _44_/a_584_47# _10_ 1.14e-20
C2369 p[2] net8 0.0127f
C2370 p[6] VPWR 0.0783f
C2371 _15_ _44_/a_93_21# 0.0168f
C2372 net19 p[9] 0.0731f
C2373 _02_ _43_/a_27_47# 1.88e-21
C2374 net6 _12_ 0.0891f
C2375 b[1] _30_/a_297_297# 3.14e-19
C2376 input12/a_27_47# p[7] 1.07e-19
C2377 _32_/a_303_47# _02_ 1.15e-20
C2378 _04_ net6 2.61e-20
C2379 net2 b[1] 0.0389f
C2380 net1 net7 0.0712f
C2381 input5/a_62_47# net7 2.04e-19
C2382 _29_/a_29_53# _35_/a_76_199# 9.88e-19
C2383 _17_ input15/a_27_47# 6.14e-19
C2384 _50_/a_27_47# _26_/a_29_53# 5.56e-19
C2385 _17_ _45_/a_27_47# 1.16e-20
C2386 net16 _22_ 0.00606f
C2387 net6 net14 2.82e-21
C2388 output18/a_27_47# b[1] 9.26e-19
C2389 p[5] p[7] 6.77e-20
C2390 net1 input13/a_27_47# 1.9e-19
C2391 net1 _49_/a_75_199# 0.00799f
C2392 net5 net10 0.0316f
C2393 _38_/a_109_47# net16 4.17e-19
C2394 p[13] net14 1.89e-19
C2395 net1 _49_/a_544_297# 0.00175f
C2396 _35_/a_226_47# _45_/a_27_47# 5.71e-21
C2397 input5/a_62_47# _44_/a_93_21# 5.05e-20
C2398 _30_/a_109_53# _05_ 0.033f
C2399 _36_/a_303_47# net5 0.00256f
C2400 _07_ _05_ 1.21e-19
C2401 _18_ _43_/a_369_47# 1.49e-19
C2402 net5 b[0] 3.39e-19
C2403 _32_/a_27_47# _05_ 2.2e-20
C2404 net13 _23_ 4.11e-19
C2405 net5 _14_ 3.89e-19
C2406 net9 p[3] 0.0375f
C2407 VPWR _43_/a_369_47# -3.75e-19
C2408 _45_/a_465_47# _10_ 3.32e-19
C2409 _42_/a_368_53# VPWR -3.03e-19
C2410 net6 _50_/a_223_47# 0.0194f
C2411 net5 _42_/a_109_93# 0.00109f
C2412 b[1] net9 0.0765f
C2413 _19_ _49_/a_315_47# 1.33e-19
C2414 net4 _52_/a_93_21# 7.93e-20
C2415 _11_ _10_ 0.176f
C2416 p[12] _22_ 2.13e-21
C2417 _19_ _27_/a_109_297# 7.54e-21
C2418 _36_/a_109_47# _23_ 3.44e-19
C2419 _12_ _35_/a_76_199# 6.84e-20
C2420 net15 net17 5.19e-19
C2421 _04_ _35_/a_76_199# 0.0269f
C2422 _35_/a_489_413# _09_ 0.0296f
C2423 p[4] VPWR 0.114f
C2424 output18/a_27_47# _02_ 4.13e-19
C2425 p[1] b[1] 0.00468f
C2426 _09_ _49_/a_201_297# 1.74e-20
C2427 _55_/a_80_21# net4 1.06e-19
C2428 _14_ _00_ 0.133f
C2429 VPWR _26_/a_183_297# -3.03e-19
C2430 net5 _50_/a_27_47# 0.0169f
C2431 _50_/a_429_93# _10_ 0.00167f
C2432 net2 _37_/a_197_47# 4.74e-20
C2433 _21_ _23_ 0.0217f
C2434 p[10] net15 0.00989f
C2435 net6 output16/a_27_47# 1.5e-19
C2436 net19 p[11] 0.00645f
C2437 net3 _19_ 0.0129f
C2438 input4/a_75_212# net6 0.0273f
C2439 input10/a_27_47# b[1] 0.00691f
C2440 _35_/a_489_413# _06_ 9.22e-19
C2441 input7/a_27_47# _19_ 3.12e-21
C2442 _25_ _12_ 1.23e-20
C2443 _17_ _11_ 0.197f
C2444 _00_ _50_/a_27_47# 0.00197f
C2445 _18_ _47_/a_81_21# 7.96e-20
C2446 net4 net3 9.28e-21
C2447 _02_ net9 0.00611f
C2448 _32_/a_27_47# _43_/a_27_47# 2.01e-20
C2449 net19 input5/a_381_47# 0.00173f
C2450 input5/a_558_47# net17 2.88e-21
C2451 _01_ _05_ 5.03e-19
C2452 _03_ _05_ 0.135f
C2453 net3 _40_/a_297_297# 2.54e-19
C2454 VPWR _47_/a_81_21# 0.00889f
C2455 net12 _34_/a_377_297# 0.00251f
C2456 _53_/a_29_53# _22_ 0.00749f
C2457 _36_/a_27_47# net8 1.52e-19
C2458 net15 _12_ 8.14e-21
C2459 _03_ p[7] 2.5e-22
C2460 _04_ net15 0.0569f
C2461 _22_ _05_ 3.33e-21
C2462 _55_/a_80_21# _15_ 0.107f
C2463 _41_/a_59_75# _47_/a_81_21# 1.5e-19
C2464 input5/a_558_47# p[10] 1.09e-19
C2465 net18 net10 3.35e-20
C2466 _14_ _27_/a_27_297# 1.66e-21
C2467 p[14] _15_ 5.32e-19
C2468 _53_/a_111_297# _10_ 2.06e-19
C2469 net13 net11 0.093f
C2470 input9/a_75_212# net13 4.4e-19
C2471 _42_/a_109_93# _27_/a_27_297# 1.35e-20
C2472 _20_ _05_ 6.79e-19
C2473 _54_/a_75_212# output18/a_27_47# 2.28e-19
C2474 net14 net15 1.07f
C2475 _04_ _43_/a_193_413# 5.67e-21
C2476 _43_/a_193_413# _12_ 7.94e-22
C2477 net19 net2 0.599f
C2478 net19 _37_/a_27_47# 0.0105f
C2479 _28_/a_109_297# net9 3.7e-19
C2480 net3 _15_ 0.224f
C2481 _38_/a_27_47# _25_ 5.76e-19
C2482 _34_/a_47_47# net10 0.0507f
C2483 _04_ input5/a_558_47# 1.25e-20
C2484 VPWR _23_ -0.00374f
C2485 p[13] b[1] 0.00201f
C2486 _55_/a_80_21# net1 1.8e-19
C2487 _32_/a_197_47# net9 6.06e-19
C2488 _01_ _43_/a_27_47# 9.77e-20
C2489 _21_ net11 0.586f
C2490 net14 _43_/a_193_413# 1.11e-19
C2491 net16 _53_/a_29_53# 2.04e-20
C2492 _32_/a_303_47# _01_ 8.58e-19
C2493 net5 _45_/a_109_297# 0.0184f
C2494 input9/a_75_212# _21_ 1.17e-21
C2495 p[11] _22_ 3.13e-20
C2496 net10 _10_ 4.45e-19
C2497 _14_ _43_/a_297_47# 9.11e-19
C2498 _38_/a_197_47# net4 7.64e-19
C2499 _22_ _43_/a_27_47# 0.091f
C2500 output19/a_27_47# input3/a_27_47# 4.77e-21
C2501 p[12] p[9] 1.4e-19
C2502 input5/a_558_47# net14 0.0325f
C2503 _36_/a_303_47# _10_ 4.09e-19
C2504 _14_ _10_ 0.0571f
C2505 _18_ _39_/a_47_47# 1.23e-19
C2506 input10/a_27_47# input12/a_27_47# 0.0154f
C2507 _29_/a_111_297# net9 8.06e-21
C2508 _29_/a_183_297# _03_ 7.36e-19
C2509 VPWR _39_/a_47_47# 0.0668f
C2510 net6 _02_ 0.00427f
C2511 _18_ _52_/a_250_297# 1.77e-19
C2512 _00_ _45_/a_109_297# 4.86e-20
C2513 net1 net3 4.25e-20
C2514 p[6] _08_ 7.08e-19
C2515 input5/a_62_47# net3 0.00164f
C2516 _20_ _32_/a_303_47# 1.54e-19
C2517 _20_ _43_/a_27_47# 0.0124f
C2518 _16_ net14 0.00266f
C2519 VPWR _52_/a_250_297# 0.019f
C2520 p[13] _02_ 7.32e-20
C2521 net9 _07_ 1.39e-20
C2522 _39_/a_377_297# _06_ 8.76e-20
C2523 _11_ _44_/a_93_21# 4.78e-20
C2524 _03_ _30_/a_297_297# 0.00117f
C2525 input7/a_27_47# net1 0.0383f
C2526 net10 _30_/a_465_297# 0.00106f
C2527 net9 _30_/a_109_53# 0.0191f
C2528 _55_/a_217_297# VPWR -0.00133f
C2529 _54_/a_75_212# input10/a_27_47# 1.17e-22
C2530 net2 _03_ 1.89e-19
C2531 _32_/a_27_47# net9 0.0136f
C2532 _06_ _52_/a_256_47# 0.00207f
C2533 _50_/a_27_47# _10_ 0.0154f
C2534 p[6] net12 0.0262f
C2535 input10/a_27_47# p[5] 0.0231f
C2536 VPWR _27_/a_205_297# 1.05e-19
C2537 net2 _01_ 2.72e-19
C2538 b[1] _35_/a_76_199# 0.00458f
C2539 net11 _33_/a_209_311# 2.49e-19
C2540 _42_/a_209_311# net17 1.04e-21
C2541 VPWR _34_/a_129_47# -9.47e-19
C2542 net8 _06_ 0.00282f
C2543 _29_/a_29_53# _26_/a_29_53# 0.00121f
C2544 net2 _22_ 1.93e-20
C2545 _17_ _14_ 0.489f
C2546 _45_/a_27_47# _52_/a_93_21# 1.18e-19
C2547 _39_/a_285_47# _23_ 1.9e-20
C2548 _42_/a_209_311# p[10] 2.37e-20
C2549 _31_/a_117_297# net8 5.91e-19
C2550 _34_/a_285_47# _06_ 0.00598f
C2551 input5/a_841_47# net1 1.33e-19
C2552 net10 _35_/a_226_47# 0.018f
C2553 _13_ _23_ 2.08e-20
C2554 _17_ _42_/a_109_93# 7.83e-20
C2555 _47_/a_81_21# _50_/a_343_93# 0.00282f
C2556 VPWR net11 0.996f
C2557 b[1] _33_/a_368_53# 4.19e-19
C2558 _20_ net2 8.83e-19
C2559 output18/a_27_47# _22_ 7.51e-19
C2560 p[14] input15/a_27_47# 7.31e-19
C2561 input9/a_75_212# VPWR 0.0641f
C2562 b[1] _25_ 0.0015f
C2563 _17_ _50_/a_27_47# 3.93e-20
C2564 net6 _50_/a_615_93# 1.43e-19
C2565 _02_ _35_/a_76_199# 5.73e-19
C2566 b[2] _23_ 2.87e-20
C2567 b[3] _06_ 9.96e-21
C2568 net15 b[1] 0.00314f
C2569 net5 _32_/a_109_47# 5.69e-21
C2570 _13_ _39_/a_47_47# 0.00117f
C2571 _03_ net9 0.149f
C2572 input6/a_27_47# net14 7.05e-19
C2573 net3 input15/a_27_47# 8.74e-20
C2574 _04_ _42_/a_209_311# 9.84e-22
C2575 _01_ net9 0.157f
C2576 input1/a_75_212# output17/a_27_47# 0.0101f
C2577 _48_/a_109_47# net11 1.74e-19
C2578 _13_ _52_/a_250_297# 5.43e-19
C2579 net7 net10 1.65e-36
C2580 _22_ net9 0.0023f
C2581 p[6] net1 3.12e-20
C2582 net5 _29_/a_29_53# 8.1e-20
C2583 _26_/a_29_53# _12_ 0.00243f
C2584 net19 net6 0.00352f
C2585 _04_ _26_/a_29_53# 2.3e-21
C2586 p[11] p[9] 0.00566f
C2587 p[7] _05_ 1.93e-19
C2588 net7 _14_ 0.00251f
C2589 p[4] net12 5.33e-19
C2590 _02_ _25_ 0.0156f
C2591 net5 net17 4.21e-21
C2592 output19/a_27_47# _14_ 1.43e-19
C2593 _42_/a_209_311# net14 0.0238f
C2594 _12_ _24_ 1.67e-19
C2595 b[2] _52_/a_250_297# 1.6e-19
C2596 net16 output18/a_27_47# 3.45e-19
C2597 input5/a_558_47# b[1] 0.00214f
C2598 net13 _35_/a_489_413# 7.36e-20
C2599 _20_ net9 0.328f
C2600 net10 input13/a_27_47# 8.86e-20
C2601 net5 _30_/a_215_297# 8.27e-21
C2602 net15 _02_ 0.0806f
C2603 _45_/a_109_297# _10_ 0.00202f
C2604 net5 p[10] 5.12e-21
C2605 _32_/a_27_47# p[13] 6.49e-20
C2606 net14 _26_/a_29_53# 1.33e-20
C2607 net13 _49_/a_201_297# 3.31e-19
C2608 _38_/a_303_47# VPWR -4.83e-19
C2609 output19/a_27_47# _42_/a_109_93# 1.56e-20
C2610 _16_ b[1] 2.21e-19
C2611 _14_ _49_/a_75_199# 6.79e-20
C2612 _15_ _26_/a_183_297# 4.63e-36
C2613 _13_ net11 2.34e-19
C2614 _14_ _44_/a_93_21# 0.04f
C2615 b[1] _30_/a_392_297# 3.99e-19
C2616 _02_ _43_/a_193_413# 9.4e-21
C2617 _40_/a_109_297# _06_ 0.00175f
C2618 _21_ _35_/a_489_413# 0.0448f
C2619 net15 _37_/a_197_47# 1.78e-19
C2620 net2 p[9] 0.00112f
C2621 b[2] net11 1.46e-19
C2622 _42_/a_109_93# _44_/a_93_21# 1.25e-19
C2623 net5 _12_ 0.983f
C2624 _50_/a_223_47# _26_/a_29_53# 0.00124f
C2625 _17_ _45_/a_109_297# 4.29e-22
C2626 _04_ net5 0.00476f
C2627 _37_/a_27_47# p[9] 0.0117f
C2628 _15_ _47_/a_81_21# 0.00332f
C2629 net6 _03_ 2.9e-20
C2630 _07_ _35_/a_76_199# 0.00226f
C2631 _23_ _08_ 1.81e-19
C2632 net3 _11_ 0.165f
C2633 _16_ _02_ 0.00564f
C2634 _31_/a_35_297# net13 1.86e-20
C2635 _54_/a_75_212# _25_ 0.0247f
C2636 input3/a_27_47# net3 0.03f
C2637 net6 _22_ 0.163f
C2638 output17/a_27_47# net8 0.0043f
C2639 net17 _31_/a_285_47# 0.00134f
C2640 _35_/a_226_47# _45_/a_109_297# 1.59e-21
C2641 _36_/a_27_47# _06_ 0.0501f
C2642 p[13] _01_ 2.02e-20
C2643 input14/a_27_47# _11_ 1.42e-19
C2644 net5 net14 0.0263f
C2645 _00_ _12_ 0.00396f
C2646 _04_ _00_ 1.98e-20
C2647 net17 _27_/a_27_297# 0.00181f
C2648 input3/a_27_47# input14/a_27_47# 5.08e-20
C2649 _18_ _43_/a_469_47# 1.59e-19
C2650 b[3] p[8] 0.00229f
C2651 net12 _23_ 2.28e-21
C2652 net2 _05_ 4.03e-20
C2653 VPWR _43_/a_469_47# -2.75e-19
C2654 net4 _39_/a_47_47# 0.0202f
C2655 _33_/a_209_311# _35_/a_489_413# 2.77e-20
C2656 p[10] _27_/a_27_297# 1.63e-19
C2657 net6 _20_ 9.69e-20
C2658 net4 _52_/a_250_297# 0.00136f
C2659 _04_ _52_/a_584_47# 2.5e-19
C2660 net14 _00_ 4.11e-20
C2661 _53_/a_29_53# output18/a_27_47# 9.46e-19
C2662 _38_/a_27_47# net5 1.76e-19
C2663 net1 _47_/a_81_21# 1.58e-21
C2664 net19 net15 0.0501f
C2665 input1/A input1/a_75_212# 0.0172f
C2666 _35_/a_226_297# _09_ 4.98e-19
C2667 _55_/a_217_297# net4 1.13e-19
C2668 _33_/a_109_93# _09_ 7.36e-20
C2669 _16_ _28_/a_109_297# 1.26e-19
C2670 net5 _50_/a_223_47# 0.00202f
C2671 _50_/a_515_93# _10_ 0.00129f
C2672 net2 _37_/a_303_47# 4.41e-19
C2673 _17_ _37_/a_109_47# 8.86e-21
C2674 VPWR _35_/a_489_413# -0.00725f
C2675 _42_/a_209_311# b[1] 5.21e-19
C2676 VPWR _49_/a_201_297# 0.0175f
C2677 _29_/a_29_53# _10_ 5.17e-19
C2678 net6 net16 8.27e-20
C2679 _04_ _27_/a_27_297# 0.0526f
C2680 _01_ _35_/a_76_199# 3.08e-21
C2681 _03_ _35_/a_76_199# 0.0733f
C2682 net19 _43_/a_193_413# 3.31e-19
C2683 _34_/a_129_47# _08_ 3.29e-19
C2684 _19_ net11 6.27e-21
C2685 net10 _52_/a_93_21# 7.84e-20
C2686 _35_/a_226_297# _06_ 1.28e-19
C2687 net5 output16/a_27_47# 4.14e-19
C2688 b[1] _26_/a_29_53# 9.93e-21
C2689 net13 net8 7.51e-20
C2690 _00_ _50_/a_223_47# 0.00738f
C2691 net18 _12_ 8.24e-19
C2692 _22_ _35_/a_76_199# 6.58e-21
C2693 _33_/a_109_93# _06_ 6.96e-19
C2694 p[11] net2 0.00557f
C2695 net19 input5/a_558_47# 2.24e-20
C2696 net9 _05_ 0.124f
C2697 net2 _43_/a_27_47# 0.01f
C2698 input4/a_75_212# net5 0.0104f
C2699 input1/a_75_212# VPWR 0.0786f
C2700 net13 _34_/a_285_47# 4.11e-20
C2701 b[1] _24_ 2.68e-19
C2702 _30_/a_215_297# _10_ 5.66e-20
C2703 net11 _08_ 8.83e-19
C2704 net9 p[7] 8.26e-19
C2705 net14 _27_/a_27_297# 0.0118f
C2706 _55_/a_217_297# _15_ 0.0474f
C2707 _55_/a_80_21# _14_ 0.0175f
C2708 _09_ _06_ 0.0965f
C2709 input5/a_381_47# net2 0.0138f
C2710 net10 _34_/a_377_297# 1.62e-19
C2711 _20_ _35_/a_76_199# 3.21e-20
C2712 _25_ _03_ 0.00422f
C2713 _15_ _27_/a_205_297# 5.5e-20
C2714 net19 _16_ 0.206f
C2715 p[14] _14_ 1.66e-20
C2716 _42_/a_209_311# _02_ 9.92e-19
C2717 net12 net11 0.358f
C2718 _21_ net8 0.00656f
C2719 _53_/a_183_297# _10_ 2.86e-19
C2720 _22_ _25_ 5.39e-19
C2721 _04_ _34_/a_47_47# 1.17e-20
C2722 net15 _03_ 4.26e-20
C2723 net6 p[12] 0.0941f
C2724 VPWR _31_/a_35_297# 0.0284f
C2725 _01_ net15 0.0314f
C2726 _02_ _26_/a_29_53# 0.0466f
C2727 _21_ _34_/a_285_47# 6.94e-20
C2728 _12_ _10_ 0.19f
C2729 p[1] p[0] 0.00812f
C2730 _04_ _10_ 9.24e-20
C2731 _29_/a_29_53# _35_/a_226_47# 2.64e-19
C2732 net15 _22_ 2.74e-19
C2733 net3 _14_ 0.0295f
C2734 _38_/a_27_47# net18 0.00997f
C2735 net6 p[9] 0.14f
C2736 _02_ _24_ 0.0232f
C2737 net5 b[1] 0.00349f
C2738 _04_ input5/a_664_47# 6.73e-21
C2739 VPWR _44_/a_250_297# 0.0233f
C2740 net2 _37_/a_27_47# 0.0692f
C2741 _32_/a_303_47# net9 0.00218f
C2742 _48_/a_27_47# _34_/a_47_47# 4.45e-21
C2743 _42_/a_109_93# net3 0.0435f
C2744 net14 _43_/a_297_47# 1.09e-21
C2745 _01_ _43_/a_193_413# 8.16e-19
C2746 _20_ net15 0.0021f
C2747 _22_ _43_/a_193_413# 0.00133f
C2748 net14 _10_ 2.4e-19
C2749 _38_/a_303_47# net4 5.95e-19
C2750 input5/a_558_47# _01_ 3.97e-20
C2751 input5/a_664_47# net14 0.0179f
C2752 input5/a_381_47# net9 3.4e-19
C2753 _48_/a_27_47# _10_ 4.55e-19
C2754 _29_/a_183_297# net9 3.51e-19
C2755 net6 _53_/a_29_53# 2.11e-20
C2756 _17_ _12_ 0.0109f
C2757 net16 _25_ 1.16e-19
C2758 _17_ _04_ 4.34e-19
C2759 _23_ _45_/a_27_47# 1.74e-19
C2760 net19 input6/a_27_47# 0.00586f
C2761 net7 _29_/a_29_53# 6.01e-19
C2762 _16_ _01_ 3.24e-19
C2763 _20_ _43_/a_193_413# 0.00161f
C2764 VPWR _52_/a_256_47# -9.47e-19
C2765 net1 net11 1.13e-19
C2766 input2/a_27_47# _31_/a_35_297# 0.00136f
C2767 _18_ net8 1.15e-21
C2768 net5 _02_ 0.233f
C2769 _38_/a_27_47# _10_ 0.0133f
C2770 _47_/a_299_297# _06_ 0.0174f
C2771 VPWR net8 0.701f
C2772 _55_/a_472_297# VPWR 0.00488f
C2773 _16_ _22_ 3.8e-19
C2774 _03_ _30_/a_392_297# 6.33e-19
C2775 _04_ input8/a_27_47# 2.36e-22
C2776 input9/a_75_212# net1 0.002f
C2777 net7 net17 0.2f
C2778 net9 _30_/a_297_297# 7.53e-19
C2779 net2 net9 3.64e-20
C2780 VPWR _27_/a_277_297# -3.63e-19
C2781 _06_ _52_/a_346_47# 0.0031f
C2782 _35_/a_226_47# _12_ 8.38e-20
C2783 _50_/a_223_47# _10_ 0.0295f
C2784 _04_ _35_/a_226_47# 0.00551f
C2785 _17_ net14 0.104f
C2786 _09_ _45_/a_193_297# 0.00961f
C2787 net2 p[1] 0.00315f
C2788 p[10] net7 0.00479f
C2789 _39_/a_47_47# _45_/a_27_47# 1.31e-19
C2790 VPWR _34_/a_285_47# -0.00233f
C2791 _29_/a_29_53# _49_/a_75_199# 1.28e-19
C2792 _55_/a_300_47# _06_ 2.5e-20
C2793 net19 _42_/a_209_311# 0.0764f
C2794 p[0] VGND 0.106f
C2795 _04_ VGND 0.472f
C2796 net9 VGND 0.717f
C2797 _03_ VGND 0.478f
C2798 net10 VGND 0.869f
C2799 _30_/a_465_297# VGND 6.42e-19
C2800 _30_/a_392_297# VGND 3.41e-19
C2801 _30_/a_297_297# VGND -5.13e-19
C2802 _30_/a_109_53# VGND 0.151f
C2803 _30_/a_215_297# VGND 0.149f
C2804 _05_ VGND 0.906f
C2805 net8 VGND 0.794f
C2806 _31_/a_285_297# VGND 1.12e-20
C2807 _31_/a_117_297# VGND -0.00177f
C2808 _31_/a_35_297# VGND 0.246f
C2809 _32_/a_303_47# VGND -4.83e-19
C2810 _32_/a_197_47# VGND 8.12e-20
C2811 _32_/a_109_47# VGND 1.05e-19
C2812 _32_/a_27_47# VGND 0.198f
C2813 _11_ VGND 0.358f
C2814 _50_/a_615_93# VGND -5.19e-19
C2815 _50_/a_515_93# VGND -4.75e-19
C2816 _50_/a_429_93# VGND 4.71e-19
C2817 _50_/a_343_93# VGND 0.171f
C2818 _50_/a_223_47# VGND 0.157f
C2819 _50_/a_27_47# VGND 0.255f
C2820 _07_ VGND 0.482f
C2821 _06_ VGND 1.88f
C2822 _33_/a_368_53# VGND 2.38e-19
C2823 _33_/a_296_53# VGND -1.43e-19
C2824 _33_/a_209_311# VGND 0.135f
C2825 _33_/a_109_93# VGND 0.145f
C2826 _08_ VGND 0.292f
C2827 net11 VGND 1.25f
C2828 _34_/a_285_47# VGND 0.0144f
C2829 _34_/a_129_47# VGND -8.76e-20
C2830 _34_/a_377_297# VGND -0.00102f
C2831 _34_/a_47_47# VGND 0.288f
C2832 _23_ VGND 0.266f
C2833 p[9] VGND 0.314f
C2834 input15/a_27_47# VGND 0.223f
C2835 _09_ VGND 0.538f
C2836 _35_/a_556_47# VGND 1.95e-19
C2837 _35_/a_226_297# VGND -4.55e-19
C2838 _35_/a_489_413# VGND 0.0246f
C2839 _35_/a_226_47# VGND 0.151f
C2840 _35_/a_76_199# VGND 0.137f
C2841 _24_ VGND 0.127f
C2842 _12_ VGND 1.2f
C2843 _52_/a_584_47# VGND -0.00112f
C2844 _52_/a_346_47# VGND -0.00175f
C2845 _52_/a_256_47# VGND -0.00161f
C2846 _52_/a_250_297# VGND 0.0246f
C2847 _52_/a_93_21# VGND 0.133f
C2848 _10_ VGND 1.75f
C2849 _36_/a_303_47# VGND 8.14e-19
C2850 _36_/a_197_47# VGND -3.75e-19
C2851 _36_/a_109_47# VGND 3.56e-19
C2852 _36_/a_27_47# VGND 0.196f
C2853 p[8] VGND 0.467f
C2854 input14/a_27_47# VGND 0.247f
C2855 _53_/a_183_297# VGND -4.34e-19
C2856 _53_/a_111_297# VGND -2.89e-19
C2857 _53_/a_29_53# VGND 0.163f
C2858 _37_/a_303_47# VGND -1.63e-19
C2859 _37_/a_197_47# VGND -4.58e-19
C2860 _37_/a_109_47# VGND -7.9e-19
C2861 _37_/a_27_47# VGND 0.16f
C2862 p[7] VGND 0.579f
C2863 input13/a_27_47# VGND 0.255f
C2864 net18 VGND 0.463f
C2865 _25_ VGND 0.39f
C2866 _54_/a_75_212# VGND 0.263f
C2867 net4 VGND 0.888f
C2868 _38_/a_303_47# VGND 1.78e-19
C2869 _38_/a_197_47# VGND 2.29e-19
C2870 _38_/a_109_47# VGND 2.3e-19
C2871 _38_/a_27_47# VGND 0.183f
C2872 net19 VGND 0.32f
C2873 _22_ VGND 0.256f
C2874 _14_ VGND 0.454f
C2875 _15_ VGND 0.485f
C2876 _55_/a_300_47# VGND -0.00109f
C2877 _55_/a_472_297# VGND -0.00188f
C2878 _55_/a_217_297# VGND -0.00225f
C2879 _55_/a_80_21# VGND 0.213f
C2880 p[6] VGND 0.365f
C2881 input12/a_27_47# VGND 0.248f
C2882 p[3] VGND 0.449f
C2883 input9/a_75_212# VGND 0.273f
C2884 _39_/a_285_47# VGND 0.0128f
C2885 _39_/a_129_47# VGND -0.00126f
C2886 _39_/a_377_297# VGND -6.28e-19
C2887 _39_/a_47_47# VGND 0.266f
C2888 p[5] VGND 0.398f
C2889 input11/a_27_47# VGND 0.235f
C2890 p[2] VGND 0.43f
C2891 input8/a_27_47# VGND 0.265f
C2892 p[4] VGND 0.717f
C2893 input10/a_27_47# VGND 0.211f
C2894 net7 VGND 0.868f
C2895 p[1] VGND 0.43f
C2896 input7/a_27_47# VGND 0.265f
C2897 p[14] VGND 0.606f
C2898 input6/a_27_47# VGND 0.205f
C2899 net5 VGND 2.03f
C2900 p[13] VGND 0.484f
C2901 input5/a_841_47# VGND 0.187f
C2902 input5/a_664_47# VGND 0.144f
C2903 input5/a_558_47# VGND 0.163f
C2904 input5/a_381_47# VGND 0.107f
C2905 input5/a_62_47# VGND 0.218f
C2906 p[12] VGND 0.72f
C2907 input4/a_75_212# VGND 0.263f
C2908 p[11] VGND 0.395f
C2909 input3/a_27_47# VGND 0.249f
C2910 net2 VGND 1.66f
C2911 p[10] VGND 0.455f
C2912 input2/a_27_47# VGND 0.194f
C2913 net1 VGND 0.849f
C2914 input1/A VGND 0.34f
C2915 VPWR VGND 37.6f
C2916 input1/a_75_212# VGND 0.268f
C2917 b[3] VGND 0.374f
C2918 output19/a_27_47# VGND 0.534f
C2919 b[2] VGND 0.593f
C2920 output18/a_27_47# VGND 0.601f
C2921 _40_/a_297_297# VGND -5.1e-19
C2922 _40_/a_191_297# VGND -9.29e-19
C2923 _40_/a_109_297# VGND -0.00181f
C2924 b[1] VGND 0.945f
C2925 net17 VGND 0.384f
C2926 output17/a_27_47# VGND 0.545f
C2927 _41_/a_145_75# VGND 3.75e-19
C2928 _41_/a_59_75# VGND 0.191f
C2929 b[0] VGND 0.708f
C2930 output16/a_27_47# VGND 0.616f
C2931 _16_ VGND 0.119f
C2932 _42_/a_368_53# VGND -4.05e-19
C2933 _42_/a_209_311# VGND 0.135f
C2934 _42_/a_109_93# VGND 0.153f
C2935 _17_ VGND 0.563f
C2936 _43_/a_369_47# VGND -8.43e-19
C2937 _43_/a_297_47# VGND -1.33e-19
C2938 _43_/a_193_413# VGND 0.122f
C2939 _43_/a_27_47# VGND 0.209f
C2940 _00_ VGND 0.516f
C2941 net6 VGND 1f
C2942 _26_/a_183_297# VGND 2.42e-19
C2943 _26_/a_111_297# VGND -2.75e-19
C2944 _26_/a_29_53# VGND 0.218f
C2945 _01_ VGND 0.244f
C2946 net14 VGND 0.958f
C2947 net3 VGND 0.784f
C2948 net15 VGND 0.673f
C2949 _27_/a_277_297# VGND -4.65e-19
C2950 _27_/a_205_297# VGND -3.36e-19
C2951 _27_/a_109_297# VGND -6.15e-19
C2952 _27_/a_27_297# VGND 0.147f
C2953 _18_ VGND 0.159f
C2954 _44_/a_584_47# VGND -0.00145f
C2955 _44_/a_346_47# VGND -0.00198f
C2956 _44_/a_256_47# VGND -0.00184f
C2957 _44_/a_250_297# VGND 0.0219f
C2958 _44_/a_93_21# VGND 0.128f
C2959 net16 VGND 0.375f
C2960 _13_ VGND 0.496f
C2961 _45_/a_465_47# VGND -8.14e-19
C2962 _45_/a_205_47# VGND -2.47e-19
C2963 _45_/a_193_297# VGND -0.00131f
C2964 _45_/a_109_297# VGND -0.00108f
C2965 _45_/a_27_47# VGND 0.187f
C2966 _28_/a_109_297# VGND -9.87e-19
C2967 net12 VGND 0.861f
C2968 net13 VGND 0.519f
C2969 _29_/a_183_297# VGND 4.41e-19
C2970 _29_/a_111_297# VGND -1.9e-19
C2971 _29_/a_29_53# VGND 0.234f
C2972 _19_ VGND 0.497f
C2973 _47_/a_384_47# VGND -2.05e-19
C2974 _47_/a_299_297# VGND 0.0344f
C2975 _47_/a_81_21# VGND 0.136f
C2976 _48_/a_181_47# VGND 3.03e-19
C2977 _48_/a_109_47# VGND 9.44e-19
C2978 _48_/a_27_47# VGND 0.232f
C2979 _21_ VGND 0.586f
C2980 _20_ VGND 0.707f
C2981 _02_ VGND 2.08f
C2982 _49_/a_315_47# VGND -0.0034f
C2983 _49_/a_208_47# VGND -0.00164f
C2984 _49_/a_544_297# VGND -0.00256f
C2985 _49_/a_201_297# VGND -5.82e-19
C2986 _49_/a_75_199# VGND 0.205f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFRTVB a_n410_n216# a_n250_n130# a_n308_n42# a_250_n42#
X0 a_250_n42# a_n250_n130# a_n308_n42# a_n410_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.5
C0 a_250_n42# a_n308_n42# 0.011f
C1 a_n250_n130# a_n308_n42# 0.0209f
C2 a_250_n42# a_n250_n130# 0.0209f
C3 a_250_n42# a_n410_n216# 0.0852f
C4 a_n308_n42# a_n410_n216# 0.0853f
C5 a_n250_n130# a_n410_n216# 1.48f
.ends

.subckt sky130_fd_pr__pfet_01v8_XQZLDL a_15_n240# w_n211_n459# a_n73_n240# a_n33_n337#
+ VSUBS
X0 a_15_n240# a_n33_n337# a_n73_n240# w_n211_n459# sky130_fd_pr__pfet_01v8 ad=0.696 pd=5.38 as=0.696 ps=5.38 w=2.4 l=0.15
C0 a_15_n240# a_n33_n337# 0.0313f
C1 a_n73_n240# a_15_n240# 0.385f
C2 a_n73_n240# a_n33_n337# 0.0313f
C3 a_15_n240# w_n211_n459# 0.163f
C4 w_n211_n459# a_n33_n337# 0.206f
C5 a_n73_n240# w_n211_n459# 0.0371f
C6 a_15_n240# VSUBS 0.11f
C7 a_n73_n240# VSUBS 0.195f
C8 a_n33_n337# VSUBS 0.139f
C9 w_n211_n459# VSUBS 1.47f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GC6 a_200_n42# w_n396_n261# a_n200_n139# a_n258_n42#
+ VSUBS
X0 a_200_n42# a_n200_n139# a_n258_n42# w_n396_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_200_n42# a_n200_n139# 0.0196f
C1 a_n258_n42# a_200_n42# 0.0134f
C2 a_n258_n42# a_n200_n139# 0.0196f
C3 a_200_n42# w_n396_n261# 0.0498f
C4 w_n396_n261# a_n200_n139# 0.73f
C5 a_n258_n42# w_n396_n261# 0.0269f
C6 a_200_n42# VSUBS 0.0338f
C7 a_n258_n42# VSUBS 0.0488f
C8 a_n200_n139# VSUBS 0.563f
C9 w_n396_n261# VSUBS 1.69f
.ends

.subckt sky130_fd_pr__nfet_01v8_ATLS57 a_15_n200# a_n73_n200# a_n33_n288# a_n141_n374#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n141_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_15_n200# a_n73_n200# 0.321f
C1 a_n33_n288# a_n73_n200# 0.0312f
C2 a_15_n200# a_n33_n288# 0.0312f
C3 a_15_n200# a_n141_n374# 0.233f
C4 a_n73_n200# a_n141_n374# 0.199f
C5 a_n33_n288# a_n141_n374# 0.341f
.ends

.subckt th13 Vp V13 Vin m1_831_275# Vn m1_559_n458#
XXM0 Vn m1_559_n458# Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vn Vin m1_559_n458# m1_831_275# sky130_fd_pr__nfet_01v8_ZFRTVB
XXM2 Vp Vp m1_831_275# Vin Vn sky130_fd_pr__pfet_01v8_XQZLDL
XXM3 V13 Vp m1_831_275# Vp Vn sky130_fd_pr__pfet_01v8_VZ9GC6
XXM4 V13 Vn m1_831_275# Vn sky130_fd_pr__nfet_01v8_ATLS57
C0 Vn m1_831_275# 0.232f
C1 Vin V13 0.0076f
C2 Vp Vin 0.176f
C3 Vin m1_559_n458# 0.181f
C4 V13 m1_831_275# 0.184f
C5 Vp m1_831_275# 0.215f
C6 m1_559_n458# m1_831_275# 0.0183f
C7 Vin m1_831_275# 0.197f
C8 Vn V13 0.0706f
C9 Vp Vn 0.206f
C10 m1_559_n458# Vn 0.152f
C11 Vp V13 0.135f
C12 Vp m1_559_n458# 0.0628f
C13 Vin Vn 0.347f
C14 m1_831_275# 0 1.05f
C15 Vin 0 1.79f
C16 V13 0 0.365f
C17 Vn 0 0.117f
C18 Vp 0 3.98f
C19 m1_559_n458# 0 0.286f
.ends

.subckt sky130_fd_pr__nfet_01v8_DD6SHA a_n33_n130# a_15_n42# a_n175_n182# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n33_n130# a_n73_n42# 0.0209f
C1 a_15_n42# a_n73_n42# 0.0699f
C2 a_15_n42# a_n33_n130# 0.0209f
C3 a_15_n42# a_n175_n182# 0.0637f
C4 a_n73_n42# a_n175_n182# 0.0716f
C5 a_n33_n130# a_n175_n182# 0.314f
.ends

.subckt sky130_fd_pr__pfet_01v8_7DPLFP w_n245_n261# a_n107_n42# a_n49_n139# a_49_n42#
+ VSUBS
X0 a_49_n42# a_n49_n139# a_n107_n42# w_n245_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.49
C0 w_n245_n261# a_n49_n139# 0.221f
C1 a_49_n42# a_n49_n139# 0.00895f
C2 a_n107_n42# a_n49_n139# 0.00895f
C3 w_n245_n261# a_49_n42# 0.0224f
C4 a_n107_n42# w_n245_n261# 0.0224f
C5 a_n107_n42# a_49_n42# 0.0396f
C6 a_49_n42# VSUBS 0.0487f
C7 a_n107_n42# VSUBS 0.0487f
C8 a_n49_n139# VSUBS 0.206f
C9 w_n245_n261# VSUBS 0.876f
.ends

.subckt sky130_fd_pr__pfet_01v8_MDPZBH a_n102_n42# a_44_n42# a_n44_n139# w_n240_n261#
+ VSUBS
X0 a_44_n42# a_n44_n139# a_n102_n42# w_n240_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.44
C0 w_n240_n261# a_n44_n139# 0.208f
C1 a_44_n42# a_n44_n139# 0.00823f
C2 a_n102_n42# a_n44_n139# 0.00823f
C3 w_n240_n261# a_44_n42# 0.0224f
C4 a_n102_n42# w_n240_n261# 0.0224f
C5 a_n102_n42# a_44_n42# 0.0423f
C6 a_44_n42# VSUBS 0.0485f
C7 a_n102_n42# VSUBS 0.0485f
C8 a_n44_n139# VSUBS 0.191f
C9 w_n240_n261# VSUBS 0.858f
.ends

.subckt th06 Vp Vin V06 Vn m1_904_n796#
XXM0 Vin m1_904_n796# Vn Vn sky130_fd_pr__nfet_01v8_DD6SHA
XXM1 Vp Vp Vin m1_904_n796# Vn sky130_fd_pr__pfet_01v8_7DPLFP
XXM2 Vp V06 m1_904_n796# Vp Vn sky130_fd_pr__pfet_01v8_MDPZBH
XXM3 Vn m1_904_n796# V06 Vn sky130_fd_pr__nfet_01v8_MYA4RC
C0 Vin m1_904_n796# 0.203f
C1 Vn m1_904_n796# 0.0382f
C2 Vp m1_904_n796# 0.197f
C3 V06 m1_904_n796# 0.157f
C4 Vn Vin 0.0188f
C5 Vin Vp 0.113f
C6 Vn Vp 0.0214f
C7 Vn V06 0.00141f
C8 V06 Vp 0.06f
C9 Vp 0 1.69f
C10 m1_904_n796# 0 0.495f
C11 V06 0 0.217f
C12 Vn 0 0.286f
C13 Vin 0 0.524f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGAKDL a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
+ VSUBS
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 w_n211_n419# a_15_n200# 0.0336f
C1 a_n33_n297# a_15_n200# 0.0293f
C2 a_n73_n200# a_15_n200# 0.321f
C3 a_n33_n297# w_n211_n419# 0.191f
C4 a_n73_n200# w_n211_n419# 0.0336f
C5 a_n33_n297# a_n73_n200# 0.0293f
C6 a_15_n200# VSUBS 0.164f
C7 a_n73_n200# VSUBS 0.164f
C8 a_n33_n297# VSUBS 0.147f
C9 w_n211_n419# VSUBS 1.14f
.ends

.subckt sky130_fd_pr__nfet_01v8_4X3CDA a_n306_n216# a_n180_n130# a_n238_n42# a_180_n42#
X0 a_180_n42# a_n180_n130# a_n238_n42# a_n306_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.8
C0 a_n238_n42# a_n180_n130# 0.0189f
C1 a_180_n42# a_n180_n130# 0.0189f
C2 a_n238_n42# a_180_n42# 0.0147f
C3 a_180_n42# a_n306_n216# 0.075f
C4 a_n238_n42# a_n306_n216# 0.075f
C5 a_n180_n130# a_n306_n216# 1.1f
.ends

.subckt sky130_fd_pr__pfet_01v8_MWB9BZ a_15_n43# w_n211_n262# a_n73_n43# a_n33_n140#
+ VSUBS
X0 a_15_n43# a_n33_n140# a_n73_n43# w_n211_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.15
C0 w_n211_n262# a_15_n43# 0.0198f
C1 a_n33_n140# a_15_n43# 0.0193f
C2 a_n73_n43# a_15_n43# 0.0715f
C3 a_n33_n140# w_n211_n262# 0.187f
C4 a_n73_n43# w_n211_n262# 0.0198f
C5 a_n33_n140# a_n73_n43# 0.0193f
C6 a_15_n43# VSUBS 0.0453f
C7 a_n73_n43# VSUBS 0.0453f
C8 a_n33_n140# VSUBS 0.143f
C9 w_n211_n262# VSUBS 0.752f
.ends

.subckt sky130_fd_pr__nfet_01v8_L9ESAD a_n175_n190# a_n73_n50# a_n33_n138# a_15_n50#
X0 a_15_n50# a_n33_n138# a_n73_n50# a_n175_n190# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_n73_n50# a_n33_n138# 0.0216f
C1 a_15_n50# a_n33_n138# 0.0216f
C2 a_n73_n50# a_15_n50# 0.0826f
C3 a_15_n50# a_n175_n190# 0.0704f
C4 a_n73_n50# a_n175_n190# 0.0797f
C5 a_n33_n138# a_n175_n190# 0.315f
.ends

.subckt th11 V11 Vin Vn m1_577_n654# Vp m1_705_187#
XXM0 Vn Vp Vn m1_577_n654# Vn sky130_fd_pr__pfet_01v8_XGAKDL
XXM1 Vn Vin m1_577_n654# m1_705_187# sky130_fd_pr__nfet_01v8_4X3CDA
XXM2 m1_705_187# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_MWB9BZ
XXM3 V11 Vp m1_705_187# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM4 Vn Vn m1_705_187# V11 sky130_fd_pr__nfet_01v8_L9ESAD
C0 m1_577_n654# m1_705_187# 0.0258f
C1 V11 Vin 2.69e-19
C2 Vp Vin 0.285f
C3 V11 Vp 0.026f
C4 Vn Vin 0.135f
C5 V11 Vn 0.00327f
C6 Vp Vn 0.0775f
C7 m1_577_n654# Vin 0.213f
C8 m1_577_n654# V11 6.11e-19
C9 m1_577_n654# Vp 0.0405f
C10 m1_577_n654# Vn 0.0457f
C11 Vin m1_705_187# 0.0649f
C12 V11 m1_705_187# 0.376f
C13 Vp m1_705_187# 0.286f
C14 Vn m1_705_187# 0.463f
C15 m1_705_187# 0 0.602f
C16 V11 0 0.404f
C17 Vn 0 0.355f
C18 Vp 0 2.61f
C19 Vin 0 1.27f
C20 m1_577_n654# 0 0.286f
.ends

.subckt sky130_fd_pr__nfet_01v8_42G4RD a_n80_n42# a_n148_n216# a_n33_n130# a_22_n42#
X0 a_22_n42# a_n33_n130# a_n80_n42# a_n148_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_22_n42# a_n80_n42# 0.0604f
C1 a_n80_n42# a_n33_n130# 0.00866f
C2 a_22_n42# a_n33_n130# 0.00866f
C3 a_22_n42# a_n148_n216# 0.0698f
C4 a_n80_n42# a_n148_n216# 0.0698f
C5 a_n33_n130# a_n148_n216# 0.321f
.ends

.subckt sky130_fd_pr__pfet_01v8_DDPLQ8 a_n77_n42# w_n215_n261# a_n33_n139# a_19_n42#
+ VSUBS
X0 a_19_n42# a_n33_n139# a_n77_n42# w_n215_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_n77_n42# a_19_n42# 0.0641f
C1 a_n77_n42# a_n33_n139# 0.0127f
C2 a_19_n42# w_n215_n261# 0.0399f
C3 a_n33_n139# w_n215_n261# 0.181f
C4 a_n77_n42# w_n215_n261# 0.017f
C5 a_n33_n139# a_19_n42# 0.0127f
C6 a_19_n42# VSUBS 0.035f
C7 a_n77_n42# VSUBS 0.05f
C8 a_n33_n139# VSUBS 0.149f
C9 w_n215_n261# VSUBS 0.797f
.ends

.subckt sky130_fd_pr__nfet_01v8_VWP3K3 a_n33_n130# a_15_n42# a_n141_182# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n141_182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_15_n42# a_n73_n42# 0.0699f
C1 a_n73_n42# a_n33_n130# 0.0209f
C2 a_15_n42# a_n33_n130# 0.0209f
C3 a_15_n42# a_n141_182# 0.0643f
C4 a_n73_n42# a_n141_182# 0.0643f
C5 a_n33_n130# a_n141_182# 0.317f
.ends

.subckt sky130_fd_pr__pfet_01v8_LZD9A4 a_n80_n42# a_22_n42# a_n33_n139# w_n218_n261#
+ VSUBS
X0 a_22_n42# a_n33_n139# a_n80_n42# w_n218_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_n80_n42# a_22_n42# 0.0604f
C1 a_n80_n42# a_n33_n139# 0.0084f
C2 a_22_n42# w_n218_n261# 0.0222f
C3 a_n33_n139# w_n218_n261# 0.185f
C4 a_n80_n42# w_n218_n261# 0.0222f
C5 a_n33_n139# a_22_n42# 0.0084f
C6 a_22_n42# VSUBS 0.0474f
C7 a_n80_n42# VSUBS 0.0474f
C8 a_n33_n139# VSUBS 0.149f
C9 w_n218_n261# VSUBS 0.775f
.ends

.subckt sky130_fd_pr__nfet_01v8_VRD6K3 a_n77_n42# a_n145_n214# a_n33_n130# a_19_n42#
X0 a_19_n42# a_n33_n130# a_n77_n42# a_n145_n214# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_19_n42# a_n77_n42# 0.0641f
C1 a_n77_n42# a_n33_n130# 0.0136f
C2 a_19_n42# a_n33_n130# 0.0136f
C3 a_19_n42# a_n145_n214# 0.0677f
C4 a_n77_n42# a_n145_n214# 0.0677f
C5 a_n33_n130# a_n145_n214# 0.32f
.ends

.subckt th04 Vp V04 Vn m1_892_n998# m1_620_n488# Vin
XXM0 m1_892_n998# Vn Vin Vn sky130_fd_pr__nfet_01v8_42G4RD
XXM1 m1_620_n488# Vp Vin m1_892_n998# Vn sky130_fd_pr__pfet_01v8_DDPLQ8
XXM2 Vp m1_620_n488# Vn Vp sky130_fd_pr__nfet_01v8_VWP3K3
XXM3 Vp V04 m1_892_n998# Vp Vn sky130_fd_pr__pfet_01v8_LZD9A4
XXM4 Vn Vn m1_892_n998# V04 sky130_fd_pr__nfet_01v8_VRD6K3
C0 Vp Vn 0.0386f
C1 Vn V04 0.0639f
C2 m1_620_n488# Vn 2.16e-19
C3 Vp V04 0.0462f
C4 m1_620_n488# Vp 0.17f
C5 m1_620_n488# V04 0.00264f
C6 m1_892_n998# Vin 0.463f
C7 Vn Vin 0.0468f
C8 Vp Vin 0.14f
C9 Vin V04 0.00141f
C10 m1_620_n488# Vin 0.0346f
C11 m1_892_n998# Vn 0.1f
C12 Vp m1_892_n998# 0.383f
C13 m1_892_n998# V04 0.13f
C14 m1_620_n488# m1_892_n998# 0.0117f
C15 Vin 0 0.679f
C16 V04 0 0.287f
C17 Vn 0 0.259f
C18 m1_892_n998# 0 0.832f
C19 Vp 0 2.13f
C20 m1_620_n488# 0 0.0632f
.ends

.subckt adc Vin Vp V01 V02 V03 V04 V08 V07 V06 V09 V10 V11 V12 V13 V14 V15 V05 Vn
+ b[1] b[2] b[3] b[0]
Xth02_0 th15_0/Vin V02 Vp th02_0/m1_983_133# th02_0/m1_571_144# Vn th02
Xth09_0 V09 Vin Vn th09_0/m1_485_n505# Vp th09_0/m1_962_372# th09
Xth14_0 V14 th15_0/Vin Vn th14_0/m1_641_n318# Vp th14_0/m1_891_419# th14
Xth07_0 Vin V07 Vp th07_0/m1_808_n892# Vn th07
Xth12_0 Vp V12 Vin th12_0/m1_394_n856# Vn th12_0/m1_529_n42# th12
Xth05_0 Vp V05 Vin th05_0/m1_752_n794# Vn th05
Xth10_0 Vp V10 Vin Vn th10_0/m1_502_n495# th10_0/m1_536_174# th10
Xth03_0 Vp V03 Vin th03_0/m1_890_n844# th03_0/m1_638_n591# Vn th03
Xth01_0 Vp th15_0/Vin V01 th01_0/m1_991_n1219# Vn th01_0/m1_571_n501# th01
Xpreamp_0 Vp Vin th15_0/Vin Vn preamp
Xth15_0 V15 th15_0/Vin th15_0/m1_597_n912# Vp th15_0/m1_849_n157# Vn th15
Xth08_0 Vin V08 th08_0/m1_477_n803# Vp Vn th08
Xtherm_0 b[0] b[2] b[3] V01 V11 V12 V13 V14 V15 V02 V03 V04 V05 V06 V07 V08 V09 V10
+ therm_0/input3/a_27_47# therm_0/_30_/a_297_297# therm_0/_43_/a_369_47# therm_0/net7
+ therm_0/_35_/a_556_47# therm_0/input13/a_27_47# therm_0/_43_/a_469_47# therm_0/_42_/a_368_53#
+ therm_0/_25_ therm_0/_30_/a_215_297# therm_0/_40_/a_191_297# therm_0/output19/a_27_47#
+ therm_0/net19 therm_0/net4 therm_0/_24_ therm_0/input10/a_27_47# therm_0/_18_ therm_0/_10_
+ therm_0/_52_/a_93_21# therm_0/_31_/a_35_297# therm_0/_07_ therm_0/input7/a_27_47#
+ therm_0/_04_ therm_0/output16/a_27_47# therm_0/input9/a_75_212# therm_0/_30_/a_109_53#
+ therm_0/_40_/a_109_297# b[1] therm_0/_42_/a_209_311# therm_0/_44_/a_584_47# therm_0/_27_/a_27_297#
+ therm_0/input1/a_75_212# therm_0/_41_/a_59_75# therm_0/input5/a_62_47# therm_0/_27_/a_277_297#
+ therm_0/net2 therm_0/input14/a_27_47# therm_0/net3 therm_0/_42_/a_296_53# therm_0/input5/a_841_47#
+ therm_0/_31_/a_285_297# therm_0/_47_/a_81_21# therm_0/_35_/a_76_199# V01 therm_0/net14
+ therm_0/_55_/a_217_297# therm_0/input5/a_381_47# therm_0/_27_/a_205_297# therm_0/_13_
+ therm_0/_34_/a_47_47# therm_0/net15 therm_0/_37_/a_109_47# therm_0/_19_ therm_0/input11/a_27_47#
+ therm_0/_23_ therm_0/net12 therm_0/_34_/a_285_47# therm_0/net18 therm_0/_49_/a_75_199#
+ therm_0/_47_/a_384_47# therm_0/net8 therm_0/net6 therm_0/net11 therm_0/_17_ therm_0/input8/a_27_47#
+ therm_0/_33_/a_209_311# therm_0/_09_ therm_0/output17/a_27_47# therm_0/_01_ therm_0/_37_/a_27_47#
+ therm_0/_38_/a_109_47# therm_0/_48_/a_109_47# therm_0/_47_/a_299_297# therm_0/_44_/a_250_297#
+ therm_0/_44_/a_93_21# therm_0/_48_/a_181_47# therm_0/_44_/a_346_47# therm_0/_37_/a_197_47#
+ therm_0/net13 therm_0/_42_/a_109_93# therm_0/_02_ therm_0/input15/a_27_47# therm_0/_43_/a_27_47#
+ therm_0/_43_/a_193_413# therm_0/_37_/a_303_47# therm_0/_55_/a_80_21# therm_0/_50_/a_515_93#
+ therm_0/input2/a_27_47# therm_0/_33_/a_109_93# therm_0/_38_/a_197_47# therm_0/input5/a_558_47#
+ therm_0/_15_ therm_0/_21_ therm_0/_50_/a_615_93# therm_0/_14_ therm_0/input12/a_27_47#
+ therm_0/_20_ therm_0/net1 therm_0/_38_/a_303_47# therm_0/_38_/a_27_47# therm_0/_40_/a_297_297#
+ therm_0/_34_/a_129_47# therm_0/_03_ therm_0/_06_ therm_0/_53_/a_29_53# therm_0/_49_/a_315_47#
+ therm_0/net16 therm_0/net10 therm_0/output18/a_27_47# therm_0/_08_ therm_0/input5/a_664_47#
+ therm_0/_16_ therm_0/_11_ therm_0/_27_/a_109_297# therm_0/_12_ therm_0/net9 therm_0/_00_
+ therm_0/_44_/a_256_47# therm_0/_05_ therm_0/_48_/a_27_47# therm_0/input6/a_27_47#
+ therm_0/net17 therm_0/_31_/a_117_297# therm_0/_50_/a_343_93# therm_0/net5 Vp Vn
+ therm_0/_29_/a_29_53# therm
Xth13_0 Vp V13 Vin th13_0/m1_831_275# Vn th13_0/m1_559_n458# th13
Xth06_0 Vp Vin V06 Vn th06_0/m1_904_n796# th06
Xth11_0 V11 Vin Vn th11_0/m1_577_n654# Vp th11_0/m1_705_187# th11
Xth04_0 Vp V04 Vn th04_0/m1_892_n998# th04_0/m1_620_n488# Vin th04
C0 V03 therm_0/input2/a_27_47# 5.03e-19
C1 V07 th08_0/m1_477_n803# 4.63e-19
C2 th01_0/m1_991_n1219# V04 2.46e-19
C3 therm_0/_02_ V06 6.08e-19
C4 therm_0/_35_/a_76_199# V07 5.17e-21
C5 V04 therm_0/_49_/a_315_47# 1.45e-20
C6 therm_0/input7/a_27_47# V04 9.09e-20
C7 therm_0/output19/a_27_47# V13 0.00421f
C8 therm_0/net2 V10 -1.73e-36
C9 V15 th10_0/m1_536_174# 0.14f
C10 V09 th12_0/m1_529_n42# 0.0422f
C11 therm_0/net19 therm_0/net14 -3.55e-33
C12 therm_0/_19_ V14 1.67e-20
C13 th01_0/m1_571_n501# V03 0.00311f
C14 th12_0/m1_529_n42# th14_0/m1_891_419# 0.0381f
C15 V14 Vin 0.00316f
C16 therm_0/net2 V12 0.00337f
C17 therm_0/input14/a_27_47# V13 1.74e-19
C18 therm_0/_48_/a_27_47# V06 3.06e-19
C19 therm_0/_19_ V02 3.37e-19
C20 V01 th04_0/m1_892_n998# 0.0457f
C21 th11_0/m1_705_187# th01_0/m1_571_n501# 9.49e-20
C22 V07 therm_0/net13 5.29e-20
C23 V03 V04 0.491f
C24 Vin V02 0.733f
C25 th15_0/Vin Vp 1.17f
C26 V13 therm_0/_37_/a_197_47# 6.97e-20
C27 V14 V02 1.37e-20
C28 b[2] therm_0/net18 3.8e-19
C29 therm_0/input8/a_27_47# Vp 1.51e-19
C30 therm_0/net14 Vp 0.00665f
C31 therm_0/_07_ V06 1.49e-19
C32 therm_0/_30_/a_215_297# V08 7.76e-20
C33 therm_0/input3/a_27_47# therm_0/net2 1.07e-32
C34 therm_0/_38_/a_197_47# b[0] 1.46e-19
C35 th13_0/m1_831_275# V15 5.89e-19
C36 therm_0/net3 V13 0.00357f
C37 therm_0/net11 b[1] 0.0013f
C38 therm_0/input6/a_27_47# V13 0.00307f
C39 b[2] therm_0/output18/a_27_47# 0.00238f
C40 therm_0/_13_ b[0] 5.29e-20
C41 V11 therm_0/net7 2.81e-20
C42 therm_0/net2 V03 8.63e-19
C43 therm_0/_27_/a_277_297# Vp 3.15e-20
C44 therm_0/_19_ Vp 0.00541f
C45 therm_0/_37_/a_109_47# V13 2.68e-21
C46 V15 th10_0/m1_502_n495# 1.36e-19
C47 Vin Vp 2.01f
C48 therm_0/input10/a_27_47# Vin 4.37e-19
C49 therm_0/net12 V08 1.17e-20
C50 therm_0/_41_/a_59_75# V13 0.00284f
C51 V14 Vp 0.107f
C52 therm_0/input11/a_27_47# Vp 6.32e-20
C53 V08 th04_0/m1_892_n998# 5.12e-19
C54 therm_0/_16_ V12 8.41e-20
C55 th11_0/m1_705_187# th02_0/m1_571_144# 1.03e-19
C56 b[1] therm_0/net17 -7.11e-33
C57 therm_0/_42_/a_109_93# V12 3.58e-19
C58 V15 th15_0/m1_597_n912# 0.00444f
C59 therm_0/_10_ V13 5.64e-19
C60 therm_0/net9 V08 7.93e-20
C61 th13_0/m1_559_n458# th15_0/Vin 0.109f
C62 b[1] V03 0.0015f
C63 Vp V02 0.298f
C64 therm_0/input15/a_27_47# V10 2.18e-20
C65 therm_0/_11_ Vp 0.00162f
C66 th11_0/m1_577_n654# V01 1.37e-21
C67 therm_0/_06_ therm_0/net18 3.55e-33
C68 V11 V12 -0.0074f
C69 V11 therm_0/_31_/a_35_297# 5.14e-20
C70 V08 therm_0/net8 1.68e-19
C71 V05 b[1] 9.42e-19
C72 therm_0/net19 Vp 6.69e-19
C73 th14_0/m1_891_419# therm_0/net5 8.26e-19
C74 therm_0/input9/a_75_212# V08 0.00104f
C75 b[3] therm_0/output19/a_27_47# 0.00611f
C76 therm_0/_14_ V13 0.00744f
C77 th15_0/m1_849_n157# th15_0/Vin 6.18e-19
C78 V11 th01_0/m1_991_n1219# 4.89e-20
C79 th12_0/m1_529_n42# th15_0/Vin 0.0262f
C80 th06_0/m1_904_n796# V08 0.00128f
C81 b[3] therm_0/input14/a_27_47# 0.00219f
C82 therm_0/_30_/a_215_297# th07_0/m1_808_n892# 4.07e-21
C83 therm_0/_17_ therm_0/_43_/a_193_413# -2.84e-32
C84 therm_0/_17_ therm_0/net15 2.84e-32
C85 th12_0/m1_529_n42# therm_0/net14 2.7e-19
C86 th13_0/m1_559_n458# Vin 0.0257f
C87 therm_0/input15/a_27_47# V15 2.79e-20
C88 therm_0/net5 therm_0/input5/a_62_47# -2.84e-32
C89 therm_0/_12_ V13 6.44e-22
C90 V04 th04_0/m1_892_n998# 0.0018f
C91 b[3] V13 0.139f
C92 therm_0/input10/a_27_47# Vp 1.73e-19
C93 V11 therm_0/net17 8.66e-20
C94 th07_0/m1_808_n892# th05_0/m1_752_n794# 1.42e-20
C95 therm_0/_30_/a_109_53# V08 2.44e-20
C96 V09 therm_0/net15 2.01e-19
C97 therm_0/output19/a_27_47# th10_0/m1_536_174# 5.9e-19
C98 V11 V03 2.67e-20
C99 therm_0/_40_/a_297_297# Vp 2.01e-20
C100 therm_0/net7 therm_0/input5/a_664_47# 2.22e-34
C101 th07_0/m1_808_n892# th04_0/m1_892_n998# 1.1e-19
C102 therm_0/_17_ V12 0.00532f
C103 therm_0/_43_/a_27_47# V13 8.99e-20
C104 therm_0/_07_ Vin 1.97e-19
C105 th15_0/m1_849_n157# Vin 0.00238f
C106 V04 therm_0/net8 0.0042f
C107 therm_0/input14/a_27_47# th10_0/m1_536_174# 1.05e-19
C108 th12_0/m1_529_n42# Vin 0.0104f
C109 th03_0/m1_638_n591# th15_0/Vin 3.89e-19
C110 th11_0/m1_705_187# V11 0.00226f
C111 th12_0/m1_529_n42# V14 1.86e-19
C112 therm_0/_31_/a_285_297# V04 2.68e-20
C113 th14_0/m1_641_n318# th11_0/m1_705_187# 5.69e-22
C114 V09 V10 0.0058f
C115 therm_0/_27_/a_27_297# V03 2.64e-19
C116 V13 th10_0/m1_536_174# 7.91e-19
C117 therm_0/_02_ Vp 1.91e-20
C118 V09 V12 0.0147f
C119 therm_0/_43_/a_469_47# V13 2.86e-20
C120 Vin th08_0/m1_477_n803# 0.0549f
C121 therm_0/output17/a_27_47# V03 6.3e-20
C122 V12 th14_0/m1_891_419# 2.97e-19
C123 b[1] th05_0/m1_752_n794# 0.00134f
C124 therm_0/input1/a_75_212# V03 9.16e-20
C125 therm_0/_44_/a_93_21# Vp 2.04e-20
C126 therm_0/input12/a_27_47# th05_0/m1_752_n794# 1.02e-20
C127 V07 therm_0/_33_/a_109_93# 2.32e-20
C128 th12_0/m1_529_n42# therm_0/net19 8.54e-21
C129 therm_0/net12 b[1] 2.56e-19
C130 th13_0/m1_559_n458# Vp 0.00128f
C131 V11 therm_0/_31_/a_117_297# 6.45e-20
C132 th07_0/m1_808_n892# th06_0/m1_904_n796# 2e-19
C133 b[1] th04_0/m1_892_n998# 4.96e-20
C134 therm_0/_33_/a_209_311# V07 5.46e-19
C135 th01_0/m1_991_n1219# th14_0/m1_891_419# 0.0018f
C136 Vin therm_0/net13 0.00225f
C137 V07 V05 -0.00237f
C138 V09 V15 0.0108f
C139 V01 V04 1.87e-19
C140 b[3] therm_0/_44_/a_250_297# 2.47e-20
C141 therm_0/net2 V13 0.00676f
C142 therm_0/_20_ V13 2.02e-20
C143 therm_0/output19/a_27_47# th10_0/m1_502_n495# 5.96e-21
C144 therm_0/net7 therm_0/input5/a_558_47# -4.44e-34
C145 th15_0/Vin therm_0/net5 1.17e-19
C146 therm_0/_40_/a_191_297# Vp 3.24e-20
C147 therm_0/_30_/a_109_53# th07_0/m1_808_n892# 2.97e-19
C148 th13_0/m1_831_275# V13 0.025f
C149 th15_0/m1_849_n157# Vp 0.0962f
C150 th12_0/m1_529_n42# Vp 0.0728f
C151 th03_0/m1_638_n591# V02 0.155f
C152 th15_0/Vin th02_0/m1_983_133# 0.0246f
C153 therm_0/net11 V06 0.004f
C154 therm_0/_30_/a_297_297# V08 2.34e-20
C155 therm_0/_04_ V04 7.55e-21
C156 therm_0/_37_/a_303_47# V13 4.34e-20
C157 therm_0/net3 therm_0/net2 5.68e-32
C158 b[1] th06_0/m1_904_n796# 4.51e-22
C159 th09_0/m1_485_n505# th02_0/m1_571_144# 0.00503f
C160 Vp th08_0/m1_477_n803# 0.0288f
C161 th11_0/m1_577_n654# th02_0/m1_571_144# 0.0183f
C162 th11_0/m1_705_187# th14_0/m1_891_419# 0.00195f
C163 V13 th15_0/m1_597_n912# 1.75e-19
C164 th09_0/m1_485_n505# th13_0/m1_831_275# 2.23e-19
C165 therm_0/_40_/a_109_297# V13 5.51e-19
C166 th03_0/m1_890_n844# th15_0/Vin 0.00307f
C167 therm_0/net5 V14 5.97e-19
C168 V04 V08 0.367f
C169 th12_0/m1_529_n42# therm_0/_15_ 6.89e-21
C170 therm_0/_10_ b[0] 6.36e-19
C171 th02_0/m1_983_133# Vin 0.0306f
C172 th03_0/m1_638_n591# Vp 0.015f
C173 b[1] V01 -2.22e-34
C174 therm_0/net1 V04 7.07e-19
C175 V07 therm_0/_30_/a_215_297# 3.38e-20
C176 therm_0/_16_ V13 1.59e-19
C177 th12_0/m1_529_n42# therm_0/_44_/a_93_21# 3.52e-20
C178 V05 V06 0.0335f
C179 b[3] th10_0/m1_536_174# 0.0209f
C180 V11 therm_0/net8 0.00138f
C181 therm_0/_48_/a_181_47# V06 8.04e-20
C182 th13_0/m1_559_n458# th12_0/m1_529_n42# 9.14e-21
C183 th07_0/m1_808_n892# V08 0.0144f
C184 th04_0/m1_620_n488# th15_0/Vin 4.08e-20
C185 therm_0/output17/a_27_47# th04_0/m1_892_n998# 6.65e-21
C186 V12 th15_0/Vin 1.05e-21
C187 th02_0/m1_983_133# V02 0.148f
C188 V07 th05_0/m1_752_n794# 8.88e-20
C189 therm_0/input1/a_75_212# th04_0/m1_892_n998# 8.62e-20
C190 therm_0/net7 Vin 0.00253f
C191 V12 therm_0/net14 5.86e-19
C192 therm_0/_49_/a_75_199# V04 1.31e-19
C193 therm_0/input15/a_27_47# V13 0.00627f
C194 V07 therm_0/net12 0.00579f
C195 therm_0/_34_/a_47_47# b[1] 2.87e-19
C196 th01_0/m1_991_n1219# th15_0/Vin -0.0283f
C197 therm_0/_20_ V08 1.54e-20
C198 therm_0/net15 V14 3.51e-20
C199 th03_0/m1_890_n844# Vin 4.79e-20
C200 V07 therm_0/net9 9.98e-20
C201 th13_0/m1_831_275# th12_0/m1_394_n856# 4.06e-20
C202 b[3] therm_0/net2 3.67e-19
C203 therm_0/_12_ b[0] 7.1e-19
C204 th15_0/Vin V15 0.113f
C205 therm_0/_06_ therm_0/_52_/a_93_21# 1.42e-32
C206 V10 Vin 0.00422f
C207 therm_0/_37_/a_27_47# V13 0.00122f
C208 th03_0/m1_890_n844# V02 0.0161f
C209 V07 therm_0/_35_/a_556_47# 3.98e-20
C210 b[1] V08 6.98e-19
C211 V11 th11_0/m1_577_n654# 1.77e-19
C212 th04_0/m1_620_n488# Vin 0.00123f
C213 th14_0/m1_641_n318# th09_0/m1_485_n505# 6.8e-20
C214 V12 Vin 4.48e-19
C215 b[1] therm_0/net1 -1.78e-33
C216 V11 V01 0.0332f
C217 therm_0/_31_/a_35_297# Vin 3.63e-19
C218 th02_0/m1_983_133# Vp 0.043f
C219 therm_0/input9/a_75_212# V07 8.08e-20
C220 V12 V14 0.00395f
C221 th15_0/Vin V03 0.161f
C222 th07_0/m1_808_n892# V04 2.45e-19
C223 V07 th06_0/m1_904_n796# 0.0101f
C224 therm_0/net11 Vin 4.33e-19
C225 th01_0/m1_991_n1219# Vin 0.0145f
C226 V03 therm_0/net14 8.33e-20
C227 therm_0/net10 V08 9.08e-20
C228 V07 therm_0/_08_ 0.00247f
C229 th11_0/m1_705_187# th15_0/Vin 0.0188f
C230 V10 therm_0/net19 0.00129f
C231 therm_0/_17_ V13 0.00307f
C232 therm_0/net2 th10_0/m1_536_174# 0.00224f
C233 therm_0/input7/a_27_47# Vin 0.00446f
C234 th05_0/m1_752_n794# V06 0.00786f
C235 therm_0/net7 Vp 4.07e-20
C236 therm_0/net6 V10 0.00123f
C237 therm_0/_20_ V04 2.62e-20
C238 therm_0/output17/a_27_47# V01 -3.55e-33
C239 V12 therm_0/net19 1.7e-19
C240 V15 Vin 0.0975f
C241 therm_0/net15 Vp 0.00272f
C242 V09 therm_0/input14/a_27_47# 7.36e-19
C243 th01_0/m1_991_n1219# V02 0.276f
C244 V07 therm_0/_30_/a_109_53# 3.03e-21
C245 therm_0/net12 V06 0.00548f
C246 therm_0/_42_/a_368_53# th12_0/m1_529_n42# 1.6e-20
C247 th03_0/m1_890_n844# Vp 0.0291f
C248 b[2] therm_0/_25_ 1.25e-19
C249 therm_0/_33_/a_109_93# Vin 1.17e-19
C250 V09 therm_0/_37_/a_197_47# 1.24e-19
C251 V09 V13 0.0209f
C252 therm_0/_19_ V03 5.68e-20
C253 therm_0/_33_/a_209_311# Vin 2.12e-19
C254 therm_0/_50_/a_343_93# V13 1.61e-20
C255 V03 Vin 0.289f
C256 V08 therm_0/_05_ 7.85e-21
C257 therm_0/_55_/a_80_21# V12 4.04e-20
C258 b[1] V04 0.00206f
C259 V10 Vp 0.065f
C260 V11 therm_0/net1 2.77e-20
C261 th04_0/m1_620_n488# Vp 0.00246f
C262 th14_0/m1_641_n318# th12_0/m1_394_n856# 0.00861f
C263 V12 Vp 0.121f
C264 V05 Vin 0.0101f
C265 th11_0/m1_705_187# Vin 0.278f
C266 V15 therm_0/net19 2.85e-20
C267 therm_0/_31_/a_35_297# Vp 2.44e-20
C268 V03 V02 0.687f
C269 therm_0/net6 V15 2.17e-20
C270 therm_0/net3 V09 3.48e-19
C271 th07_0/m1_808_n892# b[1] 7.76e-22
C272 V09 th09_0/m1_485_n505# 0.0285f
C273 therm_0/net3 th14_0/m1_891_419# 2.85e-21
C274 V07 therm_0/_04_ 1.09e-20
C275 th06_0/m1_904_n796# therm_0/input13/a_27_47# 5.34e-20
C276 V11 therm_0/input2/a_27_47# 2.03e-19
C277 th09_0/m1_485_n505# th14_0/m1_891_419# 3.27e-19
C278 therm_0/_34_/a_47_47# V07 1.77e-20
C279 th01_0/m1_991_n1219# Vp 0.0217f
C280 therm_0/net11 Vp 1.27e-20
C281 th06_0/m1_904_n796# V06 0.00888f
C282 th11_0/m1_705_187# V02 0.0253f
C283 V09 therm_0/_37_/a_109_47# 2.42e-20
C284 therm_0/input7/a_27_47# Vp 3.83e-20
C285 therm_0/net2 b[1] 3.55e-33
C286 th07_0/m1_808_n892# therm_0/net10 6.94e-21
C287 V15 Vp 0.0545f
C288 therm_0/_31_/a_117_297# Vin 2.46e-19
C289 V10 therm_0/_15_ 3.47e-36
C290 therm_0/_17_ therm_0/_44_/a_250_297# -1.42e-32
C291 V07 V08 0.376f
C292 Vp therm_0/net17 7.29e-19
C293 V12 therm_0/_15_ 0.00395f
C294 therm_0/_14_ therm_0/_17_ -1.14e-31
C295 therm_0/net14 therm_0/_42_/a_209_311# 2.84e-32
C296 V04 therm_0/_05_ 3.87e-20
C297 th15_0/Vin th04_0/m1_892_n998# 5.5e-20
C298 V11 V04 2.17e-20
C299 V03 Vp 0.401f
C300 therm_0/_44_/a_93_21# V12 4.59e-19
C301 therm_0/_42_/a_296_53# therm_0/net14 -5.55e-35
C302 therm_0/_02_ therm_0/net11 1.42e-32
C303 th12_0/m1_529_n42# therm_0/net15 2.75e-20
C304 V05 Vp 0.0176f
C305 th11_0/m1_705_187# Vp 0.0228f
C306 therm_0/_30_/a_215_297# Vin 9.95e-20
C307 b[1] therm_0/net10 4.52e-19
C308 V09 th12_0/m1_394_n856# 0.00496f
C309 therm_0/_37_/a_27_47# th10_0/m1_536_174# 3.2e-20
C310 th03_0/m1_638_n591# th02_0/m1_983_133# 3.07e-20
C311 therm_0/input5/a_381_47# th14_0/m1_891_419# 9.97e-21
C312 th14_0/m1_891_419# th12_0/m1_394_n856# 5.71e-20
C313 therm_0/output17/a_27_47# V04 1.07e-19
C314 th12_0/m1_529_n42# V10 2.39e-20
C315 th05_0/m1_752_n794# Vin 0.00961f
C316 therm_0/_34_/a_47_47# V06 0.00112f
C317 th09_0/m1_962_372# th02_0/m1_571_144# 0.0112f
C318 therm_0/input1/a_75_212# V04 5.43e-20
C319 V11 th02_0/m1_571_144# 4.75e-20
C320 V11 therm_0/net2 7.31e-20
C321 therm_0/input11/a_27_47# th05_0/m1_752_n794# 7.08e-19
C322 V09 b[3] 8.61e-19
C323 th12_0/m1_529_n42# V12 7.31e-19
C324 therm_0/input14/a_27_47# therm_0/net14 -1.42e-32
C325 therm_0/net12 Vin 0.00114f
C326 th15_0/Vin V13 0.0177f
C327 therm_0/_34_/a_129_47# b[1] 6.11e-20
C328 Vin th04_0/m1_892_n998# 0.111f
C329 th14_0/m1_891_419# therm_0/input2/a_27_47# 1.62e-21
C330 therm_0/_06_ V13 0.00596f
C331 V07 V04 2.58e-19
C332 therm_0/_06_ th06_0/m1_904_n796# 6.48e-20
C333 V07 therm_0/_09_ 8.07e-21
C334 therm_0/_00_ V13 9.74e-20
C335 therm_0/net14 V13 0.00243f
C336 therm_0/net9 Vin 2.85e-19
C337 th04_0/m1_620_n488# th08_0/m1_477_n803# 6.18e-20
C338 V06 V08 2.48e-21
C339 therm_0/_02_ therm_0/_48_/a_181_47# -5.55e-35
C340 V11 b[1] 0.00899f
C341 therm_0/output19/a_27_47# Vin 5.09e-21
C342 V02 th04_0/m1_892_n998# 2.47e-19
C343 V07 th07_0/m1_808_n892# 0.00985f
C344 th09_0/m1_485_n505# th15_0/Vin 0.113f
C345 th15_0/m1_849_n157# V15 0.0377f
C346 Vin therm_0/net8 0.00281f
C347 th12_0/m1_529_n42# V15 6.17e-20
C348 th11_0/m1_577_n654# th15_0/Vin 0.0157f
C349 therm_0/input14/a_27_47# Vin 1.03e-20
C350 V09 th10_0/m1_536_174# 0.0109f
C351 th15_0/Vin V01 0.00134f
C352 therm_0/_31_/a_285_297# Vin 1.62e-19
C353 therm_0/input9/a_75_212# Vin 8.54e-19
C354 therm_0/input3/a_27_47# th12_0/m1_529_n42# 5.38e-19
C355 therm_0/input7/a_27_47# th08_0/m1_477_n803# 4.89e-21
C356 Vin V13 0.0223f
C357 th06_0/m1_904_n796# Vin 0.0329f
C358 therm_0/_03_ V08 1.64e-19
C359 therm_0/_08_ Vin 2.42e-19
C360 therm_0/output17/a_27_47# b[1] 2.84e-32
C361 th05_0/m1_752_n794# Vp 0.00105f
C362 therm_0/_17_ therm_0/net2 -5.68e-32
C363 therm_0/_48_/a_109_47# V06 4.35e-21
C364 therm_0/input1/a_75_212# b[1] 8.88e-34
C365 th05_0/m1_752_n794# therm_0/input10/a_27_47# 5.27e-20
C366 therm_0/_42_/a_368_53# V12 7.6e-21
C367 therm_0/net12 Vp 1.27e-20
C368 therm_0/_11_ V13 0.00386f
C369 V03 th08_0/m1_477_n803# 2.7e-19
C370 Vp th04_0/m1_892_n998# 0.0342f
C371 therm_0/_30_/a_109_53# Vin 3.24e-20
C372 V07 b[1] 0.00129f
C373 th09_0/m1_485_n505# Vin 0.0284f
C374 V09 therm_0/net2 2.68e-19
C375 V09 th02_0/m1_571_144# 3.21e-19
C376 th11_0/m1_577_n654# Vin 0.0113f
C377 therm_0/net19 V13 0.00504f
C378 therm_0/_47_/a_81_21# V13 4.03e-19
C379 therm_0/net2 th14_0/m1_891_419# 0.00232f
C380 V01 Vin 0.105f
C381 therm_0/net6 V13 0.00332f
C382 V09 th13_0/m1_831_275# 0.0162f
C383 therm_0/_50_/a_515_93# V13 3.52e-23
C384 th03_0/m1_890_n844# th02_0/m1_983_133# 0.00116f
C385 therm_0/output19/a_27_47# Vp 5.68e-32
C386 V07 therm_0/net10 8.76e-20
C387 therm_0/input5/a_381_47# th15_0/Vin 1.42e-20
C388 Vp therm_0/net8 7.31e-20
C389 th12_0/m1_394_n856# th15_0/Vin 0.0129f
C390 th07_0/m1_808_n892# V06 1.26e-19
C391 th11_0/m1_577_n654# V02 3.43e-19
C392 th03_0/m1_638_n591# V03 2.96e-19
C393 therm_0/_34_/a_285_47# b[1] 1.52e-19
C394 therm_0/input14/a_27_47# Vp 0.00279f
C395 V01 V02 0.193f
C396 V09 therm_0/_37_/a_303_47# 7.76e-20
C397 therm_0/input9/a_75_212# Vp 1.45e-19
C398 V09 th10_0/m1_502_n495# 0.00223f
C399 therm_0/input8/a_27_47# V08 9.25e-20
C400 therm_0/_06_ therm_0/_53_/a_29_53# -1.42e-32
C401 therm_0/_04_ Vin 3.49e-19
C402 therm_0/_03_ V04 3.61e-20
C403 Vp V13 0.176f
C404 therm_0/_34_/a_47_47# Vin 1.73e-19
C405 th06_0/m1_904_n796# Vp 0.0244f
C406 therm_0/_04_ V14 1.51e-20
C407 therm_0/output17/a_27_47# V11 9.4e-19
C408 therm_0/input1/a_75_212# V11 1.21e-19
C409 b[3] therm_0/net14 8.66e-19
C410 therm_0/_04_ V02 3.66e-19
C411 V07 therm_0/_05_ 2.71e-21
C412 therm_0/_40_/a_297_297# V13 1.13e-19
C413 b[2] b[0] 0.00937f
C414 therm_0/net15 V10 1.24e-20
C415 th15_0/Vin th01_0/m1_571_n501# -5.68e-32
C416 therm_0/net3 Vp 0.00564f
C417 Vin V08 0.341f
C418 th09_0/m1_485_n505# Vp 0.0355f
C419 b[1] V06 0.00158f
C420 th12_0/m1_394_n856# Vin 0.0013f
C421 V12 therm_0/_43_/a_193_413# 4.53e-20
C422 therm_0/net15 V12 1.71e-19
C423 th11_0/m1_577_n654# Vp 0.0262f
C424 therm_0/net1 Vin 0.00253f
C425 th12_0/m1_529_n42# therm_0/_42_/a_209_311# 5.57e-20
C426 therm_0/net4 b[0] 1.19e-19
C427 therm_0/input12/a_27_47# V06 0.00449f
C428 therm_0/_01_ Vp 1.37e-19
C429 V01 Vp 0.124f
C430 th15_0/Vin th10_0/m1_536_174# 3.79e-20
C431 therm_0/_15_ V13 0.00684f
C432 b[3] Vin 2.69e-21
C433 therm_0/_42_/a_296_53# th12_0/m1_529_n42# 6.15e-21
C434 b[2] b[1] 0.014f
C435 Vin therm_0/input2/a_27_47# 4.93e-19
C436 V09 th09_0/m1_962_372# 8.77e-19
C437 therm_0/net14 th10_0/m1_536_174# 8.25e-20
C438 therm_0/net10 V06 0.00893f
C439 therm_0/_06_ therm_0/_09_ 1.42e-32
C440 th02_0/m1_983_133# V03 2.47e-20
C441 therm_0/net1 V02 0.00409f
C442 therm_0/input8/a_27_47# V04 0.00453f
C443 V12 V10 -0.00566f
C444 therm_0/_44_/a_93_21# V13 9.89e-20
C445 V11 th14_0/m1_891_419# 0.0727f
C446 th14_0/m1_641_n318# V09 0.00306f
C447 therm_0/_04_ Vp 0.00522f
C448 therm_0/net15 V15 1.44e-20
C449 th08_0/m1_477_n803# th04_0/m1_892_n998# 0.00506f
C450 th01_0/m1_571_n501# Vin 6.06e-19
C451 therm_0/_50_/a_615_93# V13 6.88e-20
C452 th07_0/m1_808_n892# therm_0/input8/a_27_47# 7.82e-20
C453 therm_0/_34_/a_129_47# V06 3.25e-20
C454 therm_0/net7 V03 0.0134f
C455 therm_0/_27_/a_27_297# th14_0/m1_891_419# 7.3e-21
C456 therm_0/net2 th15_0/Vin 5.84e-20
C457 th01_0/m1_991_n1219# th04_0/m1_620_n488# 7.52e-20
C458 th15_0/Vin th02_0/m1_571_144# 0.00185f
C459 V09 therm_0/_37_/a_27_47# 3.2e-19
C460 Vin th10_0/m1_536_174# 0.0136f
C461 therm_0/_40_/a_191_297# V13 2.53e-19
C462 th13_0/m1_831_275# th15_0/Vin 0.0168f
C463 V04 Vin 0.266f
C464 V15 V10 0.026f
C465 th01_0/m1_571_n501# V02 1.29e-19
C466 th13_0/m1_559_n458# th09_0/m1_485_n505# 0.00612f
C467 therm_0/output17/a_27_47# th14_0/m1_891_419# 3.28e-21
C468 therm_0/_06_ b[0] 3.27e-19
C469 th15_0/m1_849_n157# V13 0.0405f
C470 th03_0/m1_890_n844# V03 0.0141f
C471 therm_0/net2 therm_0/net14 -1.42e-32
C472 Vp V08 0.0542f
C473 therm_0/_18_ V12 9.22e-20
C474 th12_0/m1_394_n856# Vp 0.0157f
C475 therm_0/input3/a_27_47# V12 0.00164f
C476 V04 V02 3.64e-19
C477 th07_0/m1_808_n892# Vin 0.0319f
C478 b[3] Vp 0.00542f
C479 th06_0/m1_904_n796# th08_0/m1_477_n803# 2.84e-21
C480 therm_0/_06_ b[1] 7.29e-20
C481 Vp therm_0/input2/a_27_47# 5.42e-20
C482 therm_0/_17_ V09 8.68e-20
C483 th15_0/Vin th15_0/m1_597_n912# 0.0049f
C484 th04_0/m1_620_n488# V03 0.00358f
C485 therm_0/net19 th10_0/m1_536_174# 0.00606f
C486 therm_0/net3 th12_0/m1_529_n42# 0.00151f
C487 therm_0/_29_/a_29_53# V08 1.72e-20
C488 therm_0/net2 Vin 5.78e-19
C489 th02_0/m1_571_144# Vin 0.00869f
C490 therm_0/_49_/a_75_199# Vp 5.91e-20
C491 therm_0/net2 V14 0.0168f
C492 th01_0/m1_991_n1219# V03 0.0279f
C493 V07 therm_0/input13/a_27_47# 2.09e-19
C494 th13_0/m1_831_275# Vin 0.0149f
C495 therm_0/output16/a_27_47# b[0] 7.49e-20
C496 th01_0/m1_571_n501# Vp 0.0265f
C497 therm_0/_02_ V08 7.56e-21
C498 therm_0/_06_ therm_0/_23_ -2.84e-32
C499 V09 th14_0/m1_891_419# 0.00256f
C500 V07 V06 0.19f
C501 V03 therm_0/input7/a_27_47# 0.00466f
C502 th02_0/m1_571_144# V02 2.06e-20
C503 th06_0/m1_904_n796# therm_0/net13 1.1e-20
C504 therm_0/net2 V02 0.00263f
C505 V01 th08_0/m1_477_n803# 7.8e-21
C506 th11_0/m1_705_187# th01_0/m1_991_n1219# 0.00182f
C507 Vp th10_0/m1_536_174# 0.0704f
C508 therm_0/_11_ b[0] 4.2e-19
C509 b[1] Vin 0.121f
C510 Vin th10_0/m1_502_n495# 1.09e-19
C511 V04 Vp 0.066f
C512 th13_0/m1_559_n458# th12_0/m1_394_n856# 3.47e-20
C513 therm_0/input12/a_27_47# Vin 8.31e-19
C514 V03 therm_0/net17 4.77e-20
C515 Vin th15_0/m1_597_n912# 3.87e-19
C516 therm_0/_44_/a_346_47# V13 1.36e-20
C517 th09_0/m1_962_372# th15_0/Vin 0.0637f
C518 V11 th15_0/Vin 7.42e-19
C519 th14_0/m1_891_419# therm_0/input5/a_62_47# 5.09e-20
C520 b[1] V02 0.00575f
C521 therm_0/_34_/a_285_47# V06 2.04e-19
C522 th12_0/m1_529_n42# therm_0/_44_/a_250_297# 5.4e-20
C523 therm_0/_38_/a_109_47# b[0] 1.12e-19
C524 th07_0/m1_808_n892# Vp 0.0215f
C525 therm_0/net10 Vin 4.22e-19
C526 th14_0/m1_641_n318# th15_0/Vin 0.0354f
C527 therm_0/_14_ th12_0/m1_529_n42# 5.6e-21
C528 th11_0/m1_705_187# V03 1.97e-21
C529 th12_0/m1_529_n42# th12_0/m1_394_n856# 1.78e-33
C530 th02_0/m1_571_144# Vp 0.026f
C531 therm_0/net2 Vp 0.0284f
C532 Vp b[0] 4.51e-19
C533 therm_0/net5 V13 6.23e-19
C534 therm_0/_02_ V04 8.59e-21
C535 th13_0/m1_831_275# Vp 0.0388f
C536 V10 therm_0/_42_/a_209_311# -8.67e-37
C537 th08_0/m1_477_n803# V08 0.0132f
C538 Vin therm_0/_05_ 3.91e-21
C539 th09_0/m1_962_372# Vin 6.36e-19
C540 therm_0/input5/a_841_47# therm_0/net7 2.22e-34
C541 V12 therm_0/_42_/a_209_311# 2.21e-19
C542 V11 Vin 0.0701f
C543 b[1] Vp 0.00519f
C544 Vp th10_0/m1_502_n495# 0.0351f
C545 V11 V14 0.00945f
C546 th14_0/m1_641_n318# Vin 0.0621f
C547 therm_0/input12/a_27_47# Vp 9.21e-20
C548 therm_0/_42_/a_296_53# V12 6.58e-21
C549 th14_0/m1_641_n318# V14 6.65e-19
C550 V07 therm_0/_06_ 1.47e-19
C551 Vp th15_0/m1_597_n912# -7.11e-33
C552 therm_0/_40_/a_109_297# Vp 2.19e-21
C553 therm_0/net11 th05_0/m1_752_n794# 3.2e-20
C554 therm_0/_44_/a_256_47# V13 1.36e-20
C555 V11 V02 0.00259f
C556 th09_0/m1_485_n505# th02_0/m1_983_133# 0.00736f
C557 V10 therm_0/output19/a_27_47# 8.86e-19
C558 therm_0/_43_/a_193_413# V13 3.38e-19
C559 therm_0/net15 V13 0.0112f
C560 th11_0/m1_577_n654# th02_0/m1_983_133# 1.64e-19
C561 th12_0/m1_529_n42# th10_0/m1_536_174# 0.002f
C562 th01_0/m1_991_n1219# th04_0/m1_892_n998# 0.00552f
C563 therm_0/output17/a_27_47# Vin 8.69e-20
C564 therm_0/_44_/a_93_21# therm_0/net2 -1.42e-32
C565 V09 th15_0/Vin 0.201f
C566 therm_0/input1/a_75_212# Vin 6.51e-19
C567 th14_0/m1_891_419# th15_0/Vin 0.00394f
C568 V10 V13 0.00381f
C569 V09 therm_0/net14 8.76e-19
C570 V07 Vin 0.259f
C571 therm_0/output17/a_27_47# V02 0.00158f
C572 th14_0/m1_891_419# therm_0/net14 2.05e-22
C573 V04 th08_0/m1_477_n803# 0.00364f
C574 therm_0/input12/a_27_47# therm_0/_02_ -2.78e-35
C575 therm_0/_47_/a_384_47# V13 1.59e-20
C576 therm_0/input1/a_75_212# V02 0.00364f
C577 th09_0/m1_962_372# Vp 0.0369f
C578 V15 therm_0/output19/a_27_47# 2.68e-19
C579 V03 th04_0/m1_892_n998# 0.0479f
C580 V05 th05_0/m1_752_n794# 0.00814f
C581 th15_0/Vin therm_0/input5/a_62_47# 1.58e-19
C582 V11 Vp 0.179f
C583 therm_0/_02_ therm_0/net10 1.11e-34
C584 th07_0/m1_808_n892# th08_0/m1_477_n803# 4.41e-19
C585 th12_0/m1_529_n42# therm_0/net2 0.00934f
C586 th14_0/m1_641_n318# Vp 0.0569f
C587 therm_0/net3 V10 -1.39e-35
C588 th15_0/m1_849_n157# th13_0/m1_831_275# 0.0859f
C589 therm_0/_55_/a_217_297# V12 1.58e-20
C590 th12_0/m1_529_n42# th13_0/m1_831_275# 1.36e-20
C591 V10 therm_0/input6/a_27_47# 1.24e-19
C592 therm_0/_06_ V06 0.00345f
C593 therm_0/_19_ th14_0/m1_891_419# 1.7e-20
C594 therm_0/net3 V12 0.00439f
C595 V09 Vin 0.303f
C596 th14_0/m1_891_419# Vin 0.0341f
C597 V09 V14 0.0137f
C598 therm_0/_18_ V13 7.47e-20
C599 therm_0/_27_/a_27_297# Vp 5.79e-19
C600 th14_0/m1_891_419# V14 0.0958f
C601 therm_0/_38_/a_303_47# b[0] 1.51e-19
C602 V15 V13 2.37f
C603 V03 therm_0/net8 5.72e-21
C604 th04_0/m1_620_n488# V01 0.00118f
C605 therm_0/_37_/a_27_47# Vp 3.98e-19
C606 th12_0/m1_529_n42# th10_0/m1_502_n495# 8.5e-20
C607 therm_0/_21_ V08 4.8e-21
C608 therm_0/output17/a_27_47# Vp 7.75e-19
C609 therm_0/_06_ b[2] 1.78e-33
C610 therm_0/input1/a_75_212# Vp 2.57e-19
C611 therm_0/_11_ V09 3.33e-20
C612 th14_0/m1_891_419# V02 2.17e-19
C613 th01_0/m1_991_n1219# V01 0.0641f
C614 therm_0/net16 b[0] 7.31e-19
C615 therm_0/input13/a_27_47# Vin 0.00344f
C616 therm_0/input5/a_381_47# therm_0/net7 1.11e-34
C617 V12 therm_0/_10_ 6.2e-21
C618 V07 Vp 0.0734f
C619 V09 therm_0/net19 5.64e-20
C620 therm_0/input5/a_62_47# V14 0.00147f
C621 therm_0/_06_ therm_0/_24_ -2.84e-32
C622 V06 Vin 0.264f
C623 V15 therm_0/input6/a_27_47# 4.39e-20
C624 therm_0/_43_/a_369_47# V13 8.56e-20
C625 V05 th06_0/m1_904_n796# 3.54e-20
C626 therm_0/_17_ Vp 1.66e-20
C627 V12 therm_0/_44_/a_250_297# 0.001f
C628 therm_0/_14_ V10 8.67e-37
C629 therm_0/_42_/a_109_93# th12_0/m1_529_n42# 8.33e-20
C630 therm_0/_01_ V03 4.31e-20
C631 therm_0/_14_ V12 9.3e-20
C632 V03 V01 0.102f
C633 V09 Vp 0.849f
C634 th04_0/m1_620_n488# V08 3.51e-21
C635 th14_0/m1_891_419# Vp 0.0168f
C636 V12 th12_0/m1_394_n856# 3.8e-19
C637 therm_0/_31_/a_35_297# V08 1.47e-20
C638 therm_0/_03_ Vin 2.54e-19
C639 therm_0/_47_/a_299_297# V13 1.28e-19
C640 therm_0/_21_ V04 2.85e-20
C641 V11 th12_0/m1_529_n42# 9.69e-21
C642 b[3] V10 0.00495f
C643 th11_0/m1_705_187# V01 0.00427f
C644 Vp therm_0/input5/a_664_47# -2.84e-32
C645 therm_0/net12 th05_0/m1_752_n794# 2.87e-20
C646 therm_0/_38_/a_27_47# b[0] 5.6e-19
C647 th03_0/m1_890_n844# th01_0/m1_571_n501# 0.00797f
C648 therm_0/net11 V08 3.73e-20
C649 V03 therm_0/_04_ 1.22e-20
C650 therm_0/_17_ therm_0/_15_ -1.42e-32
C651 therm_0/net7 V04 2.13e-21
C652 therm_0/input13/a_27_47# Vp 1.48e-19
C653 therm_0/_44_/a_584_47# Vp 2.94e-20
C654 therm_0/_27_/a_205_297# Vp 3.97e-20
C655 therm_0/_17_ therm_0/_44_/a_93_21# 2.84e-32
C656 V06 Vp 0.0537f
C657 V06 therm_0/input10/a_27_47# 3.7e-19
C658 therm_0/_34_/a_285_47# therm_0/_02_ -1.11e-34
C659 therm_0/_27_/a_109_297# Vp 7.33e-20
C660 th15_0/Vin Vin 0.825f
C661 V10 th10_0/m1_536_174# 0.0101f
C662 th15_0/Vin V14 0.0121f
C663 b[3] V15 0.0365f
C664 V03 V08 -0.00105f
C665 therm_0/_06_ Vin 7.03e-19
C666 b[2] Vp 0.00709f
C667 V07 therm_0/_07_ 0.00369f
C668 V12 th10_0/m1_536_174# 9.23e-19
C669 th05_0/m1_752_n794# th06_0/m1_904_n796# 0.00251f
C670 therm_0/input8/a_27_47# Vin 0.00341f
C671 th13_0/m1_559_n458# V09 0.0377f
C672 therm_0/net14 Vin 6.33e-21
C673 V03 therm_0/net1 4.1e-19
C674 therm_0/_31_/a_35_297# V04 5.41e-20
C675 th15_0/Vin V02 0.652f
C676 therm_0/net12 th06_0/m1_904_n796# 2.92e-22
C677 therm_0/_17_ th12_0/m1_529_n42# 2.42e-20
C678 th11_0/m1_705_187# th12_0/m1_394_n856# 6.45e-22
C679 V04 Vn 0.773f
C680 th04_0/m1_892_n998# Vn 0.834f
C681 th04_0/m1_620_n488# Vn 0.0632f
C682 th11_0/m1_705_187# Vn 0.549f
C683 V11 Vn 0.86f
C684 Vin Vn 16.1f
C685 th11_0/m1_577_n654# Vn 0.322f
C686 th06_0/m1_904_n796# Vn 0.502f
C687 V06 Vn 0.777f
C688 th13_0/m1_831_275# Vn 1.08f
C689 V13 Vn 2.84f
C690 th13_0/m1_559_n458# Vn 0.303f
C691 therm_0/_04_ Vn 0.337f
C692 therm_0/net9 Vn 0.357f
C693 therm_0/_03_ Vn 0.36f
C694 therm_0/net10 Vn 0.422f
C695 therm_0/_30_/a_109_53# Vn 0.159f
C696 therm_0/_30_/a_215_297# Vn 0.142f
C697 therm_0/_05_ Vn 0.152f
C698 therm_0/net8 Vn 0.389f
C699 therm_0/_31_/a_285_297# Vn 0.00137f
C700 therm_0/_31_/a_35_297# Vn 0.255f
C701 therm_0/_32_/a_27_47# Vn 0.175f
C702 therm_0/_11_ Vn 0.267f
C703 therm_0/_50_/a_343_93# Vn 0.172f
C704 therm_0/_50_/a_223_47# Vn 0.141f
C705 therm_0/_50_/a_27_47# Vn 0.259f
C706 therm_0/_07_ Vn 0.288f
C707 therm_0/_06_ Vn 0.789f
C708 therm_0/_33_/a_209_311# Vn 0.143f
C709 therm_0/_33_/a_109_93# Vn 0.158f
C710 therm_0/_08_ Vn 0.131f
C711 therm_0/net11 Vn 0.771f
C712 therm_0/_34_/a_285_47# Vn 0.0174f
C713 therm_0/_34_/a_47_47# Vn 0.199f
C714 therm_0/_23_ Vn 0.106f
C715 therm_0/input15/a_27_47# Vn 0.208f
C716 therm_0/_09_ Vn 0.142f
C717 therm_0/_35_/a_489_413# Vn 0.0254f
C718 therm_0/_35_/a_226_47# Vn 0.162f
C719 therm_0/_35_/a_76_199# Vn 0.141f
C720 therm_0/_24_ Vn 0.135f
C721 therm_0/_12_ Vn 0.387f
C722 therm_0/_52_/a_250_297# Vn 0.0278f
C723 therm_0/_52_/a_93_21# Vn 0.151f
C724 therm_0/_10_ Vn 0.643f
C725 therm_0/_36_/a_27_47# Vn 0.175f
C726 therm_0/input14/a_27_47# Vn 0.208f
C727 therm_0/_53_/a_29_53# Vn 0.18f
C728 therm_0/_37_/a_27_47# Vn 0.175f
C729 therm_0/input13/a_27_47# Vn 0.208f
C730 therm_0/net18 Vn 0.207f
C731 therm_0/_25_ Vn 0.191f
C732 therm_0/_54_/a_75_212# Vn 0.21f
C733 therm_0/net4 Vn 0.324f
C734 therm_0/_38_/a_27_47# Vn 0.175f
C735 therm_0/net19 Vn 0.187f
C736 therm_0/_22_ Vn 0.215f
C737 therm_0/_14_ Vn 0.228f
C738 therm_0/_15_ Vn 0.336f
C739 therm_0/_55_/a_217_297# Vn 0.00117f
C740 therm_0/_55_/a_80_21# Vn 0.21f
C741 therm_0/input12/a_27_47# Vn 0.208f
C742 therm_0/input9/a_75_212# Vn 0.21f
C743 therm_0/_39_/a_285_47# Vn 0.0174f
C744 therm_0/_39_/a_47_47# Vn 0.199f
C745 therm_0/input11/a_27_47# Vn 0.208f
C746 therm_0/input8/a_27_47# Vn 0.208f
C747 therm_0/input10/a_27_47# Vn 0.208f
C748 therm_0/net7 Vn 0.448f
C749 therm_0/input7/a_27_47# Vn 0.208f
C750 therm_0/input6/a_27_47# Vn 0.208f
C751 therm_0/net5 Vn 0.825f
C752 therm_0/input5/a_841_47# Vn 0.0929f
C753 therm_0/input5/a_664_47# Vn 0.13f
C754 therm_0/input5/a_558_47# Vn 0.164f
C755 therm_0/input5/a_381_47# Vn 0.11f
C756 therm_0/input5/a_62_47# Vn 0.169f
C757 therm_0/input4/a_75_212# Vn 0.21f
C758 therm_0/input3/a_27_47# Vn 0.208f
C759 therm_0/net2 Vn 0.811f
C760 therm_0/input2/a_27_47# Vn 0.208f
C761 therm_0/net1 Vn 0.337f
C762 Vp Vn 82.8f
C763 therm_0/input1/a_75_212# Vn 0.21f
C764 b[3] Vn 0.43f
C765 therm_0/output19/a_27_47# Vn 0.543f
C766 b[2] Vn 0.575f
C767 therm_0/output18/a_27_47# Vn 0.543f
C768 b[1] Vn 0.438f
C769 therm_0/net17 Vn 0.172f
C770 therm_0/output17/a_27_47# Vn 0.543f
C771 therm_0/_41_/a_59_75# Vn 0.177f
C772 b[0] Vn 0.619f
C773 therm_0/output16/a_27_47# Vn 0.543f
C774 therm_0/_16_ Vn 0.125f
C775 therm_0/_42_/a_209_311# Vn 0.143f
C776 therm_0/_42_/a_109_93# Vn 0.158f
C777 therm_0/_17_ Vn 0.251f
C778 therm_0/_43_/a_193_413# Vn 0.136f
C779 therm_0/_43_/a_27_47# Vn 0.224f
C780 therm_0/_00_ Vn 0.377f
C781 therm_0/net6 Vn 0.531f
C782 therm_0/_26_/a_29_53# Vn 0.18f
C783 therm_0/_01_ Vn 0.15f
C784 therm_0/net14 Vn 0.516f
C785 therm_0/net3 Vn 0.462f
C786 therm_0/net15 Vn 0.452f
C787 therm_0/_27_/a_27_297# Vn 0.163f
C788 therm_0/_18_ Vn 0.143f
C789 therm_0/_44_/a_250_297# Vn 0.0278f
C790 therm_0/_44_/a_93_21# Vn 0.151f
C791 therm_0/net16 Vn 0.231f
C792 therm_0/_13_ Vn 0.133f
C793 therm_0/_45_/a_193_297# Vn 0.0011f
C794 therm_0/_45_/a_109_297# Vn 7.11e-19
C795 therm_0/_45_/a_27_47# Vn 0.216f
C796 therm_0/net12 Vn 0.517f
C797 therm_0/net13 Vn 0.377f
C798 therm_0/_29_/a_29_53# Vn 0.18f
C799 therm_0/_19_ Vn 0.118f
C800 therm_0/_47_/a_299_297# Vn 0.0348f
C801 therm_0/_47_/a_81_21# Vn 0.147f
C802 therm_0/_48_/a_27_47# Vn 0.177f
C803 therm_0/_21_ Vn 0.29f
C804 therm_0/_20_ Vn 0.235f
C805 therm_0/_02_ Vn 0.45f
C806 therm_0/_49_/a_201_297# Vn 0.00345f
C807 therm_0/_49_/a_75_199# Vn 0.205f
C808 th08_0/m1_477_n803# Vn 0.582f
C809 V08 Vn 0.788f
C810 V15 Vn 1.68f
C811 th15_0/m1_849_n157# Vn 1.32f
C812 th15_0/m1_597_n912# Vn 0.294f
C813 V01 Vn 1.05f
C814 th01_0/m1_991_n1219# Vn 1.24f
C815 th01_0/m1_571_n501# Vn 0.197f
C816 th15_0/Vin Vn 6.9f
C817 th03_0/m1_890_n844# Vn 1.05f
C818 V03 Vn 1.6f
C819 th03_0/m1_638_n591# Vn 0.234f
C820 th10_0/m1_536_174# Vn 0.882f
C821 V10 Vn 0.383f
C822 th10_0/m1_502_n495# Vn 0.156f
C823 th05_0/m1_752_n794# Vn 0.796f
C824 V05 Vn 1.02f
C825 th12_0/m1_529_n42# Vn 0.933f
C826 V12 Vn 0.582f
C827 th12_0/m1_394_n856# Vn 0.219f
C828 th07_0/m1_808_n892# Vn 0.523f
C829 V07 Vn 0.828f
C830 V14 Vn 0.81f
C831 th14_0/m1_891_419# Vn 1.52f
C832 th14_0/m1_641_n318# Vn 0.281f
C833 th09_0/m1_485_n505# Vn 1.24f
C834 V09 Vn 1.74f
C835 th09_0/m1_962_372# Vn 0.124f
C836 V02 Vn 1.63f
C837 th02_0/m1_983_133# Vn 1.6f
C838 th02_0/m1_571_144# Vn 0.267f
.ends

