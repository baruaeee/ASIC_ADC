magic
tech sky130A
timestamp 1703732895
<< pwell >>
rect -698 -126 698 126
<< nmos >>
rect -600 -21 600 21
<< ndiff >>
rect -629 15 -600 21
rect -629 -15 -623 15
rect -606 -15 -600 15
rect -629 -21 -600 -15
rect 600 15 629 21
rect 600 -15 606 15
rect 623 -15 629 15
rect 600 -21 629 -15
<< ndiffc >>
rect -623 -15 -606 15
rect 606 -15 623 15
<< psubdiff >>
rect -680 91 -632 108
rect 632 91 680 108
rect -680 60 -663 91
rect 663 60 680 91
rect -680 -91 -663 -60
rect 663 -91 680 -60
rect -680 -108 -632 -91
rect 632 -108 680 -91
<< psubdiffcont >>
rect -632 91 632 108
rect -680 -60 -663 60
rect 663 -60 680 60
rect -632 -108 632 -91
<< poly >>
rect -600 57 600 65
rect -600 40 -592 57
rect 592 40 600 57
rect -600 21 600 40
rect -600 -40 600 -21
rect -600 -57 -592 -40
rect 592 -57 600 -40
rect -600 -65 600 -57
<< polycont >>
rect -592 40 592 57
rect -592 -57 592 -40
<< locali >>
rect -680 91 -632 108
rect 632 91 680 108
rect -680 60 -663 91
rect 663 60 680 91
rect -600 40 -592 57
rect 592 40 600 57
rect -623 15 -606 23
rect -623 -23 -606 -15
rect 606 15 623 23
rect 606 -23 623 -15
rect -600 -57 -592 -40
rect 592 -57 600 -40
rect -680 -91 -663 -60
rect 663 -91 680 -60
rect -680 -108 -632 -91
rect 632 -108 680 -91
<< viali >>
rect -592 40 592 57
rect -623 -15 -606 15
rect 606 -15 623 15
rect -592 -57 592 -40
<< metal1 >>
rect -598 57 598 60
rect -598 40 -592 57
rect 592 40 598 57
rect -598 37 598 40
rect -626 15 -603 21
rect -626 -15 -623 15
rect -606 -15 -603 15
rect -626 -21 -603 -15
rect 603 15 626 21
rect 603 -15 606 15
rect 623 -15 626 15
rect 603 -21 626 -15
rect -598 -40 598 -37
rect -598 -57 -592 -40
rect 592 -57 598 -40
rect -598 -60 598 -57
<< properties >>
string FIXED_BBOX -671 -99 671 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 12.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
