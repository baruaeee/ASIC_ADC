magic
tech sky130A
timestamp 1704501257
<< pwell >>
rect -648 -126 648 126
<< nmos >>
rect -550 -21 550 21
<< ndiff >>
rect -579 15 -550 21
rect -579 -15 -573 15
rect -556 -15 -550 15
rect -579 -21 -550 -15
rect 550 15 579 21
rect 550 -15 556 15
rect 573 -15 579 15
rect 550 -21 579 -15
<< ndiffc >>
rect -573 -15 -556 15
rect 556 -15 573 15
<< psubdiff >>
rect -630 91 -582 108
rect 582 91 630 108
rect -630 60 -613 91
rect 613 60 630 91
rect -630 -91 -613 -60
rect 613 -91 630 -60
rect -630 -108 -582 -91
rect 582 -108 630 -91
<< psubdiffcont >>
rect -582 91 582 108
rect -630 -60 -613 60
rect 613 -60 630 60
rect -582 -108 582 -91
<< poly >>
rect -550 57 550 65
rect -550 40 -542 57
rect 542 40 550 57
rect -550 21 550 40
rect -550 -40 550 -21
rect -550 -57 -542 -40
rect 542 -57 550 -40
rect -550 -65 550 -57
<< polycont >>
rect -542 40 542 57
rect -542 -57 542 -40
<< locali >>
rect -630 91 -582 108
rect 582 91 630 108
rect -630 60 -613 91
rect 613 60 630 91
rect -550 40 -542 57
rect 542 40 550 57
rect -573 15 -556 23
rect -573 -23 -556 -15
rect 556 15 573 23
rect 556 -23 573 -15
rect -550 -57 -542 -40
rect 542 -57 550 -40
rect -630 -91 -613 -60
rect 613 -91 630 -60
rect -630 -108 -582 -91
rect 582 -108 630 -91
<< viali >>
rect -542 40 542 57
rect -573 -15 -556 15
rect 556 -15 573 15
rect -542 -57 542 -40
<< metal1 >>
rect -548 57 548 60
rect -548 40 -542 57
rect 542 40 548 57
rect -548 37 548 40
rect -576 15 -553 21
rect -576 -15 -573 15
rect -556 -15 -553 15
rect -576 -21 -553 -15
rect 553 15 576 21
rect 553 -15 556 15
rect 573 -15 576 15
rect 553 -21 576 -15
rect -548 -40 548 -37
rect -548 -57 -542 -40
rect 542 -57 548 -40
rect -548 -60 548 -57
<< properties >>
string FIXED_BBOX -621 -99 621 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 11.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
