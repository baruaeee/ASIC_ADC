magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< nwell >>
rect -354 -261 354 261
<< pmos >>
rect -158 -42 158 42
<< pdiff >>
rect -216 30 -158 42
rect -216 -30 -204 30
rect -170 -30 -158 30
rect -216 -42 -158 -30
rect 158 30 216 42
rect 158 -30 170 30
rect 204 -30 216 30
rect 158 -42 216 -30
<< pdiffc >>
rect -204 -30 -170 30
rect 170 -30 204 30
<< nsubdiff >>
rect -318 191 -222 225
rect 222 191 318 225
rect -318 129 -284 191
rect 284 129 318 191
rect -318 -191 -284 -129
rect 284 -191 318 -129
rect -318 -225 -222 -191
rect 222 -225 318 -191
<< nsubdiffcont >>
rect -222 191 222 225
rect -318 -129 -284 129
rect 284 -129 318 129
rect -222 -225 222 -191
<< poly >>
rect -158 123 158 139
rect -158 89 -142 123
rect 142 89 158 123
rect -158 42 158 89
rect -158 -89 158 -42
rect -158 -123 -142 -89
rect 142 -123 158 -89
rect -158 -139 158 -123
<< polycont >>
rect -142 89 142 123
rect -142 -123 142 -89
<< locali >>
rect -318 191 -222 225
rect 222 191 318 225
rect -318 129 -284 191
rect 284 129 318 191
rect -158 89 -142 123
rect 142 89 158 123
rect -204 30 -170 46
rect -204 -46 -170 -30
rect 170 30 204 46
rect 170 -46 204 -30
rect -158 -123 -142 -89
rect 142 -123 158 -89
rect -318 -191 -284 -129
rect 284 -191 318 -129
rect -318 -225 -222 -191
rect 222 -225 318 -191
<< viali >>
rect -142 89 142 123
rect -204 -30 -170 30
rect 170 -30 204 30
rect -142 -123 142 -89
<< metal1 >>
rect -154 123 154 129
rect -154 89 -142 123
rect 142 89 154 123
rect -154 83 154 89
rect -210 30 -164 42
rect -210 -30 -204 30
rect -170 -30 -164 30
rect -210 -42 -164 -30
rect 164 30 210 42
rect 164 -30 170 30
rect 204 -30 210 30
rect 164 -42 210 -30
rect -154 -89 154 -83
rect -154 -123 -142 -89
rect 142 -123 154 -89
rect -154 -129 154 -123
<< properties >>
string FIXED_BBOX -301 -208 301 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 1.58 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
