magic
tech sky130A
magscale 1 2
timestamp 1706239161
<< error_p >>
rect -29 123 29 129
rect -29 89 -17 123
rect -29 83 29 89
rect -29 -89 29 -83
rect -29 -123 -17 -89
rect -29 -129 29 -123
<< nwell >>
rect -224 -261 224 261
<< pmos >>
rect -28 -42 28 42
<< pdiff >>
rect -86 30 -28 42
rect -86 -30 -74 30
rect -40 -30 -28 30
rect -86 -42 -28 -30
rect 28 30 86 42
rect 28 -30 40 30
rect 74 -30 86 30
rect 28 -42 86 -30
<< pdiffc >>
rect -74 -30 -40 30
rect 40 -30 74 30
<< nsubdiff >>
rect -154 191 -92 225
rect 92 191 154 225
<< nsubdiffcont >>
rect -92 191 92 225
<< poly >>
rect -33 123 33 139
rect -33 89 -17 123
rect 17 89 33 123
rect -33 73 33 89
rect -28 42 28 73
rect -28 -73 28 -42
rect -33 -89 33 -73
rect -33 -123 -17 -89
rect 17 -123 33 -89
rect -33 -139 33 -123
<< polycont >>
rect -17 89 17 123
rect -17 -123 17 -89
<< locali >>
rect -154 191 -92 225
rect 92 191 154 225
rect -33 89 -17 123
rect 17 89 33 123
rect -74 30 -40 46
rect -74 -46 -40 -30
rect 40 30 74 46
rect 40 -46 74 -30
rect -33 -123 -17 -89
rect 17 -123 33 -89
<< viali >>
rect -17 89 17 123
rect -74 -30 -40 30
rect 40 -30 74 30
rect -17 -123 17 -89
<< metal1 >>
rect -29 123 29 129
rect -29 89 -17 123
rect 17 89 29 123
rect -29 83 29 89
rect -80 30 -34 42
rect -80 -30 -74 30
rect -40 -30 -34 30
rect -80 -42 -34 -30
rect 34 30 80 42
rect 34 -30 40 30
rect 74 -30 80 30
rect 34 -42 80 -30
rect -29 -89 29 -83
rect -29 -123 -17 -89
rect 17 -123 29 -89
rect -29 -129 29 -123
<< properties >>
string FIXED_BBOX -171 -208 171 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.28 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
