


.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n34_n198#
+ VSUBS
X0 a_15_n100# a_n34_n198# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_15_n100# w_n211_n319# 0.0808f
C1 w_n211_n319# a_n34_n198# 0.272f
C2 a_n73_n100# w_n211_n319# 0.0808f
C3 a_15_n100# a_n34_n198# 0.0287f
C4 a_n73_n100# a_15_n100# 0.162f
C5 a_n73_n100# a_n34_n198# 0.0287f
C6 a_15_n100# VSUBS 0.0484f
C7 a_n73_n100# VSUBS 0.0484f
C8 a_n34_n198# VSUBS 0.118f
C9 w_n211_n319# VSUBS 1.23f
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n34_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n34_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n34_n188# a_n73_n100# 0.0309f
C1 a_15_n100# a_n34_n188# 0.0309f
C2 a_15_n100# a_n73_n100# 0.162f
C3 a_15_n100# a_n175_n274# 0.129f
C4 a_n73_n100# a_n175_n274# 0.129f
C5 a_n34_n188# a_n175_n274# 0.373f
.ends



VDD VDD GND 1.8
.save i(vdd)
Vin Vin GND pulse(0 1.8 0ns 1ns 1ns 5ns 10ns)
.save i(vin)
x1 VDD Vin Vout GND make_symbol_Inverter
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.save all





.tran 1n 30n
.control
run
set color0=white
set color1=black
plot Vin Vout
set xbrushwidth=3
.save all
.endc
.end


**** end user architecture code
**.ends


.subckt make_symbol_Inverter Vdd Vin Vout GND

XXM1 Vdd Vout XM1/w_n211_n319# GND VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM2 GND GND Vout VSUBS sky130_fd_pr__nfet_01v8_648S5X
C0 GND Vout 0.0548f
C1 Vdd XM1/w_n211_n319# 0.0888f
C2 Vout XM1/w_n211_n319# 0.087f
C3 Vdd Vout 0.00927f
C4 GND XM1/w_n211_n319# 0.0564f
C5 Vdd GND 0.16f
C6 Vout VSUBS 0.612f
C7 GND VSUBS 1.28f
C8 Vdd VSUBS 0.39f
C9 XM1/w_n211_n319# VSUBS 1.29f
.ends

.end
