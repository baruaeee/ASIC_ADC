magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 311 29 317
rect -29 277 -17 311
rect -29 271 29 277
rect -29 -277 29 -271
rect -29 -311 -17 -277
rect -29 -317 29 -311
<< nwell >>
rect -211 -449 211 449
<< pmos >>
rect -15 -230 15 230
<< pdiff >>
rect -73 218 -15 230
rect -73 -218 -61 218
rect -27 -218 -15 218
rect -73 -230 -15 -218
rect 15 218 73 230
rect 15 -218 27 218
rect 61 -218 73 218
rect 15 -230 73 -218
<< pdiffc >>
rect -61 -218 -27 218
rect 27 -218 61 218
<< nsubdiff >>
rect -175 379 -79 413
rect 79 379 175 413
rect -175 317 -141 379
rect 141 317 175 379
rect -175 -379 -141 -317
rect 141 -379 175 -317
rect -175 -413 -79 -379
rect 79 -413 175 -379
<< nsubdiffcont >>
rect -79 379 79 413
rect -175 -317 -141 317
rect 141 -317 175 317
rect -79 -413 79 -379
<< poly >>
rect -33 311 33 327
rect -33 277 -17 311
rect 17 277 33 311
rect -33 261 33 277
rect -15 230 15 261
rect -15 -261 15 -230
rect -33 -277 33 -261
rect -33 -311 -17 -277
rect 17 -311 33 -277
rect -33 -327 33 -311
<< polycont >>
rect -17 277 17 311
rect -17 -311 17 -277
<< locali >>
rect -175 379 -79 413
rect 79 379 175 413
rect -175 317 -141 379
rect 141 317 175 379
rect -33 277 -17 311
rect 17 277 33 311
rect -61 218 -27 234
rect -61 -234 -27 -218
rect 27 218 61 234
rect 27 -234 61 -218
rect -33 -311 -17 -277
rect 17 -311 33 -277
rect -175 -379 -141 -317
rect 141 -379 175 -317
rect -175 -413 -79 -379
rect 79 -413 175 -379
<< viali >>
rect -17 277 17 311
rect -61 -218 -27 218
rect 27 -218 61 218
rect -17 -311 17 -277
<< metal1 >>
rect -29 311 29 317
rect -29 277 -17 311
rect 17 277 29 311
rect -29 271 29 277
rect -67 218 -21 230
rect -67 -218 -61 218
rect -27 -218 -21 218
rect -67 -230 -21 -218
rect 21 218 67 230
rect 21 -218 27 218
rect 61 -218 67 218
rect 21 -230 67 -218
rect -29 -277 29 -271
rect -29 -311 -17 -277
rect 17 -311 29 -277
rect -29 -317 29 -311
<< properties >>
string FIXED_BBOX -158 -396 158 396
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.3 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
