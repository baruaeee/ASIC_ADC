* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : pre_therm1                                   *
* Netlisted  : Wed Dec 11 23:18:08 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3M4_C_CDNS_733955477490                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3M4_C_CDNS_733955477490 1
** N=1 EP=1 FDC=0
.ends M3M4_C_CDNS_733955477490

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_C_CDNS_733955477491                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_C_CDNS_733955477491 1
** N=1 EP=1 FDC=0
.ends M1M2_C_CDNS_733955477491

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2M3_C_CDNS_733955477492                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2M3_C_CDNS_733955477492 1
** N=1 EP=1 FDC=0
.ends M2M3_C_CDNS_733955477492

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_C_CDNS_733955477493                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_C_CDNS_733955477493 1
** N=1 EP=1 FDC=0
.ends M1M2_C_CDNS_733955477493

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_733955477494                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_733955477494 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_733955477494

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_733955477495                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_733955477495 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_733955477495

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: PYL1CON_C_CDNS_733955477496                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt PYL1CON_C_CDNS_733955477496 1 2
** N=2 EP=2 FDC=0
.ends PYL1CON_C_CDNS_733955477496

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733955477490                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733955477490 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3.3e-07 W=8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733955477490

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733955477491                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733955477491 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733955477491

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv12f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv12f 1 2 3 4 5
** N=9 EP=5 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=465 2185 0 0 $X=300 $Y=2040
X1 4 L1M1_C_CDNS_733955477495 $T=675 3150 0 0 $X=560 $Y=2805
X2 4 L1M1_C_CDNS_733955477495 $T=810 965 0 0 $X=695 $Y=620
X3 3 6 PYL1CON_C_CDNS_733955477496 $T=465 2185 0 0 $X=280 $Y=2000
X4 2 4 3 nfet_01v8_CDNS_733955477490 $T=340 555 0 0 $X=-65 $Y=405
X5 1 4 3 pfet_01v8_CDNS_733955477491 $T=385 2785 0 0 $X=-60 $Y=2605
.ends inv12f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_733955477497                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_733955477497 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_733955477497

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733955477492                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733955477492 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=9.5e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733955477492

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733955477493                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733955477493 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733955477493

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv15f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv15f 1 2 3 4 5
** N=9 EP=5 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=700 1765 0 0 $X=535 $Y=1620
X1 4 L1M1_C_CDNS_733955477495 $T=910 3070 0 0 $X=795 $Y=2725
X2 3 6 PYL1CON_C_CDNS_733955477496 $T=700 1765 0 0 $X=515 $Y=1580
X3 4 L1M1_C_CDNS_733955477497 $T=1305 910 0 0 $X=1190 $Y=745
X4 2 4 3 nfet_01v8_CDNS_733955477492 $T=215 700 0 0 $X=-190 $Y=550
X5 1 4 3 pfet_01v8_CDNS_733955477493 $T=620 2635 0 0 $X=175 $Y=2455
.ends inv15f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733955477494                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733955477494 1 2 3
** N=7 EP=3 FDC=1
M0 2 2 1 3 pfet_01v8 L=1.5e-07 W=1e-06 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733955477494

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733955477495                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733955477495 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 pfet_01v8 L=1.05e-06 W=5.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733955477495

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: div_fixed                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt div_fixed 1 2 3 4 5
** N=8 EP=5 FDC=2
X0 2 L1M1_C_CDNS_733955477494 $T=390 585 0 0 $X=225 $Y=440
X1 3 L1M1_C_CDNS_733955477495 $T=610 1390 0 0 $X=495 $Y=1045
X2 2 6 PYL1CON_C_CDNS_733955477496 $T=405 585 0 0 $X=220 $Y=400
X3 3 L1M1_C_CDNS_733955477497 $T=1350 2690 0 90 $X=1185 $Y=2575
X4 3 2 1 pfet_01v8_CDNS_733955477494 $T=470 1900 0 180 $X=-125 $Y=720
X5 1 3 2 1 pfet_01v8_CDNS_733955477495 $T=1625 3880 1 270 $X=895 $Y=2385
.ends div_fixed

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733955477496                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733955477496 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6.75e-07 W=4.8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733955477496

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733955477497                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733955477497 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.65e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733955477497

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv14f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv14f 1 2 3 4 5 6
** N=9 EP=6 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=520 1745 0 0 $X=355 $Y=1600
X1 4 L1M1_C_CDNS_733955477495 $T=735 3095 0 0 $X=620 $Y=2750
X2 3 7 PYL1CON_C_CDNS_733955477496 $T=520 1745 0 0 $X=335 $Y=1560
X3 4 L1M1_C_CDNS_733955477497 $T=1165 915 0 0 $X=1050 $Y=750
X4 2 4 3 nfet_01v8_CDNS_733955477496 $T=350 675 0 0 $X=-55 $Y=525
X5 1 4 3 pfet_01v8_CDNS_733955477497 $T=445 2705 0 0 $X=0 $Y=2525
.ends inv14f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733955477498                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733955477498 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.6e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733955477498

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv11f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv11f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=480 1765 0 0 $X=315 $Y=1620
X1 4 L1M1_C_CDNS_733955477495 $T=750 3045 0 0 $X=635 $Y=2700
X2 3 5 PYL1CON_C_CDNS_733955477496 $T=480 1765 0 0 $X=295 $Y=1580
X3 4 L1M1_C_CDNS_733955477497 $T=1305 910 0 0 $X=1190 $Y=745
X4 2 4 3 nfet_01v8_CDNS_733955477492 $T=215 700 0 0 $X=-190 $Y=550
X5 1 4 3 pfet_01v8_CDNS_733955477498 $T=350 2610 0 0 $X=-95 $Y=2430
.ends inv11f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733955477499                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733955477499 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.55e-07 W=9.45e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733955477499

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774910                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774910 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.45e-07 W=8.65e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774910

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv10f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv10f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=500 1860 0 0 $X=335 $Y=1715
X1 4 L1M1_C_CDNS_733955477495 $T=720 1035 0 0 $X=605 $Y=690
X2 4 L1M1_C_CDNS_733955477495 $T=770 3090 0 0 $X=655 $Y=2745
X3 3 5 PYL1CON_C_CDNS_733955477496 $T=500 1860 0 0 $X=315 $Y=1675
X4 2 4 3 nfet_01v8_CDNS_733955477499 $T=425 555 0 0 $X=20 $Y=405
X5 1 4 3 pfet_01v8_CDNS_7339554774910 $T=385 2670 0 0 $X=-60 $Y=2490
.ends inv10f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774911                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774911 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=9.9e-07 W=4.9e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774911

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774912                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774912 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.65e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774912

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv08f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv08f 1 2 3 4 5 6
** N=9 EP=6 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=155 1745 0 0 $X=-10 $Y=1600
X1 4 L1M1_C_CDNS_733955477495 $T=665 3170 0 0 $X=550 $Y=2825
X2 3 7 PYL1CON_C_CDNS_733955477496 $T=155 1745 0 0 $X=-30 $Y=1560
X3 4 L1M1_C_CDNS_733955477497 $T=1035 1870 0 90 $X=870 $Y=1755
X4 2 4 3 nfet_01v8_CDNS_7339554774911 $T=1280 740 0 90 $X=640 $Y=335
X5 1 4 3 pfet_01v8_CDNS_7339554774912 $T=360 2755 0 0 $X=-85 $Y=2575
.ends inv08f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774913                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774913 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=6.95e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774913

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774914                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774914 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=4e-07 W=6.5e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774914

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv05f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv05f 1 2 3 4 5 6
** N=9 EP=6 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=510 1810 0 0 $X=345 $Y=1665
X1 4 L1M1_C_CDNS_733955477495 $T=650 3170 0 0 $X=535 $Y=2825
X2 4 L1M1_C_CDNS_733955477495 $T=855 960 0 0 $X=740 $Y=615
X3 3 7 PYL1CON_C_CDNS_733955477496 $T=510 1810 0 0 $X=325 $Y=1625
X4 1 4 3 pfet_01v8_CDNS_7339554774913 $T=360 2825 0 0 $X=-85 $Y=2645
X5 2 4 3 nfet_01v8_CDNS_7339554774914 $T=315 630 0 0 $X=-90 $Y=480
.ends inv05f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774915                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774915 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.5e-07 W=8e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774915

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774916                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774916 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=2.85e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774916

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv02f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv02f 1 2 3 4 5 6
** N=9 EP=6 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=460 1630 0 0 $X=295 $Y=1485
X1 4 L1M1_C_CDNS_733955477495 $T=725 3245 0 0 $X=610 $Y=2900
X2 3 7 PYL1CON_C_CDNS_733955477496 $T=460 1630 0 0 $X=275 $Y=1445
X3 4 L1M1_C_CDNS_733955477497 $T=740 850 0 0 $X=625 $Y=685
X4 1 4 3 pfet_01v8_CDNS_7339554774915 $T=335 2855 0 0 $X=-110 $Y=2675
X5 2 4 3 nfet_01v8_CDNS_7339554774916 $T=315 640 0 0 $X=-90 $Y=490
.ends inv02f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774917                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774917 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3e-07 W=9.8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774917

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774918                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774918 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.55e-07 W=5.7e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774918

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv07f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv07f 1 2 3 4 5 6
** N=9 EP=6 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=435 2320 0 0 $X=270 $Y=2175
X1 4 L1M1_C_CDNS_733955477495 $T=755 940 0 0 $X=640 $Y=595
X2 3 7 PYL1CON_C_CDNS_733955477496 $T=435 2320 0 0 $X=250 $Y=2135
X3 4 L1M1_C_CDNS_733955477497 $T=655 3235 0 0 $X=540 $Y=3070
X4 2 4 3 nfet_01v8_CDNS_7339554774917 $T=315 460 0 0 $X=-90 $Y=310
X5 1 4 3 pfet_01v8_CDNS_7339554774918 $T=360 2950 0 0 $X=-85 $Y=2770
.ends inv07f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774919                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774919 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.9e-07 W=6.2e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774919

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774920                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774920 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6e-07 W=7.05e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774920

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv04f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv04f 1 2 3 4 5 6
** N=9 EP=6 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=575 1030 0 0 $X=410 $Y=885
X1 4 L1M1_C_CDNS_733955477495 $T=710 2960 0 0 $X=595 $Y=2615
X2 4 L1M1_C_CDNS_733955477495 $T=1025 1070 0 0 $X=910 $Y=725
X3 3 7 PYL1CON_C_CDNS_733955477496 $T=575 1030 0 0 $X=390 $Y=845
X4 1 4 3 pfet_01v8_CDNS_7339554774919 $T=380 2650 0 0 $X=-65 $Y=2470
X5 2 4 3 nfet_01v8_CDNS_7339554774920 $T=280 715 0 0 $X=-125 $Y=565
.ends inv04f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774921                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774921 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=5.5e-07 W=5.4e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774921

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774922                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774922 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.6e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774922

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv13f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv13f 1 2 3 4 5 6 7
** N=9 EP=7 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=465 1790 0 0 $X=300 $Y=1645
X1 4 L1M1_C_CDNS_733955477495 $T=685 3120 0 0 $X=570 $Y=2775
X2 3 8 PYL1CON_C_CDNS_733955477496 $T=465 1790 0 0 $X=280 $Y=1605
X3 4 L1M1_C_CDNS_733955477497 $T=1050 915 0 0 $X=935 $Y=750
X4 2 4 3 nfet_01v8_CDNS_7339554774921 $T=360 720 0 0 $X=-45 $Y=570
X5 1 4 3 pfet_01v8_CDNS_7339554774922 $T=385 2685 0 0 $X=-60 $Y=2505
.ends inv13f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774923                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774923 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.1e-06 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774923

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774924                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774924 1 2 3
** N=9 EP=3 FDC=2
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.7e-07 $X=0 $Y=0 $dt=8
M1 1 3 2 1 pfet_01v8 L=1.5e-07 W=7.7e-07 $X=430 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774924

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv09f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv09f 1 2 3 4 5
** N=9 EP=5 FDC=3
X0 3 L1M1_C_CDNS_733955477494 $T=20 2075 0 0 $X=-145 $Y=1930
X1 3 6 PYL1CON_C_CDNS_733955477496 $T=20 2075 0 0 $X=-165 $Y=1890
X2 4 L1M1_C_CDNS_733955477497 $T=670 1935 0 90 $X=505 $Y=1820
X3 4 L1M1_C_CDNS_733955477497 $T=690 3225 0 0 $X=575 $Y=3060
X4 2 4 3 nfet_01v8_CDNS_7339554774923 $T=905 695 0 90 $X=335 $Y=290
X5 1 4 3 pfet_01v8_CDNS_7339554774924 $T=400 2840 0 0 $X=-45 $Y=2660
.ends inv09f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774925                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774925 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3.2e-07 W=7.25e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774925

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774926                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774926 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=4.35e-07 W=5.6e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774926

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv06f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv06f 1 2 3 4 5 6 7 8
** N=9 EP=8 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=555 2320 0 0 $X=390 $Y=2175
X1 4 L1M1_C_CDNS_733955477495 $T=855 1035 0 0 $X=740 $Y=690
X2 3 9 PYL1CON_C_CDNS_733955477496 $T=555 2320 0 0 $X=370 $Y=2135
X3 4 L1M1_C_CDNS_733955477497 $T=910 3285 0 0 $X=795 $Y=3120
X4 2 4 3 nfet_01v8_CDNS_7339554774925 $T=395 685 0 0 $X=-10 $Y=535
X5 1 4 3 pfet_01v8_CDNS_7339554774926 $T=335 3005 0 0 $X=-110 $Y=2825
.ends inv06f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774927                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774927 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=3.5e-07 W=6.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774927

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774928                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774928 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=4.5e-07 W=6.4e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774928

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv03f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv03f 1 2 3 4 5
** N=9 EP=5 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=510 1870 0 0 $X=345 $Y=1725
X1 4 L1M1_C_CDNS_733955477495 $T=825 3370 0 0 $X=710 $Y=3025
X2 4 L1M1_C_CDNS_733955477495 $T=880 960 0 0 $X=765 $Y=615
X3 3 6 PYL1CON_C_CDNS_733955477496 $T=510 1870 0 0 $X=325 $Y=1685
X4 1 4 3 pfet_01v8_CDNS_7339554774927 $T=335 3045 0 0 $X=-110 $Y=2865
X5 2 4 3 nfet_01v8_CDNS_7339554774928 $T=290 640 0 0 $X=-115 $Y=490
.ends inv03f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774929                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774929 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6.5e-07 W=4.45e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774929

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774930                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774930 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=6.3e-07 W=7.9e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774930

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv01f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv01f 1 2 3 4 5 6
** N=9 EP=6 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=575 1630 0 0 $X=410 $Y=1485
X1 4 L1M1_C_CDNS_733955477495 $T=1065 3205 0 0 $X=950 $Y=2860
X2 3 7 PYL1CON_C_CDNS_733955477496 $T=575 1630 0 0 $X=390 $Y=1445
X3 4 L1M1_C_CDNS_733955477497 $T=1085 695 0 0 $X=970 $Y=530
X4 2 4 3 nfet_01v8_CDNS_7339554774929 $T=295 475 0 0 $X=-110 $Y=325
X5 1 4 3 pfet_01v8_CDNS_7339554774930 $T=295 2820 0 0 $X=-150 $Y=2640
.ends inv01f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339554774931                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339554774931 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 pfet_01v8 L=2.5e-07 W=5.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339554774931

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774932                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774932 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 nfet_01v8 L=5.5e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774932

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: preamp1F                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt preamp1F 1 2 3 4 5
** N=9 EP=5 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=810 990 0 0 $X=645 $Y=845
X1 4 L1M1_C_CDNS_733955477495 $T=725 1970 0 0 $X=610 $Y=1625
X2 3 6 PYL1CON_C_CDNS_733955477496 $T=810 990 0 0 $X=625 $Y=805
X3 4 2 3 1 pfet_01v8_CDNS_7339554774931 $T=840 2840 0 90 $X=110 $Y=2395
X4 4 1 3 2 nfet_01v8_CDNS_7339554774932 $T=610 1275 0 270 $X=460 $Y=320
.ends preamp1F

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_733955477498                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_733955477498 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_733955477498

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339554774933                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339554774933 1 2 3 4
** N=10 EP=4 FDC=1
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=1.02e-06 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339554774933

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: preampF                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt preampF 1 2 3 4 5 6
** N=9 EP=6 FDC=2
X0 3 L1M1_C_CDNS_733955477494 $T=415 2135 0 0 $X=250 $Y=1990
X1 3 7 PYL1CON_C_CDNS_733955477496 $T=415 2135 0 0 $X=230 $Y=1950
X2 4 L1M1_C_CDNS_733955477497 $T=1100 3570 0 90 $X=935 $Y=3455
X3 4 2 3 1 pfet_01v8_CDNS_733955477495 $T=825 3430 0 270 $X=645 $Y=1935
X4 1 L1M1_C_CDNS_733955477498 $T=130 995 0 0 $X=15 $Y=470
X5 4 L1M1_C_CDNS_733955477498 $T=570 995 0 0 $X=455 $Y=470
X6 4 1 3 2 nfet_01v8_CDNS_7339554774933 $T=430 485 1 180 $X=-125 $Y=335
.ends preampF

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pre_therm1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pre_therm1 2 6 7 14 16 18 3 5 8 11
+ 10 12 15 17 19
** N=37 EP=15 FDC=37
X0 1 M3M4_C_CDNS_733955477490 $T=10420 4140 0 0 $X=10055 $Y=3950
X1 1 M3M4_C_CDNS_733955477490 $T=10420 12420 0 0 $X=10055 $Y=12230
X2 2 M1M2_C_CDNS_733955477491 $T=-550 6305 0 0 $X=-680 $Y=6145
X3 2 M1M2_C_CDNS_733955477491 $T=390 2575 0 90 $X=230 $Y=2445
X4 2 M1M2_C_CDNS_733955477491 $T=530 6015 0 90 $X=370 $Y=5885
X5 3 M1M2_C_CDNS_733955477491 $T=900 7460 0 90 $X=740 $Y=7330
X6 2 M1M2_C_CDNS_733955477491 $T=2010 5985 0 0 $X=1880 $Y=5825
X7 4 M1M2_C_CDNS_733955477491 $T=2260 2040 0 0 $X=2130 $Y=1880
X8 5 M1M2_C_CDNS_733955477491 $T=2400 7525 0 0 $X=2270 $Y=7365
X9 6 M1M2_C_CDNS_733955477491 $T=2730 685 0 0 $X=2600 $Y=525
X10 2 M1M2_C_CDNS_733955477491 $T=3360 6510 0 0 $X=3230 $Y=6350
X11 4 M1M2_C_CDNS_733955477491 $T=3665 2040 0 0 $X=3535 $Y=1880
X12 7 M1M2_C_CDNS_733955477491 $T=4015 845 0 0 $X=3885 $Y=685
X13 8 M1M2_C_CDNS_733955477491 $T=4260 6685 0 0 $X=4130 $Y=6525
X14 9 M1M2_C_CDNS_733955477491 $T=4635 10115 0 0 $X=4505 $Y=9955
X15 10 M1M2_C_CDNS_733955477491 $T=4865 11555 0 0 $X=4735 $Y=11395
X16 2 M1M2_C_CDNS_733955477491 $T=4920 5985 0 0 $X=4790 $Y=5825
X17 2 M1M2_C_CDNS_733955477491 $T=5230 1015 0 0 $X=5100 $Y=855
X18 11 M1M2_C_CDNS_733955477491 $T=5625 6620 0 0 $X=5495 $Y=6460
X19 9 M1M2_C_CDNS_733955477491 $T=6200 10115 0 0 $X=6070 $Y=9955
X20 12 M1M2_C_CDNS_733955477491 $T=6540 11510 0 0 $X=6410 $Y=11350
X21 13 M1M2_C_CDNS_733955477491 $T=6835 1845 0 0 $X=6705 $Y=1685
X22 9 M1M2_C_CDNS_733955477491 $T=6995 6120 0 0 $X=6865 $Y=5960
X23 14 M1M2_C_CDNS_733955477491 $T=7165 775 0 0 $X=7035 $Y=615
X24 15 M1M2_C_CDNS_733955477491 $T=7610 4890 0 90 $X=7450 $Y=4760
X25 9 M1M2_C_CDNS_733955477491 $T=8375 6465 0 0 $X=8245 $Y=6305
X26 13 M1M2_C_CDNS_733955477491 $T=8420 1055 0 0 $X=8290 $Y=895
X27 16 M1M2_C_CDNS_733955477491 $T=8940 885 0 0 $X=8810 $Y=725
X28 17 M1M2_C_CDNS_733955477491 $T=8975 5590 0 90 $X=8815 $Y=5460
X29 13 M1M2_C_CDNS_733955477491 $T=9860 1845 0 0 $X=9730 $Y=1685
X30 9 M1M2_C_CDNS_733955477491 $T=9900 6480 0 90 $X=9740 $Y=6350
X31 18 M1M2_C_CDNS_733955477491 $T=10550 745 0 90 $X=10390 $Y=615
X32 19 M1M2_C_CDNS_733955477491 $T=10615 7430 0 90 $X=10455 $Y=7300
X33 20 M2M3_C_CDNS_733955477492 $T=9415 8280 0 0 $X=9050 $Y=8095
X34 20 M2M3_C_CDNS_733955477492 $T=9640 0 0 0 $X=9275 $Y=-185
X35 1 M2M3_C_CDNS_733955477492 $T=10415 4140 0 0 $X=10050 $Y=3955
X36 1 M2M3_C_CDNS_733955477492 $T=10415 12420 0 0 $X=10050 $Y=12235
X37 20 M1M2_C_CDNS_733955477493 $T=9410 8280 0 0 $X=9120 $Y=8120
X38 20 M1M2_C_CDNS_733955477493 $T=9635 0 0 0 $X=9345 $Y=-160
X39 1 M1M2_C_CDNS_733955477493 $T=10465 4140 0 0 $X=10175 $Y=3980
X40 1 M1M2_C_CDNS_733955477493 $T=10465 12420 0 0 $X=10175 $Y=12260
X41 1 20 9 15 21 inv12f $T=6585 8280 1 0 $X=6405 $Y=3835
X42 1 20 22 23 24 inv15f $T=7525 8280 0 0 $X=7335 $Y=8015
X43 2 20 9 25 26 div_fixed $T=0 8280 0 0 $X=-180 $Y=8015
X44 1 20 9 19 27 28 inv14f $T=9405 8280 1 0 $X=9225 $Y=3835
X45 1 20 9 12 inv11f $T=5775 8280 0 0 $X=5585 $Y=8015
X46 1 20 9 10 inv10f $T=4080 8280 0 0 $X=3900 $Y=8015
X47 1 20 2 8 29 30 inv08f $T=3260 8280 1 0 $X=3080 $Y=3835
X48 1 20 13 18 27 28 inv05f $T=9405 0 0 0 $X=9225 $Y=-265
X49 1 20 4 7 29 30 inv02f $T=3260 0 0 0 $X=3080 $Y=-265
X50 1 20 2 5 31 32 inv07f $T=1630 8280 1 0 $X=1450 $Y=3835
X51 1 20 13 16 33 34 inv04f $T=7900 0 0 0 $X=7720 $Y=-265
X52 1 20 9 17 33 24 34 inv13f $T=7965 8280 1 0 $X=7785 $Y=3835
X53 1 20 2 11 35 inv09f $T=4955 8280 1 0 $X=4765 $Y=3835
X54 1 20 2 3 36 25 37 26 inv06f $T=0 8280 1 0 $X=-180 $Y=3835
X55 1 20 13 14 21 inv03f $T=6270 0 0 0 $X=6090 $Y=-265
X56 1 20 4 6 31 32 inv01f $T=1630 0 0 0 $X=1450 $Y=-265
X57 1 20 2 13 35 preamp1F $T=4640 0 0 0 $X=4460 $Y=-265
X58 1 20 2 4 36 37 preampF $T=0 0 0 0 $X=-180 $Y=-265
.ends pre_therm1
