magic
tech sky130A
timestamp 1704877912
<< pwell >>
rect -142 -129 142 129
<< nmos >>
rect -44 -24 44 24
<< ndiff >>
rect -73 18 -44 24
rect -73 -18 -67 18
rect -50 -18 -44 18
rect -73 -24 -44 -18
rect 44 18 73 24
rect 44 -18 50 18
rect 67 -18 73 18
rect 44 -24 73 -18
<< ndiffc >>
rect -67 -18 -50 18
rect 50 -18 67 18
<< psubdiff >>
rect -124 94 -76 111
rect 76 94 124 111
rect -124 63 -107 94
rect 107 63 124 94
rect -124 -94 -107 -63
rect 107 -94 124 -63
rect -124 -111 -76 -94
rect 76 -111 124 -94
<< psubdiffcont >>
rect -76 94 76 111
rect -124 -63 -107 63
rect 107 -63 124 63
rect -76 -111 76 -94
<< poly >>
rect -44 60 44 68
rect -44 43 -36 60
rect 36 43 44 60
rect -44 24 44 43
rect -44 -43 44 -24
rect -44 -60 -36 -43
rect 36 -60 44 -43
rect -44 -68 44 -60
<< polycont >>
rect -36 43 36 60
rect -36 -60 36 -43
<< locali >>
rect -124 94 -76 111
rect 76 94 124 111
rect -124 63 -107 94
rect 107 63 124 94
rect -44 43 -36 60
rect 36 43 44 60
rect -67 18 -50 26
rect -67 -26 -50 -18
rect 50 18 67 26
rect 50 -26 67 -18
rect -44 -60 -36 -43
rect 36 -60 44 -43
rect -124 -94 -107 -63
rect 107 -94 124 -63
rect -124 -111 -76 -94
rect 76 -111 124 -94
<< viali >>
rect -36 43 36 60
rect -67 -18 -50 18
rect 50 -18 67 18
rect -36 -60 36 -43
<< metal1 >>
rect -42 60 42 63
rect -42 43 -36 60
rect 36 43 42 60
rect -42 40 42 43
rect -70 18 -47 24
rect -70 -18 -67 18
rect -50 -18 -47 18
rect -70 -24 -47 -18
rect 47 18 70 24
rect 47 -18 50 18
rect 67 -18 70 18
rect 47 -24 70 -18
rect -42 -43 42 -40
rect -42 -60 -36 -43
rect 36 -60 42 -43
rect -42 -63 42 -60
<< properties >>
string FIXED_BBOX -115 -102 115 102
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.48 l 0.88 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
