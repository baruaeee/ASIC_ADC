magic
tech sky130A
magscale 1 2
timestamp 1708346635
<< checkpaint >>
rect 0 2427 2628 2676
rect -1313 2241 2668 2427
rect -1313 2152 3125 2241
rect -1313 2133 3864 2152
rect -1313 -925 4261 2133
rect -1313 -2460 2668 -925
<< error_s >>
rect 946 547 999 1069
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use preamp  x2
timestamp 1708346635
transform 1 0 0 0 1 0
box -53 -1200 1408 1167
use sky130_fd_pr__pfet_01v8_LDQF7K  XM0
timestamp 0
transform 1 0 2776 0 1 604
box -225 -269 225 269
use sky130_fd_pr__nfet_01v8_HZA4VB  XM1
timestamp 0
transform 1 0 2208 0 1 640
box -396 -252 396 252
use sky130_fd_pr__pfet_01v8_GEY2B5  XM2
timestamp 0
transform 1 0 1590 0 1 711
box -275 -270 275 270
use sky130_fd_pr__pfet_01v8_KQKFM4  XM3
timestamp 0
transform 1 0 473 0 1 808
box -526 -261 526 261
use sky130_fd_pr__nfet_01v8_5NW376  XM4
timestamp 0
transform 1 0 1157 0 1 955
box -211 -461 211 461
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 V15
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
