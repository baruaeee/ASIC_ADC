magic
tech sky130A
magscale 1 2
timestamp 1706211875
<< error_s >>
rect 200 966 230 1008
rect 286 966 316 1008
rect 155 950 189 958
rect 241 950 275 958
rect 327 950 361 958
rect 155 924 189 932
rect 241 924 275 932
rect 327 924 361 932
rect 155 912 167 924
rect 200 882 230 924
rect 286 882 316 924
rect 349 912 361 924
<< locali >>
rect 405 2419 413 2453
rect 447 2419 455 2453
rect 405 605 455 2419
rect 405 571 413 605
rect 447 571 455 605
<< viali >>
rect 413 2419 447 2453
rect 413 571 447 605
<< metal1 >>
rect 396 2453 464 2464
rect 396 2419 413 2453
rect 447 2419 464 2453
rect 396 2408 464 2419
rect 312 1622 376 1624
rect 312 1570 318 1622
rect 370 1570 376 1622
rect 312 1568 376 1570
rect 312 1454 376 1456
rect 312 1402 318 1454
rect 370 1402 376 1454
rect 312 1400 376 1402
rect 396 605 464 616
rect 396 571 413 605
rect 447 571 464 605
rect 396 560 464 571
<< via1 >>
rect 318 1570 370 1622
rect 318 1402 370 1454
<< metal2 >>
rect 316 1622 372 1628
rect 316 1570 318 1622
rect 370 1570 372 1622
rect 316 1454 372 1570
rect 316 1402 318 1454
rect 370 1402 372 1454
rect 316 1396 372 1402
use NMOS_S_1127905_X1_Y1_1706205215_1706205215  NMOS_S_1127905_X1_Y1_1706205215_1706205215_0
timestamp 1706211875
transform -1 0 516 0 -1 1512
box 52 56 395 1482
use PMOS_S_77083866_X1_Y1_1706205216_1706205215  PMOS_S_77083866_X1_Y1_1706205216_1706205215_0
timestamp 1706211875
transform -1 0 516 0 1 1512
box 0 0 516 1512
<< end >>
