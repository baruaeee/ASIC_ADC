VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
  MACRO oaTaper STRING ;
END PROPERTYDEFINITIONS

MACRO pre_therm
  CLASS CORE ;
  ORIGIN 0 -0.005 ;
  FOREIGN pre_therm 0 0.005 ;
  SIZE 12.57 BY 12.415 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y15
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 9.5 11.005 10.155 11.695 ;
        RECT 9.895 9.025 10.155 11.695 ;
      LAYER met2 ;
        RECT 10.46 11.35 10.96 11.85 ;
        RECT 9.5 11.35 10.96 11.67 ;
      LAYER via ;
        RECT 9.555 11.435 9.705 11.585 ;
    END
  END Y15
  PIN Y14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 11.635 7.3 11.955 7.56 ;
        RECT 11.635 4.84 11.865 7.56 ;
        RECT 11.205 4.84 11.865 5.53 ;
      LAYER met2 ;
        RECT 12.07 7.18 12.57 7.68 ;
        RECT 11.635 7.3 12.57 7.56 ;
      LAYER via ;
        RECT 11.72 7.355 11.87 7.505 ;
    END
  END Y14
  PIN Y13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 9.995 5.46 10.315 5.72 ;
        RECT 10.08 4.815 10.31 7.56 ;
        RECT 9.715 4.815 10.31 5.505 ;
      LAYER met2 ;
        RECT 12.07 5.46 12.57 5.96 ;
        RECT 9.995 5.46 12.57 5.72 ;
      LAYER via ;
        RECT 10.08 5.515 10.23 5.665 ;
    END
  END Y13
  PIN Y12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.46 6.97 8.95 7.66 ;
        RECT 8.69 4.76 8.95 7.66 ;
        RECT 8.325 4.765 8.95 5.455 ;
        RECT 8.63 4.76 8.95 5.455 ;
      LAYER met2 ;
        RECT 12.07 4.64 12.57 5.14 ;
        RECT 8.63 4.76 12.57 5.02 ;
      LAYER via ;
        RECT 8.715 4.815 8.865 4.965 ;
    END
  END Y12
  PIN Y11
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.59 10.98 8.405 11.67 ;
        RECT 8.145 9.025 8.405 11.67 ;
      LAYER met2 ;
        RECT 7.85 10.545 11.18 10.995 ;
        RECT 10.68 9.295 11.18 10.995 ;
        RECT 7.59 11.35 8.11 11.67 ;
        RECT 7.85 10.545 8.11 11.67 ;
      LAYER via ;
        RECT 7.645 11.435 7.795 11.585 ;
    END
  END Y11
  PIN Y10
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.915 11.025 6.615 11.715 ;
        RECT 6.355 8.97 6.615 11.715 ;
        RECT 5.865 8.97 6.615 9.66 ;
      LAYER met2 ;
        RECT 5.915 11.215 6.415 11.715 ;
        RECT 5.915 11.025 6.175 11.715 ;
      LAYER via ;
        RECT 5.97 11.48 6.12 11.63 ;
    END
  END Y10
  PIN Y09
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.64 5.83 7.57 6.09 ;
        RECT 6.64 5.83 6.97 6.46 ;
        RECT 6.71 4.89 6.94 6.46 ;
        RECT 6.675 5.83 6.935 6.78 ;
      LAYER met2 ;
        RECT 4.37 7.38 6.935 7.64 ;
        RECT 6.675 6.46 6.935 7.64 ;
        RECT 3.32 10.675 4.63 10.935 ;
        RECT 4.37 7.38 4.63 10.935 ;
        RECT 3.32 10.555 3.82 11.055 ;
      LAYER via ;
        RECT 6.73 6.545 6.88 6.695 ;
    END
  END Y09
  PIN Y08
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.31 4.765 5.64 6.525 ;
        RECT 5.31 4.765 5.57 6.845 ;
        RECT 4.99 4.765 5.64 5.455 ;
      LAYER met2 ;
        RECT 3.91 6.92 5.57 7.18 ;
        RECT 5.31 6.525 5.57 7.18 ;
        RECT 3.12 9.52 4.17 9.78 ;
        RECT 3.91 6.92 4.17 9.78 ;
        RECT 3.12 9.4 3.62 9.9 ;
      LAYER via ;
        RECT 5.365 6.61 5.515 6.76 ;
    END
  END Y08
  PIN Y07
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.45 6.995 4.15 7.685 ;
        RECT 3.92 4.88 4.15 7.685 ;
        RECT 3.35 4.88 4.15 5.21 ;
      LAYER met2 ;
        RECT 2.435 8.785 3.71 9.105 ;
        RECT 3.45 7.365 3.71 9.105 ;
        RECT 2.435 8.705 2.935 9.205 ;
      LAYER via ;
        RECT 3.505 7.45 3.655 7.6 ;
    END
  END Y07
  PIN Y06
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.92 6.9 2.62 7.59 ;
        RECT 2.39 4.83 2.62 7.59 ;
        RECT 1.975 4.83 2.62 5.16 ;
      LAYER met2 ;
        RECT 1.92 7.33 2.63 7.59 ;
        RECT 2.13 7.09 2.63 7.59 ;
      LAYER via ;
        RECT 2.005 7.385 2.155 7.535 ;
    END
  END Y06
  PIN Y05
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 11.12 2.825 11.89 3.515 ;
        RECT 11.66 0.615 11.89 3.515 ;
        RECT 11.325 0.615 11.89 1.305 ;
      LAYER met2 ;
        RECT 12.07 0.495 12.57 0.995 ;
        RECT 11.57 0.615 12.57 0.875 ;
      LAYER via ;
        RECT 11.655 0.67 11.805 0.82 ;
    END
  END Y05
  PIN Y04
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 9.675 2.615 10.555 3.305 ;
        RECT 10.325 0.725 10.555 3.305 ;
        RECT 9.99 0.725 10.555 1.415 ;
      LAYER met2 ;
        RECT 9.87 0.35 10.37 0.725 ;
        RECT 9.99 0.35 10.25 1.045 ;
      LAYER via ;
        RECT 10.045 0.81 10.195 0.96 ;
    END
  END Y04
  PIN Y03
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.16 3.07 8.945 3.695 ;
        RECT 8.715 0.615 8.945 3.695 ;
        RECT 8.215 0.615 8.945 1.305 ;
        RECT 8.16 3.045 8.39 3.695 ;
      LAYER met2 ;
        RECT 8.215 0.615 8.475 0.935 ;
      LAYER via ;
        RECT 8.27 0.7 8.42 0.85 ;
    END
  END Y03
  PIN Y02
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.05 2.9 5.795 3.59 ;
        RECT 5.565 0.685 5.795 3.59 ;
        RECT 5.065 0.685 5.795 1.015 ;
      LAYER met2 ;
        RECT 4.56 0.685 5.325 1.005 ;
        RECT 4.56 0.685 4.82 1.185 ;
      LAYER via ;
        RECT 5.12 0.77 5.27 0.92 ;
    END
  END Y02
  PIN Y01
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.76 2.86 4.28 3.55 ;
        RECT 4.055 0.525 4.28 3.55 ;
        RECT 3.78 0.525 4.28 1.025 ;
    END
  END Y01
  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
        RECT 10.455 -0.165 11.185 0.165 ;
        RECT 10.23 8.115 10.96 8.445 ;
        RECT 10.455 -0.165 10.785 8.445 ;
      LAYER met1 ;
        RECT 1.18 -0.2 11.965 0.2 ;
        RECT 1.18 8.08 11.965 8.48 ;
        RECT 1.455 8.08 1.685 9.01 ;
      LAYER met2 ;
        RECT 10.48 -0.185 11.16 0.185 ;
        RECT 10.255 8.095 10.935 8.465 ;
      LAYER via ;
        RECT 10.355 8.205 10.505 8.355 ;
        RECT 10.58 -0.075 10.73 0.075 ;
        RECT 10.675 8.205 10.825 8.355 ;
        RECT 10.9 -0.075 11.05 0.075 ;
      LAYER via2 ;
        RECT 10.295 8.18 10.495 8.38 ;
        RECT 10.52 -0.1 10.72 0.1 ;
        RECT 10.695 8.18 10.895 8.38 ;
        RECT 10.92 -0.1 11.12 0.1 ;
    END
  END VSS
  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 11.235 12.255 11.965 12.585 ;
        RECT 11.635 3.975 11.965 12.585 ;
        RECT 11.235 3.975 11.965 4.305 ;
      LAYER met3 ;
        RECT 11.24 3.95 11.96 4.33 ;
        RECT 11.23 3.975 11.96 4.305 ;
        RECT 11.24 12.23 11.96 12.61 ;
        RECT 11.23 12.255 11.96 12.585 ;
      LAYER met1 ;
        RECT 10.585 3.9 11.965 4.38 ;
        RECT 1.055 3.94 11.965 4.34 ;
        RECT 7.765 3.9 10.525 4.34 ;
        RECT 9.08 3.9 10.46 4.38 ;
        RECT 8.945 3.9 10.46 4.345 ;
        RECT 7.45 3.94 8.83 4.38 ;
        RECT 2.81 3.94 7.2 4.38 ;
        RECT 4.44 3.9 5.82 4.38 ;
        RECT 2.81 3.9 4.19 4.38 ;
        RECT 1.055 3.9 2.56 4.38 ;
        RECT 1.055 0.47 1.425 1.52 ;
        RECT 1.055 0.47 1.255 4.38 ;
        RECT 5.26 12.22 11.965 12.62 ;
        RECT 5.26 12.22 6.64 12.66 ;
      LAYER met2 ;
        RECT 11.255 3.955 11.935 4.325 ;
        RECT 11.255 12.235 11.935 12.605 ;
      LAYER via ;
        RECT 11.41 12.345 11.56 12.495 ;
        RECT 11.41 4.065 11.56 4.215 ;
        RECT 11.73 12.345 11.88 12.495 ;
        RECT 11.73 4.065 11.88 4.215 ;
      LAYER via2 ;
        RECT 11.295 12.32 11.495 12.52 ;
        RECT 11.295 4.04 11.495 4.24 ;
        RECT 11.695 12.32 11.895 12.52 ;
        RECT 11.695 4.04 11.895 4.24 ;
      LAYER via3 ;
        RECT 11.3 12.32 11.5 12.52 ;
        RECT 11.3 4.04 11.5 4.24 ;
        RECT 11.7 12.32 11.9 12.52 ;
        RECT 11.7 4.04 11.9 4.24 ;
    END
  END VDD
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.28 0.805 6.835 1.175 ;
        RECT 5.97 6.02 6.34 6.39 ;
        RECT 5.97 5.825 6.23 6.39 ;
        RECT 4.41 6.35 4.78 6.72 ;
        RECT 3.06 5.775 3.43 6.145 ;
        RECT 1.55 5.775 1.92 6.145 ;
        RECT 1.41 1.855 1.78 2.705 ;
        RECT 1.085 10.615 1.525 11.995 ;
        RECT 0.5 10.615 1.525 10.875 ;
        RECT 0.5 10.555 0.76 10.875 ;
      LAYER met2 ;
        RECT 5.525 0.855 6.54 1.175 ;
        RECT 0 5.885 6.23 6.145 ;
        RECT 1.87 5.825 6.23 6.145 ;
        RECT 0.5 2.445 5.785 2.705 ;
        RECT 5.525 0.855 5.785 2.705 ;
        RECT 4.41 5.825 4.67 6.67 ;
        RECT 0.5 2.445 0.76 10.875 ;
        RECT 0 5.765 0.76 6.265 ;
      LAYER via ;
        RECT 0.555 10.64 0.705 10.79 ;
        RECT 1.495 2.5 1.645 2.65 ;
        RECT 1.635 5.94 1.785 6.09 ;
        RECT 3.115 5.91 3.265 6.06 ;
        RECT 4.465 6.435 4.615 6.585 ;
        RECT 6.025 5.91 6.175 6.06 ;
        RECT 6.335 0.94 6.485 1.09 ;
    END
  END IN
  OBS
    LAYER mcon ;
      RECT 11.665 7.28 11.835 7.45 ;
      RECT 11.42 -0.085 11.59 0.085 ;
      RECT 11.42 4.055 11.59 4.225 ;
      RECT 11.42 8.195 11.59 8.365 ;
      RECT 11.355 0.695 11.525 0.865 ;
      RECT 11.355 1.055 11.525 1.225 ;
      RECT 11.235 4.92 11.405 5.09 ;
      RECT 11.235 5.28 11.405 5.45 ;
      RECT 11.15 2.905 11.32 3.075 ;
      RECT 11.15 3.265 11.32 3.435 ;
      RECT 11.02 6.45 11.19 6.62 ;
      RECT 11.01 1.725 11.18 1.895 ;
      RECT 10.96 -0.085 11.13 0.085 ;
      RECT 10.96 4.055 11.13 4.225 ;
      RECT 10.96 8.195 11.13 8.365 ;
      RECT 10.11 7.28 10.28 7.45 ;
      RECT 10.02 0.805 10.19 0.975 ;
      RECT 10.02 1.165 10.19 1.335 ;
      RECT 9.98 8.195 10.15 8.365 ;
      RECT 9.925 9.105 10.095 9.275 ;
      RECT 9.915 -0.085 10.085 0.085 ;
      RECT 9.915 4.055 10.085 4.225 ;
      RECT 9.745 4.895 9.915 5.065 ;
      RECT 9.745 5.255 9.915 5.425 ;
      RECT 9.705 2.695 9.875 2.865 ;
      RECT 9.705 3.055 9.875 3.225 ;
      RECT 9.57 0.945 9.74 1.115 ;
      RECT 9.54 12.335 9.71 12.505 ;
      RECT 9.53 11.085 9.7 11.255 ;
      RECT 9.53 11.445 9.7 11.615 ;
      RECT 9.525 6.405 9.695 6.575 ;
      RECT 9.52 8.195 9.69 8.365 ;
      RECT 9.455 -0.085 9.625 0.085 ;
      RECT 9.455 4.055 9.625 4.225 ;
      RECT 9.32 9.96 9.49 10.13 ;
      RECT 9.08 8.195 9.25 8.365 ;
      RECT 9.08 12.335 9.25 12.505 ;
      RECT 8.645 4.055 8.815 4.225 ;
      RECT 8.6 8.195 8.77 8.365 ;
      RECT 8.49 7.05 8.66 7.22 ;
      RECT 8.49 7.41 8.66 7.58 ;
      RECT 8.355 4.865 8.525 5.035 ;
      RECT 8.355 5.225 8.525 5.395 ;
      RECT 8.285 -0.085 8.455 0.085 ;
      RECT 8.285 4.055 8.455 4.225 ;
      RECT 8.245 0.695 8.415 0.865 ;
      RECT 8.245 1.055 8.415 1.225 ;
      RECT 8.19 3.105 8.36 3.275 ;
      RECT 8.19 3.465 8.36 3.635 ;
      RECT 8.175 9.105 8.345 9.275 ;
      RECT 8.15 8.195 8.32 8.365 ;
      RECT 8.145 6.01 8.315 6.18 ;
      RECT 7.875 1.785 8.045 1.955 ;
      RECT 7.825 -0.085 7.995 0.085 ;
      RECT 7.825 4.055 7.995 4.225 ;
      RECT 7.79 8.195 7.96 8.365 ;
      RECT 7.79 12.335 7.96 12.505 ;
      RECT 7.62 11.06 7.79 11.23 ;
      RECT 7.62 11.42 7.79 11.59 ;
      RECT 7.35 9.96 7.52 10.13 ;
      RECT 7.33 8.195 7.5 8.365 ;
      RECT 7.33 12.335 7.5 12.505 ;
      RECT 7.115 4.055 7.285 4.225 ;
      RECT 6.97 8.195 7.14 8.365 ;
      RECT 6.74 4.97 6.91 5.14 ;
      RECT 6.72 6.26 6.89 6.43 ;
      RECT 6.655 -0.085 6.825 0.085 ;
      RECT 6.655 4.055 6.825 4.225 ;
      RECT 6.545 0.905 6.715 1.075 ;
      RECT 6.51 8.195 6.68 8.365 ;
      RECT 6.46 1.705 6.63 1.875 ;
      RECT 6.46 2.065 6.63 2.235 ;
      RECT 6.195 -0.085 6.365 0.085 ;
      RECT 6.195 4.055 6.365 4.225 ;
      RECT 6.095 8.195 6.265 8.365 ;
      RECT 6.095 12.335 6.265 12.505 ;
      RECT 6.07 6.12 6.24 6.29 ;
      RECT 5.945 11.105 6.115 11.275 ;
      RECT 5.945 11.465 6.115 11.635 ;
      RECT 5.895 9.05 6.065 9.22 ;
      RECT 5.895 9.41 6.065 9.58 ;
      RECT 5.675 10.055 5.845 10.225 ;
      RECT 5.635 8.195 5.805 8.365 ;
      RECT 5.635 12.335 5.805 12.505 ;
      RECT 5.39 6.325 5.56 6.495 ;
      RECT 5.275 -0.085 5.445 0.085 ;
      RECT 5.275 4.055 5.445 4.225 ;
      RECT 5.275 8.195 5.445 8.365 ;
      RECT 5.095 0.765 5.265 0.935 ;
      RECT 5.08 2.98 5.25 3.15 ;
      RECT 5.08 3.34 5.25 3.51 ;
      RECT 5.02 4.845 5.19 5.015 ;
      RECT 5.02 5.205 5.19 5.375 ;
      RECT 4.815 -0.085 4.985 0.085 ;
      RECT 4.815 1.545 4.985 1.715 ;
      RECT 4.815 4.055 4.985 4.225 ;
      RECT 4.815 8.195 4.985 8.365 ;
      RECT 4.51 6.45 4.68 6.62 ;
      RECT 3.81 0.61 3.98 0.78 ;
      RECT 3.79 2.94 3.96 3.11 ;
      RECT 3.79 3.3 3.96 3.47 ;
      RECT 3.645 -0.085 3.815 0.085 ;
      RECT 3.645 4.055 3.815 4.225 ;
      RECT 3.645 8.195 3.815 8.365 ;
      RECT 3.48 7.075 3.65 7.245 ;
      RECT 3.48 7.435 3.65 7.605 ;
      RECT 3.38 4.96 3.55 5.13 ;
      RECT 3.3 1.545 3.47 1.715 ;
      RECT 3.185 -0.085 3.355 0.085 ;
      RECT 3.185 4.055 3.355 4.225 ;
      RECT 3.185 8.195 3.355 8.365 ;
      RECT 3.16 5.875 3.33 6.045 ;
      RECT 2.445 10.885 2.615 11.055 ;
      RECT 2.195 3.485 2.365 3.655 ;
      RECT 2.015 -0.085 2.185 0.085 ;
      RECT 2.015 4.055 2.185 4.225 ;
      RECT 2.015 8.195 2.185 8.365 ;
      RECT 2.005 4.91 2.175 5.08 ;
      RECT 1.95 6.98 2.12 7.15 ;
      RECT 1.95 7.34 2.12 7.51 ;
      RECT 1.705 9.405 1.875 9.575 ;
      RECT 1.705 9.765 1.875 9.935 ;
      RECT 1.665 0.55 1.835 0.72 ;
      RECT 1.665 0.91 1.835 1.08 ;
      RECT 1.665 1.27 1.835 1.44 ;
      RECT 1.65 5.875 1.82 6.045 ;
      RECT 1.555 -0.085 1.725 0.085 ;
      RECT 1.555 4.055 1.725 4.225 ;
      RECT 1.555 8.195 1.725 8.365 ;
      RECT 1.51 2.05 1.68 2.22 ;
      RECT 1.485 8.78 1.655 8.95 ;
      RECT 1.24 10.99 1.41 11.16 ;
      RECT 1.24 11.45 1.41 11.62 ;
      RECT 1.225 0.55 1.395 0.72 ;
      RECT 1.225 0.91 1.395 1.08 ;
      RECT 1.225 1.27 1.395 1.44 ;
    LAYER met1 ;
      RECT 10.91 1.625 11.17 2.005 ;
      RECT 10.91 1.625 11.28 1.995 ;
      RECT 6.435 1.57 6.66 2.47 ;
      RECT 7.775 1.685 8.145 2.325 ;
      RECT 6.43 1.645 6.66 2.295 ;
      RECT 6.43 1.685 8.145 2.005 ;
      RECT 7.25 9.86 7.51 10.275 ;
      RECT 7.25 9.86 7.62 10.23 ;
      RECT 2.365 9.325 2.695 11.085 ;
      RECT 2.365 9.955 5.945 10.325 ;
      RECT 1.675 9.325 2.695 10.015 ;
      RECT 2.135 0.47 2.425 3.685 ;
      RECT 3.2 1.35 3.57 2.2 ;
      RECT 2.135 1.35 3.57 1.67 ;
      RECT 1.635 0.47 2.425 1.52 ;
      RECT 10.92 6.35 11.29 6.72 ;
      RECT 9.47 0.845 9.84 1.215 ;
      RECT 9.425 6.305 9.795 6.675 ;
      RECT 9.22 9.86 9.59 10.23 ;
      RECT 8.045 5.91 8.415 6.28 ;
      RECT 4.715 1.35 5.085 2.2 ;
    LAYER via ;
      RECT 11.005 6.405 11.155 6.555 ;
      RECT 10.965 1.77 11.115 1.92 ;
      RECT 9.525 0.98 9.675 1.13 ;
      RECT 9.48 6.39 9.63 6.54 ;
      RECT 9.275 9.995 9.425 10.145 ;
      RECT 8.1 6.045 8.25 6.195 ;
      RECT 7.94 1.77 8.09 1.92 ;
      RECT 7.305 10.04 7.455 10.19 ;
      RECT 5.74 10.04 5.89 10.19 ;
      RECT 4.77 1.965 4.92 2.115 ;
      RECT 3.365 1.965 3.515 2.115 ;
    LAYER met2 ;
      RECT 5.685 9.955 7.595 10.275 ;
      RECT 7.335 5.96 7.595 10.275 ;
      RECT 5.685 9.955 9.48 10.23 ;
      RECT 9.22 9.91 9.48 10.23 ;
      RECT 9.425 5.96 9.685 6.625 ;
      RECT 9.425 6.35 11.24 6.61 ;
      RECT 7.335 5.96 9.685 6.28 ;
      RECT 7.885 1.685 11.17 2.005 ;
      RECT 9.47 0.895 9.73 2.005 ;
      RECT 3.31 1.88 4.975 2.2 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END pre_therm

END LIBRARY
