magic
tech sky130A
magscale 1 2
timestamp 1706462747
<< error_p >>
rect -29 131 29 137
rect -29 97 -17 131
rect -29 91 29 97
rect -29 -97 29 -91
rect -29 -131 -17 -97
rect -29 -137 29 -131
<< nwell >>
rect -225 -269 225 269
<< pmos >>
rect -29 -50 29 50
<< pdiff >>
rect -87 38 -29 50
rect -87 -38 -75 38
rect -41 -38 -29 38
rect -87 -50 -29 -38
rect 29 38 87 50
rect 29 -38 41 38
rect 75 -38 87 38
rect 29 -50 87 -38
<< pdiffc >>
rect -75 -38 -41 38
rect 41 -38 75 38
<< nsubdiff >>
rect -189 137 -155 199
rect -189 -199 -155 -137
<< nsubdiffcont >>
rect -189 -137 -155 137
<< poly >>
rect -33 131 33 147
rect -33 97 -17 131
rect 17 97 33 131
rect -33 81 33 97
rect -29 50 29 81
rect -29 -81 29 -50
rect -33 -97 33 -81
rect -33 -131 -17 -97
rect 17 -131 33 -97
rect -33 -147 33 -131
<< polycont >>
rect -17 97 17 131
rect -17 -131 17 -97
<< locali >>
rect -189 137 -155 199
rect -33 97 -17 131
rect 17 97 33 131
rect -75 38 -41 54
rect -75 -54 -41 -38
rect 41 38 75 54
rect 41 -54 75 -38
rect -33 -131 -17 -97
rect 17 -131 33 -97
rect -189 -199 -155 -137
<< viali >>
rect -17 97 17 131
rect -75 -38 -41 38
rect 41 -38 75 38
rect -17 -131 17 -97
<< metal1 >>
rect -29 131 29 137
rect -29 97 -17 131
rect 17 97 29 131
rect -29 91 29 97
rect -81 38 -35 50
rect -81 -38 -75 38
rect -41 -38 -35 38
rect -81 -50 -35 -38
rect 35 38 81 50
rect 35 -38 41 38
rect 75 -38 81 38
rect 35 -50 81 -38
rect -29 -97 29 -91
rect -29 -131 -17 -97
rect 17 -131 29 -97
rect -29 -137 29 -131
<< properties >>
string FIXED_BBOX -172 -216 172 216
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 0.285 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
