* NGSPICE file created from th04.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_42G4RD a_n80_n42# a_n148_n216# a_n33_n130# a_22_n42#
X0 a_22_n42# a_n33_n130# a_n80_n42# a_n148_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_n80_n42# a_22_n42# 0.0604f
C1 a_n33_n130# a_22_n42# 0.00866f
C2 a_n33_n130# a_n80_n42# 0.00866f
C3 a_22_n42# a_n148_n216# 0.0698f
C4 a_n80_n42# a_n148_n216# 0.0698f
C5 a_n33_n130# a_n148_n216# 0.321f
.ends

.subckt sky130_fd_pr__pfet_01v8_DDPLQ8 a_n77_n42# w_n215_n261# a_n33_n139# a_19_n42#
+ VSUBS
X0 a_19_n42# a_n33_n139# a_n77_n42# w_n215_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_n33_n139# a_n77_n42# 0.0127f
C1 a_19_n42# w_n215_n261# 0.0399f
C2 a_19_n42# a_n77_n42# 0.0641f
C3 w_n215_n261# a_n77_n42# 0.017f
C4 a_19_n42# a_n33_n139# 0.0127f
C5 w_n215_n261# a_n33_n139# 0.181f
C6 a_19_n42# VSUBS 0.035f
C7 a_n77_n42# VSUBS 0.05f
C8 a_n33_n139# VSUBS 0.149f
C9 w_n215_n261# VSUBS 0.797f
.ends

.subckt sky130_fd_pr__nfet_01v8_VWP3K3 a_n33_n130# a_15_n42# a_n141_182# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n141_182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n42# a_15_n42# 0.0699f
C1 a_n33_n130# a_15_n42# 0.0209f
C2 a_n33_n130# a_n73_n42# 0.0209f
C3 a_15_n42# a_n141_182# 0.0643f
C4 a_n73_n42# a_n141_182# 0.0643f
C5 a_n33_n130# a_n141_182# 0.317f
.ends

.subckt sky130_fd_pr__pfet_01v8_LZD9A4 a_n80_n42# a_22_n42# a_n33_n139# w_n218_n261#
+ VSUBS
X0 a_22_n42# a_n33_n139# a_n80_n42# w_n218_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_n33_n139# a_n80_n42# 0.0084f
C1 a_22_n42# w_n218_n261# 0.0222f
C2 a_22_n42# a_n80_n42# 0.0604f
C3 w_n218_n261# a_n80_n42# 0.0222f
C4 a_22_n42# a_n33_n139# 0.0084f
C5 w_n218_n261# a_n33_n139# 0.185f
C6 a_22_n42# VSUBS 0.0474f
C7 a_n80_n42# VSUBS 0.0474f
C8 a_n33_n139# VSUBS 0.149f
C9 w_n218_n261# VSUBS 0.775f
.ends

.subckt sky130_fd_pr__nfet_01v8_VRD6K3 a_n77_n42# a_n145_n214# a_n33_n130# a_19_n42#
X0 a_19_n42# a_n33_n130# a_n77_n42# a_n145_n214# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_n77_n42# a_19_n42# 0.0641f
C1 a_n33_n130# a_19_n42# 0.0136f
C2 a_n33_n130# a_n77_n42# 0.0136f
C3 a_19_n42# a_n145_n214# 0.0677f
C4 a_n77_n42# a_n145_n214# 0.0677f
C5 a_n33_n130# a_n145_n214# 0.32f
.ends

.subckt th04 Vp V04 Vin Vn
XXM0 m1_892_n998# Vn Vin Vn sky130_fd_pr__nfet_01v8_42G4RD
XXM1 m1_620_n488# Vp Vin m1_892_n998# Vn sky130_fd_pr__pfet_01v8_DDPLQ8
XXM2 Vp m1_620_n488# Vn Vp sky130_fd_pr__nfet_01v8_VWP3K3
XXM3 Vp V04 m1_892_n998# Vp Vn sky130_fd_pr__pfet_01v8_LZD9A4
XXM4 Vn Vn m1_892_n998# V04 sky130_fd_pr__nfet_01v8_VRD6K3
C0 m1_892_n998# V04 0.13f
C1 Vin V04 0.00141f
C2 Vp m1_892_n998# 0.383f
C3 Vp Vin 0.14f
C4 m1_892_n998# Vin 0.463f
C5 m1_620_n488# V04 0.00264f
C6 Vp m1_620_n488# 0.17f
C7 m1_892_n998# m1_620_n488# 0.0117f
C8 m1_620_n488# Vin 0.0346f
C9 Vp V04 0.0462f
C10 Vin Vn 0.726f
C11 m1_892_n998# Vn 0.932f
C12 V04 Vn 0.351f
C13 Vp Vn 2.17f
C14 m1_620_n488# Vn 0.0634f
.ends

