magic
tech sky130A
magscale 1 2
timestamp 1706233216
<< pwell >>
rect -309 -252 309 252
<< nmos >>
rect -113 -42 113 42
<< ndiff >>
rect -171 30 -113 42
rect -171 -30 -159 30
rect -125 -30 -113 30
rect -171 -42 -113 -30
rect 113 30 171 42
rect 113 -30 125 30
rect 159 -30 171 30
rect 113 -42 171 -30
<< ndiffc >>
rect -159 -30 -125 30
rect 125 -30 159 30
<< psubdiff >>
rect -239 -216 -177 -182
rect 177 -216 239 -182
<< psubdiffcont >>
rect -177 -216 177 -182
<< poly >>
rect -113 114 113 130
rect -113 80 -97 114
rect 97 80 113 114
rect -113 42 113 80
rect -113 -80 113 -42
rect -113 -114 -97 -80
rect 97 -114 113 -80
rect -113 -130 113 -114
<< polycont >>
rect -97 80 97 114
rect -97 -114 97 -80
<< locali >>
rect -113 80 -97 114
rect 97 80 113 114
rect -159 30 -125 46
rect -159 -46 -125 -30
rect 125 30 159 46
rect 125 -46 159 -30
rect -113 -114 -97 -80
rect 97 -114 113 -80
rect -239 -216 -177 -182
rect 177 -216 239 -182
<< viali >>
rect -97 80 97 114
rect -159 -30 -125 30
rect 125 -30 159 30
rect -97 -114 97 -80
<< metal1 >>
rect -109 114 109 120
rect -109 80 -97 114
rect 97 80 109 114
rect -109 74 109 80
rect -165 30 -119 42
rect -165 -30 -159 30
rect -125 -30 -119 30
rect -165 -42 -119 -30
rect 119 30 165 42
rect 119 -30 125 30
rect 159 -30 165 30
rect 119 -42 165 -30
rect -109 -80 109 -74
rect -109 -114 -97 -80
rect 97 -114 109 -80
rect -109 -120 109 -114
<< properties >>
string FIXED_BBOX -256 -199 256 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 1.13 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
