//Verilog HDL for "ADC", "TB_single" "functional"


module TB_single ( );

endmodule
