magic
tech sky130A
magscale 1 2
timestamp 1704387395
<< error_p >>
rect -29 118 29 124
rect -29 84 -17 118
rect -29 78 29 84
rect -29 -84 29 -78
rect -29 -118 -17 -84
rect -29 -124 29 -118
<< pwell >>
rect -211 -256 211 256
<< nmos >>
rect -15 -46 15 46
<< ndiff >>
rect -73 34 -15 46
rect -73 -34 -61 34
rect -27 -34 -15 34
rect -73 -46 -15 -34
rect 15 34 73 46
rect 15 -34 27 34
rect 61 -34 73 34
rect 15 -46 73 -34
<< ndiffc >>
rect -61 -34 -27 34
rect 27 -34 61 34
<< psubdiff >>
rect -175 186 -79 220
rect 79 186 175 220
rect -175 124 -141 186
rect 141 124 175 186
rect -175 -186 -141 -124
rect 141 -186 175 -124
rect -175 -220 -79 -186
rect 79 -220 175 -186
<< psubdiffcont >>
rect -79 186 79 220
rect -175 -124 -141 124
rect 141 -124 175 124
rect -79 -220 79 -186
<< poly >>
rect -33 118 33 134
rect -33 84 -17 118
rect 17 84 33 118
rect -33 68 33 84
rect -15 46 15 68
rect -15 -68 15 -46
rect -33 -84 33 -68
rect -33 -118 -17 -84
rect 17 -118 33 -84
rect -33 -134 33 -118
<< polycont >>
rect -17 84 17 118
rect -17 -118 17 -84
<< locali >>
rect -175 186 -79 220
rect 79 186 175 220
rect -175 124 -141 186
rect 141 124 175 186
rect -33 84 -17 118
rect 17 84 33 118
rect -61 34 -27 50
rect -61 -50 -27 -34
rect 27 34 61 50
rect 27 -50 61 -34
rect -33 -118 -17 -84
rect 17 -118 33 -84
rect -175 -186 -141 -124
rect 141 -186 175 -124
rect -175 -220 -79 -186
rect 79 -220 175 -186
<< viali >>
rect -17 84 17 118
rect -61 -34 -27 34
rect 27 -34 61 34
rect -17 -118 17 -84
<< metal1 >>
rect -29 118 29 124
rect -29 84 -17 118
rect 17 84 29 118
rect -29 78 29 84
rect -67 34 -21 46
rect -67 -34 -61 34
rect -27 -34 -21 34
rect -67 -46 -21 -34
rect 21 34 67 46
rect 21 -34 27 34
rect 61 -34 67 34
rect 21 -46 67 -34
rect -29 -84 29 -78
rect -29 -118 -17 -84
rect 17 -118 29 -84
rect -29 -124 29 -118
<< properties >>
string FIXED_BBOX -158 -203 158 203
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.46 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
