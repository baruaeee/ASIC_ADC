magic
tech sky130A
timestamp 1706241174
<< pwell >>
rect -188 -126 188 126
<< nmos >>
rect -90 -21 90 21
<< ndiff >>
rect -119 15 -90 21
rect -119 -15 -113 15
rect -96 -15 -90 15
rect -119 -21 -90 -15
rect 90 15 119 21
rect 90 -15 96 15
rect 113 -15 119 15
rect 90 -21 119 -15
<< ndiffc >>
rect -113 -15 -96 15
rect 96 -15 113 15
<< psubdiff >>
rect -153 -108 -122 -91
rect 122 -108 151 -91
<< psubdiffcont >>
rect -122 -108 122 -91
<< poly >>
rect -90 57 90 65
rect -90 40 -82 57
rect 82 40 90 57
rect -90 21 90 40
rect -90 -40 90 -21
rect -90 -57 -82 -40
rect 82 -57 90 -40
rect -90 -65 90 -57
<< polycont >>
rect -82 40 82 57
rect -82 -57 82 -40
<< locali >>
rect -90 40 -82 57
rect 82 40 90 57
rect -113 15 -96 23
rect -113 -23 -96 -15
rect 96 15 113 23
rect 96 -23 113 -15
rect -90 -57 -82 -40
rect 82 -57 90 -40
rect -153 -108 -122 -91
rect 122 -108 151 -91
<< viali >>
rect -82 40 82 57
rect -113 -15 -96 15
rect 96 -15 113 15
rect -82 -57 82 -40
<< metal1 >>
rect -88 57 88 60
rect -88 40 -82 57
rect 82 40 88 57
rect -88 37 88 40
rect -116 15 -93 21
rect -116 -15 -113 15
rect -96 -15 -93 15
rect -116 -21 -93 -15
rect 93 15 116 21
rect 93 -15 96 15
rect 113 -15 116 15
rect 93 -21 116 -15
rect -88 -40 88 -37
rect -88 -57 -82 -40
rect 82 -57 88 -40
rect -88 -60 88 -57
<< properties >>
string FIXED_BBOX -161 -99 161 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 1.8 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
