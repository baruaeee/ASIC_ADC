magic
tech sky130A
magscale 1 2
timestamp 1705440736
<< locali >>
rect 672 250 826 324
rect 588 66 698 102
rect 588 -778 624 66
rect 1058 -643 1128 -558
rect 588 -814 710 -778
<< viali >>
rect 1058 -679 1128 -643
<< metal1 >>
rect 976 622 1176 790
rect 718 586 1202 622
rect 718 322 754 586
rect 828 374 896 430
rect 1166 338 1202 586
rect 1260 370 1322 432
rect 718 286 822 322
rect 718 284 782 286
rect 786 284 822 286
rect 718 248 822 284
rect 904 252 984 330
rect 934 226 984 252
rect 1166 282 1260 338
rect 1166 246 1266 282
rect 1320 256 1414 332
rect 1356 228 1414 256
rect 572 164 898 200
rect 572 -328 608 164
rect 948 -4 984 226
rect 1276 -4 1312 212
rect 394 -458 608 -328
rect 718 -40 1312 -4
rect 1378 42 1414 228
rect 718 -340 754 -40
rect 812 -304 882 -250
rect 1242 -304 1278 -40
rect 1378 -158 1590 42
rect 718 -376 824 -340
rect 718 -382 786 -376
rect 788 -382 824 -376
rect 718 -418 824 -382
rect 878 -414 958 -336
rect 906 -424 958 -414
rect 394 -494 882 -458
rect 394 -528 594 -494
rect 774 -978 810 -922
rect 922 -926 958 -424
rect 1146 -418 1236 -336
rect 1378 -354 1414 -158
rect 1292 -416 1414 -354
rect 1146 -442 1206 -418
rect 1146 -612 1182 -442
rect 1234 -514 1296 -452
rect 1126 -637 1182 -612
rect 1046 -643 1182 -637
rect 1046 -679 1058 -643
rect 1128 -646 1182 -643
rect 1128 -679 1272 -646
rect 1046 -682 1272 -679
rect 1046 -685 1140 -682
rect 1102 -978 1138 -924
rect 774 -1014 1138 -978
rect 774 -1016 980 -1014
rect 944 -1116 980 -1016
rect 1236 -1116 1272 -682
rect 1344 -1116 1544 -952
rect 944 -1152 1544 -1116
use sky130_fd_pr__pfet_01v8_XGS3BL  XM0
timestamp 1704310947
transform 0 -1 957 1 0 -953
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_L7T3GD  XM1
timestamp 1704336338
transform 1 0 849 0 1 -378
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_QPDSQG  XM2
timestamp 1704336338
transform 1 0 863 0 1 293
box -225 -261 225 261
use sky130_fd_pr__pfet_01v8_M479BZ  XM3
timestamp 1704336338
transform 1 0 1293 0 1 293
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_L7T3GD  XM4
timestamp 1704336338
transform 1 0 1265 0 1 -378
box -211 -252 211 252
<< labels >>
flabel metal1 394 -528 594 -328 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 976 590 1176 790 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 1390 -158 1590 42 0 FreeSans 256 0 0 0 V10
port 1 nsew
flabel metal1 1344 -1152 1544 -952 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
