magic
tech sky130A
magscale 1 2
timestamp 1706529083
<< nwell >>
rect 2878 -1714 3806 -1488
rect 3808 -1708 4222 -1544
rect 4646 -1708 4894 -1528
rect 3808 -1714 4894 -1708
rect 2878 -1754 4894 -1714
rect 2878 -1756 3866 -1754
rect 2878 -1768 3824 -1756
rect 2878 -1840 3806 -1768
rect 4214 -1796 4894 -1754
rect 4214 -1912 4890 -1796
rect 2952 -4424 3304 -4242
<< pwell >>
rect 4210 -758 4260 -696
<< locali >>
rect 3673 -2476 3770 -2438
<< viali >>
rect 3639 -2476 3673 -2438
rect 3554 -3395 3588 -3361
<< metal1 >>
rect 3103 -17 3155 -11
rect 2398 -38 2450 -32
rect 2319 -81 2398 -47
rect 2319 -511 2353 -81
rect 2398 -96 2450 -90
rect 2964 -63 3103 -26
rect 2964 -511 2998 -63
rect 3103 -75 3155 -69
rect 1766 -545 4843 -511
rect 3028 -598 3072 -545
rect 5118 -559 5218 -528
rect 4957 -593 5443 -559
rect 1538 -1162 1638 -1062
rect 1585 -1327 1619 -1162
rect 2945 -1842 2979 -1651
rect 3028 -1714 3065 -598
rect 5118 -628 5218 -593
rect 4156 -698 4256 -660
rect 4156 -702 4308 -698
rect 4156 -754 4209 -702
rect 4261 -754 4308 -702
rect 4156 -758 4308 -754
rect 4156 -760 4256 -758
rect 5409 -769 5443 -593
rect 5144 -1135 5244 -1092
rect 4943 -1169 5244 -1135
rect 5144 -1192 5244 -1169
rect 4054 -1270 4106 -1264
rect 4054 -1328 4106 -1322
rect 3138 -1355 3190 -1349
rect 3138 -1413 3190 -1407
rect 5340 -1354 5417 -1295
rect 5340 -1391 5420 -1354
rect 5340 -1392 5404 -1391
rect 3022 -1720 3074 -1714
rect 3022 -1778 3074 -1772
rect 1747 -2502 1781 -2325
rect 1700 -2602 1800 -2502
rect 1786 -2956 1823 -2879
rect 1774 -3008 1780 -2956
rect 1832 -3008 1838 -2956
rect 2151 -3012 2203 -3006
rect 2151 -3070 2203 -3064
rect 3331 -3095 3365 -1445
rect 3581 -1591 3615 -1545
rect 4822 -1604 4834 -1598
rect 4814 -1636 4862 -1604
rect 4786 -1669 4886 -1636
rect 5340 -1669 5377 -1392
rect 4217 -1703 5377 -1669
rect 4786 -1736 4886 -1703
rect 4151 -1992 4157 -1940
rect 4209 -1992 4215 -1940
rect 3620 -2324 3626 -2272
rect 3678 -2276 3684 -2272
rect 3678 -2315 3878 -2276
rect 3678 -2324 3684 -2315
rect 5064 -2360 5164 -2324
rect 4956 -2416 5286 -2360
rect 5064 -2424 5164 -2416
rect 3538 -2438 3590 -2432
rect 3633 -2438 3679 -2426
rect 3633 -2447 3639 -2438
rect 3590 -2476 3639 -2447
rect 3673 -2476 3679 -2438
rect 3590 -2481 3679 -2476
rect 3633 -2488 3679 -2481
rect 3538 -2496 3590 -2490
rect 5230 -2772 5286 -2416
rect 5315 -3005 5407 -2971
rect 5315 -3025 5349 -3005
rect 4624 -3059 5349 -3025
rect 3614 -3072 3786 -3059
rect 3331 -3129 3601 -3095
rect 3614 -3116 3788 -3072
rect 3627 -3122 3788 -3116
rect 2145 -3304 2151 -3252
rect 2203 -3304 2209 -3252
rect 3331 -3549 3365 -3129
rect 3521 -3270 3555 -3249
rect 3486 -3322 3492 -3270
rect 3544 -3322 3555 -3270
rect 3501 -3333 3555 -3322
rect 3501 -3343 3595 -3333
rect 3501 -3361 3597 -3343
rect 3501 -3395 3554 -3361
rect 3588 -3395 3597 -3361
rect 3501 -3403 3597 -3395
rect 3548 -3407 3594 -3403
rect 3159 -3583 3365 -3549
rect 2634 -3649 2734 -3600
rect 2634 -3683 2853 -3649
rect 2634 -3700 2734 -3683
rect 3159 -3955 3193 -3583
rect 4920 -3600 5020 -3500
rect 3269 -3673 3786 -3636
rect 3269 -3739 3306 -3673
rect 4931 -3687 4965 -3600
rect 4781 -3721 4965 -3687
rect 3257 -3791 3263 -3739
rect 3315 -3791 3321 -3739
rect 3015 -3989 3193 -3955
rect 3015 -4400 3049 -3989
rect 3082 -4348 3088 -4296
rect 3140 -4305 3146 -4296
rect 3140 -4339 3255 -4305
rect 3140 -4348 3146 -4339
rect 3372 -4370 3424 -4364
rect 3015 -4487 3059 -4400
rect 3372 -4428 3424 -4422
rect 2933 -5452 2939 -5400
rect 2991 -5452 2997 -5400
rect 3025 -5817 3059 -4487
rect 4112 -5022 4212 -4922
rect 3874 -5508 3911 -5490
rect 3240 -5537 3292 -5531
rect 3863 -5545 3911 -5508
rect 3292 -5582 3954 -5545
rect 3824 -5586 3911 -5582
rect 3240 -5595 3292 -5589
rect 3025 -5851 3283 -5817
rect 3080 -6454 3086 -6402
rect 3141 -6454 3147 -6402
rect 4740 -6440 4840 -6340
rect 3080 -6455 3209 -6454
rect 3080 -6456 3232 -6455
rect 3080 -6464 3401 -6456
rect 3079 -6498 3401 -6464
rect 3202 -6499 3401 -6498
<< via1 >>
rect 2398 -90 2450 -38
rect 3103 -69 3155 -17
rect 4209 -754 4261 -702
rect 4054 -1322 4106 -1270
rect 3138 -1407 3190 -1355
rect 3022 -1772 3074 -1720
rect 1780 -3008 1832 -2956
rect 2151 -3064 2203 -3012
rect 4157 -1992 4209 -1940
rect 3626 -2324 3678 -2272
rect 3538 -2490 3590 -2438
rect 2151 -3304 2203 -3252
rect 3492 -3322 3544 -3270
rect 3263 -3791 3315 -3739
rect 3088 -4348 3140 -4296
rect 3372 -4422 3424 -4370
rect 2939 -5452 2991 -5400
rect 3240 -5589 3292 -5537
rect 3086 -6454 3141 -6402
<< metal2 >>
rect 3190 -16 3246 -7
rect 2434 -36 2490 -27
rect 2392 -90 2398 -38
rect 3097 -69 3103 -17
rect 3155 -21 3161 -17
rect 3155 -66 3190 -21
rect 3155 -69 3161 -66
rect 3190 -81 3246 -72
rect 2434 -101 2490 -92
rect 4209 -702 4261 -696
rect 4209 -760 4218 -754
rect 4252 -760 4261 -754
rect 4048 -1322 4054 -1270
rect 4106 -1279 4112 -1270
rect 4106 -1313 4252 -1279
rect 4106 -1322 4112 -1313
rect 3100 -1355 3198 -1354
rect 3100 -1364 3138 -1355
rect 2688 -1407 3138 -1364
rect 3190 -1407 3198 -1355
rect 2688 -1408 3198 -1407
rect 3016 -1772 3022 -1720
rect 3074 -1729 3080 -1720
rect 3074 -1763 3669 -1729
rect 3074 -1772 3080 -1763
rect 3635 -2266 3669 -1763
rect 4055 -1743 4089 -1322
rect 4055 -1777 4200 -1743
rect 4166 -1934 4200 -1777
rect 4157 -1940 4209 -1934
rect 4157 -1998 4209 -1992
rect 3626 -2272 3678 -2266
rect 3626 -2330 3678 -2324
rect 3626 -2331 3663 -2330
rect 3481 -2492 3490 -2436
rect 3546 -2438 3555 -2436
rect 3590 -2490 3596 -2438
rect 3546 -2492 3555 -2490
rect 1780 -2956 1832 -2950
rect 1780 -3014 1832 -3008
rect 3405 -2961 3766 -2927
rect 1783 -3043 1828 -3014
rect 1768 -3099 1777 -3043
rect 1833 -3099 1842 -3043
rect 2145 -3064 2151 -3012
rect 2203 -3064 2209 -3012
rect 3405 -3023 3439 -2961
rect 2795 -3057 3439 -3023
rect 2160 -3246 2194 -3064
rect 2151 -3252 2203 -3246
rect 2151 -3310 2203 -3304
rect 3263 -3739 3315 -3733
rect 3263 -3797 3315 -3791
rect 3266 -3826 3311 -3797
rect 3251 -3882 3260 -3826
rect 3316 -3882 3325 -3826
rect 3088 -4296 3140 -4290
rect 3077 -4376 3086 -4320
rect 3142 -4376 3151 -4320
rect 3405 -4370 3439 -3057
rect 3481 -3288 3490 -3232
rect 3546 -3288 3555 -3232
rect 3492 -3328 3544 -3322
rect 3366 -4422 3372 -4370
rect 3424 -4413 3439 -4370
rect 3424 -4422 3430 -4413
rect 2929 -5365 2938 -5309
rect 2994 -5365 3003 -5309
rect 2943 -5394 2988 -5365
rect 2939 -5400 2991 -5394
rect 2939 -5458 2991 -5452
rect 2944 -5545 2981 -5458
rect 3234 -5545 3240 -5537
rect 2944 -5582 3240 -5545
rect 3234 -5589 3240 -5582
rect 3292 -5589 3298 -5537
rect 3076 -6411 3085 -6355
rect 3141 -6411 3150 -6355
rect 3086 -6460 3141 -6454
<< via2 >>
rect 2434 -38 2490 -36
rect 2434 -90 2450 -38
rect 2450 -90 2490 -38
rect 3190 -72 3246 -16
rect 2434 -92 2490 -90
rect 3490 -2438 3546 -2436
rect 3490 -2490 3538 -2438
rect 3538 -2490 3546 -2438
rect 3490 -2492 3546 -2490
rect 1777 -3099 1833 -3043
rect 3260 -3882 3316 -3826
rect 3086 -4348 3088 -4320
rect 3088 -4348 3140 -4320
rect 3140 -4348 3142 -4320
rect 3086 -4376 3142 -4348
rect 3490 -3270 3546 -3232
rect 3490 -3288 3492 -3270
rect 3492 -3288 3544 -3270
rect 3544 -3288 3546 -3270
rect 2938 -5365 2994 -5309
rect 3085 -6402 3141 -6355
rect 3085 -6411 3086 -6402
rect 3086 -6411 3141 -6402
<< metal3 >>
rect 3100 -10 3164 -6
rect 3100 -11 3228 -10
rect 3100 -12 3251 -11
rect 2429 -34 2495 -31
rect 2429 -36 2749 -34
rect 2429 -92 2434 -36
rect 2490 -92 2749 -36
rect 3164 -16 3251 -12
rect 3164 -72 3190 -16
rect 3246 -72 3251 -16
rect 3164 -76 3251 -72
rect 3100 -77 3251 -76
rect 3100 -80 3224 -77
rect 3100 -82 3164 -80
rect 2429 -94 2749 -92
rect 2429 -97 2495 -94
rect 3485 -2436 3551 -2431
rect 3485 -2492 3490 -2436
rect 3546 -2492 3551 -2436
rect 3485 -2497 3551 -2492
rect 1767 -3017 1773 -2953
rect 1837 -3017 1843 -2953
rect 1769 -3043 1839 -3017
rect 1769 -3077 1777 -3043
rect 1772 -3099 1777 -3077
rect 1833 -3081 1839 -3043
rect 1833 -3099 1838 -3081
rect 1772 -3104 1838 -3099
rect 3488 -3227 3548 -2497
rect 3485 -3232 3551 -3227
rect 3485 -3288 3490 -3232
rect 3546 -3288 3551 -3232
rect 3485 -3293 3551 -3288
rect 3250 -3800 3256 -3736
rect 3320 -3800 3326 -3736
rect 3252 -3826 3322 -3800
rect 3252 -3860 3260 -3826
rect 3255 -3882 3260 -3860
rect 3316 -3864 3322 -3826
rect 3316 -3882 3321 -3864
rect 3255 -3887 3321 -3882
rect 3081 -4320 3147 -4315
rect 3081 -4376 3086 -4320
rect 3142 -4376 3147 -4320
rect 3081 -4381 3147 -4376
rect 2933 -5309 2999 -5304
rect 2933 -5327 2938 -5309
rect 2932 -5365 2938 -5327
rect 2994 -5331 2999 -5309
rect 2994 -5365 3002 -5331
rect 2932 -5391 3002 -5365
rect 2928 -5455 2934 -5391
rect 2998 -5455 3004 -5391
rect 3084 -6253 3144 -4381
rect 3083 -6350 3144 -6253
rect 3080 -6355 3146 -6350
rect 3080 -6411 3085 -6355
rect 3141 -6411 3146 -6355
rect 3080 -6416 3146 -6411
<< via3 >>
rect 3100 -76 3164 -12
rect 1773 -3017 1837 -2953
rect 3256 -3800 3320 -3736
rect 2934 -5455 2998 -5391
<< metal4 >>
rect 3099 -12 3165 -11
rect 3099 -14 3100 -12
rect 3060 -74 3100 -14
rect 3099 -76 3100 -74
rect 3164 -14 3165 -12
rect 3164 -74 3274 -14
rect 3164 -76 3165 -74
rect 3099 -77 3165 -76
rect 1775 -2952 1835 -2913
rect 1772 -2953 1838 -2952
rect 1772 -3017 1773 -2953
rect 1837 -3017 1838 -2953
rect 1772 -3018 1838 -3017
rect 1775 -3100 1835 -3018
rect 1774 -3160 3318 -3100
rect 3258 -3735 3318 -3160
rect 3255 -3736 3321 -3735
rect 3255 -3800 3256 -3736
rect 3320 -3800 3321 -3736
rect 3255 -3801 3321 -3800
rect 3258 -4106 3318 -3801
rect 2936 -4166 3318 -4106
rect 2936 -5390 2996 -4166
rect 2933 -5391 2999 -5390
rect 2933 -5455 2934 -5391
rect 2998 -5455 2999 -5391
rect 2933 -5456 2999 -5455
rect 2936 -5495 2996 -5456
use preamp  preamp_0
timestamp 1706402911
transform -1 0 4522 0 -1 -374
box 394 136 1494 1340
use th01  th01_0
timestamp 1706270854
transform 1 0 2870 0 -1 -6940
box 316 -1456 1968 6
use th09  th09_0
timestamp 1706479318
transform 1 0 1406 0 -1 -3900
box 368 -754 1692 524
use th10  th10_0
timestamp 1706270854
transform 1 0 3944 0 -1 -1282
box 270 -794 1168 452
use th11  th11_0
timestamp 1706241174
transform 1 0 2720 0 1 -4710
box 466 -880 1630 468
use th12  th12_0
timestamp 1706270854
transform 1 0 3422 0 1 -1986
box 278 -1078 1572 236
use th13  th13_0
timestamp 1706474503
transform -1 0 3736 0 1 -2482
box 438 -680 2042 646
use th14  th14_0
timestamp 1706473616
transform 1 0 2994 0 -1 -3516
box 524 -532 1974 728
use th15  th15_0
timestamp 1706464016
transform -1 0 3478 0 -1 -1688
box 482 -1164 1936 152
<< labels >>
flabel metal1 5118 -628 5218 -528 0 FreeSans 256 180 0 0 Vn
port 17 nsew
flabel metal1 4156 -760 4256 -660 0 FreeSans 256 0 0 0 Vin
port 0 nsew
flabel metal1 4786 -1736 4886 -1636 0 FreeSans 256 0 0 0 Vp
port 1 nsew
flabel metal1 5144 -1192 5244 -1092 0 FreeSans 256 180 0 0 V10
port 10 nsew
flabel metal1 5064 -2424 5164 -2324 0 FreeSans 256 180 0 0 V12
port 12 nsew
flabel metal1 4920 -3600 5020 -3500 0 FreeSans 256 180 0 0 V14
port 14 nsew
flabel metal1 1538 -1162 1638 -1062 0 FreeSans 256 180 0 0 V15
port 15 nsew
flabel metal1 4112 -5022 4212 -4922 0 FreeSans 256 0 0 0 V11
port 11 nsew
flabel metal1 4740 -6440 4840 -6340 0 FreeSans 256 0 0 0 V01
port 2 nsew
flabel metal1 1700 -2602 1800 -2502 0 FreeSans 256 180 0 0 V13
port 13 nsew
flabel metal1 2634 -3700 2734 -3600 0 FreeSans 256 0 0 0 V09
port 9 nsew
<< end >>
