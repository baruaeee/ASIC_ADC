magic
tech sky130A
magscale 1 2
timestamp 1706211875
<< nwell >>
rect 0 0 516 1512
<< pmos >>
rect 200 525 230 609
rect 286 525 316 609
<< pdiff >>
rect 147 575 200 609
rect 147 541 155 575
rect 189 541 200 575
rect 147 525 200 541
rect 230 575 286 609
rect 230 541 241 575
rect 275 541 286 575
rect 230 525 286 541
rect 316 575 369 609
rect 316 541 327 575
rect 361 541 369 575
rect 316 525 369 541
<< pdiffc >>
rect 155 541 189 575
rect 241 541 275 575
rect 327 541 361 575
<< nsubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
<< nsubdiffcont >>
rect 241 1327 275 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 609 230 897
rect 286 609 316 897
rect 200 252 230 525
rect 286 252 316 525
<< polycont >>
rect 241 907 275 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 147 575 197 773
rect 147 541 155 575
rect 189 541 197 575
rect 147 185 197 541
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 575 283 773
rect 233 541 241 575
rect 275 541 283 575
rect 233 101 283 541
rect 233 67 241 101
rect 275 67 283 101
rect 319 575 369 773
rect 319 541 327 575
rect 361 541 369 575
rect 319 185 369 541
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
<< viali >>
rect 241 1327 275 1361
rect 241 907 275 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
<< metal1 >>
rect 52 1361 292 1372
rect 52 1327 241 1361
rect 275 1327 292 1361
rect 52 1316 292 1327
rect 52 941 292 952
rect 52 907 241 941
rect 275 907 292 941
rect 52 896 292 907
rect 138 185 378 196
rect 138 151 155 185
rect 189 151 327 185
rect 361 151 378 185
rect 138 140 378 151
rect 52 101 292 112
rect 52 67 241 101
rect 275 67 292 101
rect 52 56 292 67
<< end >>
