magic
tech sky130A
timestamp 1706239161
<< pwell >>
rect -121 -126 121 126
<< nmos >>
rect -23 -21 23 21
<< ndiff >>
rect -52 15 -23 21
rect -52 -15 -46 15
rect -29 -15 -23 15
rect -52 -21 -23 -15
rect 23 15 52 21
rect 23 -15 29 15
rect 46 -15 52 15
rect 23 -21 52 -15
<< ndiffc >>
rect -46 -15 -29 15
rect 29 -15 46 15
<< psubdiff >>
rect -103 60 -86 91
rect -103 -91 -86 -60
<< psubdiffcont >>
rect -103 -60 -86 60
<< poly >>
rect -23 57 23 65
rect -23 40 -15 57
rect 15 40 23 57
rect -23 21 23 40
rect -23 -40 23 -21
rect -23 -57 -15 -40
rect 15 -57 23 -40
rect -23 -65 23 -57
<< polycont >>
rect -15 40 15 57
rect -15 -57 15 -40
<< locali >>
rect -103 60 -86 91
rect -23 40 -15 57
rect 15 40 23 57
rect -46 15 -29 23
rect -46 -23 -29 -15
rect 29 15 46 23
rect 29 -23 46 -15
rect -23 -57 -15 -40
rect 15 -57 23 -40
rect -103 -91 -86 -60
<< viali >>
rect -15 40 15 57
rect -46 -15 -29 15
rect 29 -15 46 15
rect -15 -57 15 -40
<< metal1 >>
rect -21 57 21 60
rect -21 40 -15 57
rect 15 40 21 57
rect -21 37 21 40
rect -49 15 -26 21
rect -49 -15 -46 15
rect -29 -15 -26 15
rect -49 -21 -26 -15
rect 26 15 49 21
rect 26 -15 29 15
rect 46 -15 49 15
rect 26 -21 49 -15
rect -21 -40 21 -37
rect -21 -57 -15 -40
rect 15 -57 21 -40
rect -21 -60 21 -57
<< properties >>
string FIXED_BBOX -94 -99 94 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.46 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
