magic
tech sky130A
magscale 1 2
timestamp 1706216322
<< nwell >>
rect -332 -263 332 263
<< pmos >>
rect -136 -44 136 44
<< pdiff >>
rect -194 32 -136 44
rect -194 -32 -182 32
rect -148 -32 -136 32
rect -194 -44 -136 -32
rect 136 32 194 44
rect 136 -32 148 32
rect 182 -32 194 32
rect 136 -44 194 -32
<< pdiffc >>
rect -182 -32 -148 32
rect 148 -32 182 32
<< nsubdiff >>
rect -262 193 -200 227
rect 200 193 262 227
<< nsubdiffcont >>
rect -200 193 200 227
<< poly >>
rect -136 125 136 141
rect -136 91 -120 125
rect 120 91 136 125
rect -136 44 136 91
rect -136 -91 136 -44
rect -136 -125 -120 -91
rect 120 -125 136 -91
rect -136 -141 136 -125
<< polycont >>
rect -120 91 120 125
rect -120 -125 120 -91
<< locali >>
rect -262 193 -200 227
rect 200 193 262 227
rect -136 91 -120 125
rect 120 91 136 125
rect -182 32 -148 48
rect -182 -48 -148 -32
rect 148 32 182 48
rect 148 -48 182 -32
rect -136 -125 -120 -91
rect 120 -125 136 -91
<< viali >>
rect -120 91 120 125
rect -182 -32 -148 32
rect 148 -32 182 32
rect -120 -125 120 -91
<< metal1 >>
rect -132 125 132 131
rect -132 91 -120 125
rect 120 91 132 125
rect -132 85 132 91
rect -188 32 -142 44
rect -188 -32 -182 32
rect -148 -32 -142 32
rect -188 -44 -142 -32
rect 142 32 188 44
rect 142 -32 148 32
rect 182 -32 188 32
rect 142 -44 188 -32
rect -132 -91 132 -85
rect -132 -125 -120 -91
rect 120 -125 132 -91
rect -132 -131 132 -125
<< properties >>
string FIXED_BBOX -279 -210 279 210
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.44 l 1.36 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
