magic
tech sky130A
magscale 1 2
timestamp 1704730646
<< error_p >>
rect -29 172 29 178
rect -29 138 -17 172
rect -29 132 29 138
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect -29 -178 29 -172
<< pwell >>
rect -226 -310 226 310
<< nmos >>
rect -30 -100 30 100
<< ndiff >>
rect -88 88 -30 100
rect -88 -88 -76 88
rect -42 -88 -30 88
rect -88 -100 -30 -88
rect 30 88 88 100
rect 30 -88 42 88
rect 76 -88 88 88
rect 30 -100 88 -88
<< ndiffc >>
rect -76 -88 -42 88
rect 42 -88 76 88
<< psubdiff >>
rect -190 240 -94 274
rect 94 240 190 274
rect -190 178 -156 240
rect 156 178 190 240
rect -190 -240 -156 -178
rect 156 -240 190 -178
rect -190 -274 -94 -240
rect 94 -274 190 -240
<< psubdiffcont >>
rect -94 240 94 274
rect -190 -178 -156 178
rect 156 -178 190 178
rect -94 -274 94 -240
<< poly >>
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -33 122 33 138
rect -30 100 30 122
rect -30 -122 30 -100
rect -33 -138 33 -122
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -188 33 -172
<< polycont >>
rect -17 138 17 172
rect -17 -172 17 -138
<< locali >>
rect -190 240 -94 274
rect 94 240 190 274
rect -190 178 -156 240
rect 156 178 190 240
rect -33 138 -17 172
rect 17 138 33 172
rect -76 88 -42 104
rect -76 -104 -42 -88
rect 42 88 76 104
rect 42 -104 76 -88
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -190 -240 -156 -178
rect 156 -240 190 -178
rect -190 -274 -94 -240
rect 94 -274 190 -240
<< viali >>
rect -17 138 17 172
rect -76 -88 -42 88
rect 42 -88 76 88
rect -17 -172 17 -138
<< metal1 >>
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect -82 88 -36 100
rect -82 -88 -76 88
rect -42 -88 -36 88
rect -82 -100 -36 -88
rect 36 88 82 100
rect 36 -88 42 88
rect 76 -88 82 88
rect 36 -100 82 -88
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect 17 -172 29 -138
rect -29 -178 29 -172
<< properties >>
string FIXED_BBOX -173 -257 173 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
