magic
tech sky130A
magscale 1 2
timestamp 1706233216
<< error_p >>
rect -29 148 29 154
rect -29 114 -17 148
rect -29 108 29 114
rect -29 -114 29 -108
rect -29 -148 -17 -114
rect -29 -154 29 -148
<< nwell >>
rect -212 -286 212 286
<< pmos >>
rect -16 -67 16 67
<< pdiff >>
rect -74 55 -16 67
rect -74 -55 -62 55
rect -28 -55 -16 55
rect -74 -67 -16 -55
rect 16 55 74 67
rect 16 -55 28 55
rect 62 -55 74 55
rect 16 -67 74 -55
<< pdiffc >>
rect -62 -55 -28 55
rect 28 -55 62 55
<< nsubdiff >>
rect 142 154 176 216
rect 142 -216 176 -154
<< nsubdiffcont >>
rect 142 -154 176 154
<< poly >>
rect -33 148 33 164
rect -33 114 -17 148
rect 17 114 33 148
rect -33 98 33 114
rect -16 67 16 98
rect -16 -98 16 -67
rect -33 -114 33 -98
rect -33 -148 -17 -114
rect 17 -148 33 -114
rect -33 -164 33 -148
<< polycont >>
rect -17 114 17 148
rect -17 -148 17 -114
<< locali >>
rect 142 154 176 216
rect -33 114 -17 148
rect 17 114 33 148
rect -62 55 -28 71
rect -62 -71 -28 -55
rect 28 55 62 71
rect 28 -71 62 -55
rect -33 -148 -17 -114
rect 17 -148 33 -114
rect 142 -216 176 -154
<< viali >>
rect -17 114 17 148
rect -62 -55 -28 55
rect 28 -55 62 55
rect -17 -148 17 -114
<< metal1 >>
rect -29 148 29 154
rect -29 114 -17 148
rect 17 114 29 148
rect -29 108 29 114
rect -68 55 -22 67
rect -68 -55 -62 55
rect -28 -55 -22 55
rect -68 -67 -22 -55
rect 22 55 68 67
rect 22 -55 28 55
rect 62 -55 68 55
rect 22 -67 68 -55
rect -29 -114 29 -108
rect -29 -148 -17 -114
rect 17 -148 29 -114
rect -29 -154 29 -148
<< properties >>
string FIXED_BBOX -159 -233 159 233
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.668 l 0.16 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
