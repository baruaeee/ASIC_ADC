magic
tech sky130A
magscale 1 2
timestamp 1702941826
<< checkpaint >>
rect -944 2205 6968 2258
rect 9734 2205 12686 2286
rect -944 2117 12686 2205
rect -944 2064 18025 2117
rect 20791 2064 23733 6909
rect -944 -766 23733 2064
rect 4395 -819 23733 -766
rect 9734 -872 23733 -819
rect 10113 -925 23733 -872
rect 15452 -978 23733 -925
rect 20791 -1031 23733 -978
<< error_s >>
rect 299 998 333 1016
rect 299 962 369 998
rect 316 928 387 962
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 928
rect 316 547 369 583
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_KGSDF3  XM1
timestamp 0
transform 1 0 158 0 1 3266
box -211 -2719 211 2719
use sky130_fd_pr__pfet_01v8_SKYSXJ  XM2
timestamp 0
transform 1 0 11210 0 1 707
box -216 -319 216 319
use sky130_fd_pr__nfet_01v8_YYPCPJ  XM3
timestamp 0
transform 1 0 3012 0 1 746
box -2696 -252 2696 252
use sky130_fd_pr__nfet_01v8_YYPCPJ  XM4
timestamp 0
transform 1 0 8351 0 1 693
box -2696 -252 2696 252
use sky130_fd_pr__pfet_01v8_KVC9YE  XM7
timestamp 0
transform 1 0 14069 0 1 596
box -2696 -261 2696 261
use sky130_fd_pr__pfet_01v8_KVC9YE  XM9
timestamp 0
transform 1 0 19408 0 1 543
box -2696 -261 2696 261
use sky130_fd_pr__nfet_01v8_3STNDZ  XM10
timestamp 0
transform 1 0 22262 0 1 2939
box -211 -2710 211 2710
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
