* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : pre_therm                                    *
* Netlisted  : Mon Dec  9 01:54:35 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_C_CDNS_733705663440                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_C_CDNS_733705663440 1
** N=1 EP=1 FDC=0
.ends M1M2_C_CDNS_733705663440

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2M3_C_CDNS_733705663441                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2M3_C_CDNS_733705663441 1
** N=1 EP=1 FDC=0
.ends M2M3_C_CDNS_733705663441

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_C_CDNS_733705663442                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_C_CDNS_733705663442 1
** N=1 EP=1 FDC=0
.ends M1M2_C_CDNS_733705663442

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3M4_C_CDNS_733705663443                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3M4_C_CDNS_733705663443 1
** N=1 EP=1 FDC=0
.ends M3M4_C_CDNS_733705663443

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: PYL1CON_C_CDNS_733705663444                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt PYL1CON_C_CDNS_733705663444 1 2
** N=2 EP=2 FDC=0
.ends PYL1CON_C_CDNS_733705663444

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_733705663445                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_733705663445 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_733705663445

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_733705663446                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_733705663446 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_733705663446

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_733705663447                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_733705663447 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_733705663447

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733705663440                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733705663440 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6.5e-07 W=4.45e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733705663440

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733705663441                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733705663441 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=6.3e-07 W=7.9e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733705663441

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv01f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv01f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=575 1630 0 0 $X=390 $Y=1445
X1 3 L1M1_C_CDNS_733705663445 $T=575 1630 0 0 $X=410 $Y=1485
X2 4 L1M1_C_CDNS_733705663446 $T=1065 3205 0 0 $X=950 $Y=2860
X3 4 L1M1_C_CDNS_733705663447 $T=1085 695 0 0 $X=970 $Y=530
X4 2 4 3 nfet_01v8_CDNS_733705663440 $T=295 475 0 0 $X=-110 $Y=325
X5 1 4 3 pfet_01v8_CDNS_733705663441 $T=295 2820 0 0 $X=-150 $Y=2640
.ends inv01f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_733705663448                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_733705663448 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_733705663448

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733705663442                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733705663442 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 pfet_01v8 L=1.05e-06 W=5.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733705663442

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733705663443                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733705663443 1 2 3 4
** N=10 EP=4 FDC=1
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=1.02e-06 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733705663443

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: preampF                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt preampF 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=415 2135 0 0 $X=230 $Y=1950
X1 3 L1M1_C_CDNS_733705663445 $T=415 2135 0 0 $X=250 $Y=1990
X2 4 L1M1_C_CDNS_733705663447 $T=1100 3570 0 90 $X=935 $Y=3455
X3 1 L1M1_C_CDNS_733705663448 $T=130 995 0 0 $X=15 $Y=470
X4 4 L1M1_C_CDNS_733705663448 $T=570 995 0 0 $X=455 $Y=470
X5 4 2 3 1 pfet_01v8_CDNS_733705663442 $T=825 3430 0 270 $X=645 $Y=1935
X6 4 1 3 2 nfet_01v8_CDNS_733705663443 $T=430 485 1 180 $X=-125 $Y=335
.ends preampF

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733705663444                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733705663444 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.5e-07 W=8e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733705663444

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733705663445                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733705663445 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=2.85e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733705663445

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv02f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv02f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=460 1630 0 0 $X=275 $Y=1445
X1 3 L1M1_C_CDNS_733705663445 $T=460 1630 0 0 $X=295 $Y=1485
X2 4 L1M1_C_CDNS_733705663446 $T=725 3245 0 0 $X=610 $Y=2900
X3 4 L1M1_C_CDNS_733705663447 $T=740 850 0 0 $X=625 $Y=685
X4 1 4 3 pfet_01v8_CDNS_733705663444 $T=335 2855 0 0 $X=-110 $Y=2675
X5 2 4 3 nfet_01v8_CDNS_733705663445 $T=315 640 0 0 $X=-90 $Y=490
.ends inv02f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733705663446                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733705663446 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 pfet_01v8 L=2.5e-07 W=5.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733705663446

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733705663447                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733705663447 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 nfet_01v8 L=5.5e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733705663447

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: preamp1F                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt preamp1F 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=810 990 0 0 $X=625 $Y=805
X1 3 L1M1_C_CDNS_733705663445 $T=810 990 0 0 $X=645 $Y=845
X2 4 L1M1_C_CDNS_733705663446 $T=725 1970 0 0 $X=610 $Y=1625
X3 4 2 3 1 pfet_01v8_CDNS_733705663446 $T=840 2840 0 90 $X=110 $Y=2395
X4 4 1 3 2 nfet_01v8_CDNS_733705663447 $T=610 1275 0 270 $X=460 $Y=320
.ends preamp1F

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733705663448                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733705663448 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=3.5e-07 W=6.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733705663448

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733705663449                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733705663449 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=4.5e-07 W=6.4e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733705663449

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv03f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv03f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=510 1870 0 0 $X=325 $Y=1685
X1 3 L1M1_C_CDNS_733705663445 $T=510 1870 0 0 $X=345 $Y=1725
X2 4 L1M1_C_CDNS_733705663446 $T=825 3370 0 0 $X=710 $Y=3025
X3 4 L1M1_C_CDNS_733705663446 $T=880 960 0 0 $X=765 $Y=615
X4 1 4 3 pfet_01v8_CDNS_733705663448 $T=335 3045 0 0 $X=-110 $Y=2865
X5 2 4 3 nfet_01v8_CDNS_733705663449 $T=290 640 0 0 $X=-115 $Y=490
.ends inv03f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634410                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634410 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.9e-07 W=6.2e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634410

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634411                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634411 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6e-07 W=7.05e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634411

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv04f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv04f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=575 1030 0 0 $X=390 $Y=845
X1 3 L1M1_C_CDNS_733705663445 $T=575 1030 0 0 $X=410 $Y=885
X2 4 L1M1_C_CDNS_733705663446 $T=710 2960 0 0 $X=595 $Y=2615
X3 4 L1M1_C_CDNS_733705663446 $T=1025 1070 0 0 $X=910 $Y=725
X4 1 4 3 pfet_01v8_CDNS_7337056634410 $T=380 2650 0 0 $X=-65 $Y=2470
X5 2 4 3 nfet_01v8_CDNS_7337056634411 $T=280 715 0 0 $X=-125 $Y=565
.ends inv04f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634412                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634412 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=6.95e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634412

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634413                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634413 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=4e-07 W=6.5e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634413

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv05f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv05f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=510 1810 0 0 $X=325 $Y=1625
X1 3 L1M1_C_CDNS_733705663445 $T=510 1810 0 0 $X=345 $Y=1665
X2 4 L1M1_C_CDNS_733705663446 $T=650 3170 0 0 $X=535 $Y=2825
X3 4 L1M1_C_CDNS_733705663446 $T=855 960 0 0 $X=740 $Y=615
X4 1 4 3 pfet_01v8_CDNS_7337056634412 $T=360 2825 0 0 $X=-85 $Y=2645
X5 2 4 3 nfet_01v8_CDNS_7337056634413 $T=315 630 0 0 $X=-90 $Y=480
.ends inv05f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634414                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634414 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3.2e-07 W=7.25e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634414

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634415                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634415 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=4.35e-07 W=5.6e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634415

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv06f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv06f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=555 2320 0 0 $X=370 $Y=2135
X1 3 L1M1_C_CDNS_733705663445 $T=555 2320 0 0 $X=390 $Y=2175
X2 4 L1M1_C_CDNS_733705663446 $T=855 1035 0 0 $X=740 $Y=690
X3 4 L1M1_C_CDNS_733705663447 $T=910 3285 0 0 $X=795 $Y=3120
X4 2 4 3 nfet_01v8_CDNS_7337056634414 $T=395 685 0 0 $X=-10 $Y=535
X5 1 4 3 pfet_01v8_CDNS_7337056634415 $T=335 3005 0 0 $X=-110 $Y=2825
.ends inv06f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634416                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634416 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3e-07 W=9.8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634416

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634417                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634417 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.55e-07 W=5.7e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634417

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv07f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv07f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=435 2320 0 0 $X=250 $Y=2135
X1 3 L1M1_C_CDNS_733705663445 $T=435 2320 0 0 $X=270 $Y=2175
X2 4 L1M1_C_CDNS_733705663446 $T=755 940 0 0 $X=640 $Y=595
X3 4 L1M1_C_CDNS_733705663447 $T=655 3235 0 0 $X=540 $Y=3070
X4 2 4 3 nfet_01v8_CDNS_7337056634416 $T=315 460 0 0 $X=-90 $Y=310
X5 1 4 3 pfet_01v8_CDNS_7337056634417 $T=360 2950 0 0 $X=-85 $Y=2770
.ends inv07f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634418                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634418 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=9.9e-07 W=4.9e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634418

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634419                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634419 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.65e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634419

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv08f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv08f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=155 1745 0 0 $X=-30 $Y=1560
X1 3 L1M1_C_CDNS_733705663445 $T=155 1745 0 0 $X=-10 $Y=1600
X2 4 L1M1_C_CDNS_733705663446 $T=665 3170 0 0 $X=550 $Y=2825
X3 4 L1M1_C_CDNS_733705663447 $T=1035 1870 0 90 $X=870 $Y=1755
X4 2 4 3 nfet_01v8_CDNS_7337056634418 $T=1280 740 0 90 $X=640 $Y=335
X5 1 4 3 pfet_01v8_CDNS_7337056634419 $T=360 2755 0 0 $X=-85 $Y=2575
.ends inv08f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634420                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634420 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.1e-06 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634420

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634421                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634421 1 2 3
** N=9 EP=3 FDC=2
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.7e-07 $X=0 $Y=0 $dt=8
M1 1 3 2 1 pfet_01v8 L=1.5e-07 W=7.7e-07 $X=430 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634421

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv09f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv09f 1 2 3 4
** N=9 EP=4 FDC=3
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=20 2075 0 0 $X=-165 $Y=1890
X1 3 L1M1_C_CDNS_733705663445 $T=20 2075 0 0 $X=-145 $Y=1930
X2 4 L1M1_C_CDNS_733705663447 $T=670 1935 0 90 $X=505 $Y=1820
X3 4 L1M1_C_CDNS_733705663447 $T=690 3225 0 0 $X=575 $Y=3060
X4 2 4 3 nfet_01v8_CDNS_7337056634420 $T=905 695 0 90 $X=335 $Y=290
X5 1 4 3 pfet_01v8_CDNS_7337056634421 $T=400 2840 0 0 $X=-45 $Y=2660
.ends inv09f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634422                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634422 1 2 3
** N=7 EP=3 FDC=1
M0 2 2 1 3 pfet_01v8 L=1.5e-07 W=1e-06 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634422

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: div_fixed                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt div_fixed 1 2 3
** N=8 EP=3 FDC=2
X0 2 4 PYL1CON_C_CDNS_733705663444 $T=405 585 0 0 $X=220 $Y=400
X1 2 L1M1_C_CDNS_733705663445 $T=390 585 0 0 $X=225 $Y=440
X2 3 L1M1_C_CDNS_733705663446 $T=610 1390 0 0 $X=495 $Y=1045
X3 3 L1M1_C_CDNS_733705663447 $T=1350 2690 0 90 $X=1185 $Y=2575
X4 1 3 2 1 pfet_01v8_CDNS_733705663442 $T=1625 3880 1 270 $X=895 $Y=2385
X5 3 2 1 pfet_01v8_CDNS_7337056634422 $T=470 1900 0 180 $X=-125 $Y=720
.ends div_fixed

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634423                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634423 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.55e-07 W=9.45e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634423

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634424                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634424 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.45e-07 W=8.65e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634424

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv10f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv10f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=500 1860 0 0 $X=315 $Y=1675
X1 3 L1M1_C_CDNS_733705663445 $T=500 1860 0 0 $X=335 $Y=1715
X2 4 L1M1_C_CDNS_733705663446 $T=720 1035 0 0 $X=605 $Y=690
X3 4 L1M1_C_CDNS_733705663446 $T=770 3090 0 0 $X=655 $Y=2745
X4 2 4 3 nfet_01v8_CDNS_7337056634423 $T=425 555 0 0 $X=20 $Y=405
X5 1 4 3 pfet_01v8_CDNS_7337056634424 $T=385 2670 0 0 $X=-60 $Y=2490
.ends inv10f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634425                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634425 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=9.5e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634425

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634426                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634426 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.6e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634426

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv11f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv11f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=480 1765 0 0 $X=295 $Y=1580
X1 3 L1M1_C_CDNS_733705663445 $T=480 1765 0 0 $X=315 $Y=1620
X2 4 L1M1_C_CDNS_733705663446 $T=750 3045 0 0 $X=635 $Y=2700
X3 4 L1M1_C_CDNS_733705663447 $T=1305 910 0 0 $X=1190 $Y=745
X4 2 4 3 nfet_01v8_CDNS_7337056634425 $T=215 700 0 0 $X=-190 $Y=550
X5 1 4 3 pfet_01v8_CDNS_7337056634426 $T=350 2610 0 0 $X=-95 $Y=2430
.ends inv11f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634427                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634427 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3.3e-07 W=8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634427

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634428                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634428 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634428

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv12f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv12f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=465 2185 0 0 $X=280 $Y=2000
X1 3 L1M1_C_CDNS_733705663445 $T=465 2185 0 0 $X=300 $Y=2040
X2 4 L1M1_C_CDNS_733705663446 $T=675 3150 0 0 $X=560 $Y=2805
X3 4 L1M1_C_CDNS_733705663446 $T=810 965 0 0 $X=695 $Y=620
X4 2 4 3 nfet_01v8_CDNS_7337056634427 $T=340 555 0 0 $X=-65 $Y=405
X5 1 4 3 pfet_01v8_CDNS_7337056634428 $T=385 2785 0 0 $X=-60 $Y=2605
.ends inv12f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634429                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634429 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=5.5e-07 W=5.4e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634429

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634430                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634430 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.6e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634430

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv13f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv13f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=465 1790 0 0 $X=280 $Y=1605
X1 3 L1M1_C_CDNS_733705663445 $T=465 1790 0 0 $X=300 $Y=1645
X2 4 L1M1_C_CDNS_733705663446 $T=685 3120 0 0 $X=570 $Y=2775
X3 4 L1M1_C_CDNS_733705663447 $T=1050 915 0 0 $X=935 $Y=750
X4 2 4 3 nfet_01v8_CDNS_7337056634429 $T=360 720 0 0 $X=-45 $Y=570
X5 1 4 3 pfet_01v8_CDNS_7337056634430 $T=385 2685 0 0 $X=-60 $Y=2505
.ends inv13f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634431                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634431 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6.75e-07 W=4.8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634431

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634432                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634432 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.65e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634432

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv14f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv14f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=520 1745 0 0 $X=335 $Y=1560
X1 3 L1M1_C_CDNS_733705663445 $T=520 1745 0 0 $X=355 $Y=1600
X2 4 L1M1_C_CDNS_733705663446 $T=735 3095 0 0 $X=620 $Y=2750
X3 4 L1M1_C_CDNS_733705663447 $T=1165 915 0 0 $X=1050 $Y=750
X4 2 4 3 nfet_01v8_CDNS_7337056634431 $T=350 675 0 0 $X=-55 $Y=525
X5 1 4 3 pfet_01v8_CDNS_7337056634432 $T=445 2705 0 0 $X=0 $Y=2525
.ends inv14f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634433                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634433 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634433

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv15f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv15f 1 2 3 4
** N=9 EP=4 FDC=2
X0 3 5 PYL1CON_C_CDNS_733705663444 $T=700 1765 0 0 $X=515 $Y=1580
X1 3 L1M1_C_CDNS_733705663445 $T=700 1765 0 0 $X=535 $Y=1620
X2 4 L1M1_C_CDNS_733705663446 $T=910 3070 0 0 $X=795 $Y=2725
X3 4 L1M1_C_CDNS_733705663447 $T=1305 910 0 0 $X=1190 $Y=745
X4 2 4 3 nfet_01v8_CDNS_7337056634425 $T=215 700 0 0 $X=-190 $Y=550
X5 1 4 3 pfet_01v8_CDNS_7337056634433 $T=620 2635 0 0 $X=175 $Y=2455
.ends inv15f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pre_therm                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pre_therm 1 20 21 5 6 4 7 10 14 16
+ 11 13 9 12 15 17 18 19
** N=21 EP=18 FDC=37
X0 1 M1M2_C_CDNS_733705663440 $T=-685 1245 0 0 $X=-815 $Y=1085
X1 1 M1M2_C_CDNS_733705663440 $T=145 12545 0 0 $X=15 $Y=12385
X2 1 M1M2_C_CDNS_733705663440 $T=360 6515 0 0 $X=230 $Y=6355
X3 2 M1M2_C_CDNS_733705663440 $T=1095 7550 0 0 $X=965 $Y=7390
X4 3 M1M2_C_CDNS_733705663440 $T=2265 2075 0 90 $X=2105 $Y=1945
X5 2 M1M2_C_CDNS_733705663440 $T=2260 7550 0 0 $X=2130 $Y=7390
X6 4 M1M2_C_CDNS_733705663440 $T=2705 1035 0 0 $X=2575 $Y=875
X7 5 M1M2_C_CDNS_733705663440 $T=2840 8375 0 0 $X=2710 $Y=8215
X8 2 M1M2_C_CDNS_733705663440 $T=3885 7550 0 0 $X=3755 $Y=7390
X9 3 M1M2_C_CDNS_733705663440 $T=4000 1265 0 0 $X=3870 $Y=1105
X10 6 M1M2_C_CDNS_733705663440 $T=4235 8215 0 0 $X=4105 $Y=8055
X11 7 M1M2_C_CDNS_733705663440 $T=4520 1145 0 0 $X=4390 $Y=985
X12 8 M1M2_C_CDNS_733705663440 $T=4565 11390 0 90 $X=4405 $Y=11260
X13 9 M1M2_C_CDNS_733705663440 $T=5155 12860 0 0 $X=5025 $Y=12700
X14 1 M1M2_C_CDNS_733705663440 $T=5350 7260 0 90 $X=5190 $Y=7130
X15 3 M1M2_C_CDNS_733705663440 $T=5705 2075 0 90 $X=5545 $Y=1945
X16 10 M1M2_C_CDNS_733705663440 $T=6090 1145 0 0 $X=5960 $Y=985
X17 8 M1M2_C_CDNS_733705663440 $T=6190 11390 0 90 $X=6030 $Y=11260
X18 11 M1M2_C_CDNS_733705663440 $T=6245 7100 0 0 $X=6115 $Y=6940
X19 12 M1M2_C_CDNS_733705663440 $T=6500 12815 0 0 $X=6370 $Y=12655
X20 1 M1M2_C_CDNS_733705663440 $T=7015 6930 0 90 $X=6855 $Y=6800
X21 1 M1M2_C_CDNS_733705663440 $T=7515 2895 0 90 $X=7355 $Y=2765
X22 13 M1M2_C_CDNS_733705663440 $T=7635 7080 0 0 $X=7505 $Y=6920
X23 14 M1M2_C_CDNS_733705663440 $T=7830 1145 0 0 $X=7700 $Y=985
X24 8 M1M2_C_CDNS_733705663440 $T=7870 11390 0 90 $X=7710 $Y=11260
X25 15 M1M2_C_CDNS_733705663440 $T=8120 12815 0 0 $X=7990 $Y=12655
X26 1 M1M2_C_CDNS_733705663440 $T=9135 2895 0 90 $X=8975 $Y=2765
X27 8 M1M2_C_CDNS_733705663440 $T=9130 7340 0 0 $X=9000 $Y=7180
X28 16 M1M2_C_CDNS_733705663440 $T=9470 1145 0 0 $X=9340 $Y=985
X29 8 M1M2_C_CDNS_733705663440 $T=9500 11390 0 90 $X=9340 $Y=11260
X30 17 M1M2_C_CDNS_733705663440 $T=9760 12815 0 0 $X=9630 $Y=12655
X31 18 M1M2_C_CDNS_733705663440 $T=9845 8180 0 0 $X=9715 $Y=8020
X32 8 M1M2_C_CDNS_733705663440 $T=11005 7340 0 0 $X=10875 $Y=7180
X33 19 M1M2_C_CDNS_733705663440 $T=11710 7340 0 90 $X=11550 $Y=7210
X34 20 M2M3_C_CDNS_733705663441 $T=1140 13975 0 0 $X=775 $Y=13790
X35 21 M2M3_C_CDNS_733705663441 $T=1615 9305 0 0 $X=1250 $Y=9120
X36 21 M2M3_C_CDNS_733705663441 $T=1855 0 0 0 $X=1490 $Y=-185
X37 20 M2M3_C_CDNS_733705663441 $T=2840 4650 0 0 $X=2475 $Y=4465
X38 21 M2M3_C_CDNS_733705663441 $T=10560 0 0 0 $X=10195 $Y=-185
X39 21 M2M3_C_CDNS_733705663441 $T=10560 9320 0 0 $X=10195 $Y=9135
X40 20 M2M3_C_CDNS_733705663441 $T=11565 4660 0 0 $X=11200 $Y=4475
X41 20 M2M3_C_CDNS_733705663441 $T=11565 13980 0 0 $X=11200 $Y=13795
X42 20 M1M2_C_CDNS_733705663442 $T=1145 13970 0 0 $X=855 $Y=13810
X43 21 M1M2_C_CDNS_733705663442 $T=1615 9300 0 0 $X=1325 $Y=9140
X44 21 M1M2_C_CDNS_733705663442 $T=1855 -5 0 0 $X=1565 $Y=-165
X45 20 M1M2_C_CDNS_733705663442 $T=2820 4650 0 0 $X=2530 $Y=4490
X46 21 M1M2_C_CDNS_733705663442 $T=10560 0 0 0 $X=10270 $Y=-160
X47 21 M1M2_C_CDNS_733705663442 $T=10560 9320 0 0 $X=10270 $Y=9160
X48 20 M1M2_C_CDNS_733705663442 $T=11615 4655 0 0 $X=11325 $Y=4495
X49 20 M1M2_C_CDNS_733705663442 $T=11615 13975 0 0 $X=11325 $Y=13815
X50 20 M3M4_C_CDNS_733705663443 $T=1140 13975 0 0 $X=775 $Y=13785
X51 20 M3M4_C_CDNS_733705663443 $T=2835 4655 0 0 $X=2470 $Y=4465
X52 20 M3M4_C_CDNS_733705663443 $T=11570 4660 0 0 $X=11205 $Y=4470
X53 20 M3M4_C_CDNS_733705663443 $T=11570 13980 0 0 $X=11205 $Y=13790
X54 20 21 2 5 inv01f $T=1740 9060 1 0 $X=1560 $Y=4615
X55 20 21 1 2 preampF $T=0 9060 1 0 $X=-180 $Y=4615
X56 20 21 2 6 inv02f $T=3480 9060 1 0 $X=3300 $Y=4615
X57 20 21 1 3 preamp1F $T=0 255 0 0 $X=-180 $Y=-10
X58 20 21 3 4 inv03f $T=1740 260 0 0 $X=1560 $Y=-5
X59 20 21 3 7 inv04f $T=3480 260 0 0 $X=3300 $Y=-5
X60 20 21 3 10 inv05f $T=5220 260 0 0 $X=5040 $Y=-5
X61 20 21 1 14 inv06f $T=6960 260 0 0 $X=6780 $Y=-5
X62 20 21 1 16 inv07f $T=8700 260 0 0 $X=8520 $Y=-5
X63 20 21 1 11 inv08f $T=5220 9060 1 0 $X=5040 $Y=4615
X64 20 21 1 13 inv09f $T=6970 9060 1 0 $X=6780 $Y=4615
X65 1 21 8 div_fixed $T=0 9580 0 0 $X=-180 $Y=9315
X66 20 21 8 9 inv10f $T=4040 9585 0 0 $X=3860 $Y=9320
X67 20 21 8 12 inv11f $T=5735 9585 0 0 $X=5545 $Y=9320
X68 20 21 8 15 inv12f $T=7430 9580 0 0 $X=7250 $Y=9315
X69 20 21 8 17 inv13f $T=9060 9580 0 0 $X=8880 $Y=9315
X70 20 21 8 18 inv14f $T=8665 9060 1 0 $X=8485 $Y=4615
X71 20 21 8 19 inv15f $T=10360 9060 1 0 $X=10170 $Y=4615
.ends pre_therm
