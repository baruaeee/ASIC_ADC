magic
tech sky130A
magscale 1 2
timestamp 1696192394
<< nwell >>
rect -211 -319 211 319
<< pmos >>
rect -15 -100 15 100
<< pdiff >>
rect -73 88 -15 100
rect -73 -88 -61 88
rect -27 -88 -15 88
rect -73 -100 -15 -88
rect 15 88 73 100
rect 15 -88 27 88
rect 61 -88 73 88
rect 15 -100 73 -88
<< pdiffc >>
rect -61 -88 -27 88
rect 27 -88 61 88
<< nsubdiff >>
rect -175 249 -79 283
rect 79 249 175 283
rect -175 187 -141 249
rect 141 187 175 249
rect -175 -249 -141 -187
rect 141 -249 175 -187
rect -175 -283 -79 -249
rect 79 -283 175 -249
<< nsubdiffcont >>
rect -79 249 79 283
rect -175 -187 -141 187
rect 141 -187 175 187
rect -79 -283 79 -249
<< poly >>
rect -34 188 34 198
rect -34 154 -18 188
rect 18 154 34 188
rect -34 130 34 154
rect -15 100 15 130
rect -15 -130 15 -100
rect -34 -154 34 -130
rect -34 -188 -18 -154
rect 18 -188 34 -154
rect -34 -198 34 -188
<< polycont >>
rect -18 154 18 188
rect -18 -188 18 -154
<< locali >>
rect -175 249 -79 283
rect 79 249 175 283
rect -175 187 -141 249
rect -34 188 34 198
rect -34 154 -18 188
rect 18 154 34 188
rect -34 146 34 154
rect 141 187 175 249
rect -61 88 -27 104
rect -61 -104 -27 -88
rect 27 88 61 104
rect 27 -104 61 -88
rect -175 -249 -141 -187
rect -34 -154 34 -148
rect -34 -188 -18 -154
rect 18 -188 34 -154
rect -34 -198 34 -188
rect 141 -249 175 -187
rect -175 -283 -79 -249
rect 79 -283 175 -249
<< viali >>
rect -18 154 18 188
rect -61 -88 -27 88
rect 27 -88 61 88
rect -18 -188 18 -154
<< metal1 >>
rect -34 188 34 198
rect -34 154 -18 188
rect 18 154 34 188
rect -34 146 34 154
rect -67 88 -21 100
rect -67 -88 -61 88
rect -27 -88 -21 88
rect -67 -100 -21 -88
rect 21 88 67 100
rect 21 -88 27 88
rect 61 -88 67 88
rect 21 -100 67 -88
rect -34 -154 34 -148
rect -34 -188 -18 -154
rect 18 -188 34 -154
rect -34 -198 34 -188
<< properties >>
string FIXED_BBOX -158 -266 158 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
