magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect 22233 5511 22291 5517
rect 22233 5477 22245 5511
rect 22233 5471 22291 5477
<< error_s >>
rect 299 998 333 1016
rect 299 962 369 998
rect 316 928 387 962
rect 5637 928 5672 962
rect 11030 956 11065 963
rect 11030 945 11064 956
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 928
rect 5638 909 5672 928
rect 316 547 369 583
rect 5657 530 5672 909
rect 5691 875 5726 909
rect 5691 530 5725 875
rect 5691 496 5706 530
rect 10994 477 11064 945
rect 11181 888 11239 894
rect 11181 854 11193 888
rect 11181 848 11239 854
rect 11356 821 11390 875
rect 11181 560 11239 566
rect 11181 526 11193 560
rect 11181 520 11239 526
rect 10994 441 11047 477
rect 11375 424 11390 821
rect 11409 787 11444 821
rect 16694 787 16729 821
rect 22087 804 22121 822
rect 11409 424 11443 787
rect 16695 768 16729 787
rect 11409 390 11424 424
rect 16714 371 16729 768
rect 16748 734 16783 768
rect 16748 371 16782 734
rect 16748 337 16763 371
rect 22051 318 22121 804
rect 22233 401 22291 407
rect 22233 367 22245 401
rect 22233 361 22291 367
rect 22051 282 22104 318
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_KGSDF3  XM1
timestamp 1703732895
transform 1 0 158 0 1 3266
box -211 -2719 211 2719
use sky130_fd_pr__pfet_01v8_SKYSXJ  XM2
timestamp 1703732895
transform 1 0 11210 0 1 707
box -216 -319 216 319
use sky130_fd_pr__nfet_01v8_YYPCPJ  XM3
timestamp 1703732895
transform 1 0 3012 0 1 746
box -2696 -252 2696 252
use sky130_fd_pr__nfet_01v8_YYPCPJ  XM4
timestamp 1703732895
transform 1 0 8351 0 1 693
box -2696 -252 2696 252
use sky130_fd_pr__pfet_01v8_KVC9YE  XM7
timestamp 1703732895
transform 1 0 14069 0 1 596
box -2696 -261 2696 261
use sky130_fd_pr__pfet_01v8_KVC9YE  XM9
timestamp 1703732895
transform 1 0 19408 0 1 543
box -2696 -261 2696 261
use sky130_fd_pr__nfet_01v8_3STNDZ  XM10
timestamp 1703732895
transform 1 0 22262 0 1 2939
box -211 -2710 211 2710
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
