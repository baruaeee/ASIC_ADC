* NGSPICE file created from th12.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_P28Q2U a_n33_n232# a_15_n135# w_n211_n354# a_n73_n135#
+ VSUBS
X0 a_15_n135# a_n33_n232# a_n73_n135# w_n211_n354# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.28 as=0.391 ps=3.28 w=1.35 l=0.15
C0 a_n33_n232# a_n73_n135# 0.0258f
C1 a_n33_n232# w_n211_n354# 0.19f
C2 a_n33_n232# a_15_n135# 0.0258f
C3 a_n73_n135# w_n211_n354# 0.0279f
C4 a_n73_n135# a_15_n135# 0.218f
C5 a_15_n135# w_n211_n354# 0.0279f
C6 a_15_n135# VSUBS 0.115f
C7 a_n73_n135# VSUBS 0.115f
C8 a_n33_n232# VSUBS 0.146f
C9 w_n211_n354# VSUBS 0.983f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZMY3VB a_n348_n42# a_n290_n130# a_n450_n182# a_290_n42#
X0 a_290_n42# a_n290_n130# a_n348_n42# a_n450_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.9
C0 a_n348_n42# a_290_n42# 0.00961f
C1 a_n348_n42# a_n290_n130# 0.0217f
C2 a_290_n42# a_n290_n130# 0.0217f
C3 a_290_n42# a_n450_n182# 0.076f
C4 a_n348_n42# a_n450_n182# 0.0839f
C5 a_n290_n130# a_n450_n182# 1.6f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n33_n197# a_n73_n100# 0.0236f
C1 a_n33_n197# w_n211_n319# 0.189f
C2 a_n33_n197# a_15_n100# 0.0236f
C3 a_n73_n100# w_n211_n319# 0.0248f
C4 a_n73_n100# a_15_n100# 0.162f
C5 a_15_n100# w_n211_n319# 0.0248f
C6 a_15_n100# VSUBS 0.0885f
C7 a_n73_n100# VSUBS 0.0885f
C8 a_n33_n197# VSUBS 0.145f
C9 w_n211_n319# VSUBS 0.894f
.ends

.subckt sky130_fd_pr__pfet_01v8_WV9GCW a_n158_n42# w_n296_n261# a_n100_n139# a_100_n42#
+ VSUBS
X0 a_100_n42# a_n100_n139# a_n158_n42# w_n296_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1
C0 a_n100_n139# a_n158_n42# 0.0144f
C1 a_n100_n139# w_n296_n261# 0.346f
C2 a_n100_n139# a_100_n42# 0.0144f
C3 a_n158_n42# w_n296_n261# 0.0224f
C4 a_n158_n42# a_100_n42# 0.024f
C5 a_100_n42# w_n296_n261# 0.0224f
C6 a_100_n42# VSUBS 0.0504f
C7 a_n158_n42# VSUBS 0.0504f
C8 a_n100_n139# VSUBS 0.353f
C9 w_n296_n261# VSUBS 1.06f
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n141_240# a_n33_n188# a_15_n100#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n141_240# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n73_n100# a_15_n100# 0.162f
C1 a_n73_n100# a_n33_n188# 0.0254f
C2 a_15_n100# a_n33_n188# 0.0254f
C3 a_15_n100# a_n141_240# 0.113f
C4 a_n73_n100# a_n141_240# 0.113f
C5 a_n33_n188# a_n141_240# 0.322f
.ends

.subckt th12 Vp V12 Vin Vn
XXM0 Vn Vn Vp m1_394_n856# Vn sky130_fd_pr__pfet_01v8_P28Q2U
XXM1 m1_529_n42# Vin Vn m1_394_n856# sky130_fd_pr__nfet_01v8_ZMY3VB
XXM2 m1_529_n42# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM3 Vp Vp m1_529_n42# V12 Vn sky130_fd_pr__pfet_01v8_WV9GCW
XXM4 V12 Vn m1_529_n42# Vn sky130_fd_pr__nfet_01v8_648S5X
C0 Vn Vin 0.135f
C1 Vp Vin 0.238f
C2 m1_529_n42# V12 0.0929f
C3 V12 m1_394_n856# 4.74e-19
C4 m1_529_n42# m1_394_n856# 0.0134f
C5 Vn V12 0.0234f
C6 Vp V12 0.0454f
C7 Vn m1_529_n42# 0.254f
C8 Vn m1_394_n856# 0.0338f
C9 Vp m1_529_n42# 0.322f
C10 Vp m1_394_n856# 0.04f
C11 Vn Vp 0.132f
C12 Vin V12 0.00205f
C13 Vin m1_529_n42# 0.0965f
C14 Vin m1_394_n856# 0.321f
C15 Vn 0 0.29f
C16 Vp 0 2.88f
C17 m1_529_n42# 0 0.861f
C18 V12 0 0.359f
C19 m1_394_n856# 0 0.215f
C20 Vin 0 1.9f
.ends

