magic
tech sky130A
magscale 1 2
timestamp 1704962958
<< pwell >>
rect -493 -258 493 258
<< nmos >>
rect -297 -48 297 48
<< ndiff >>
rect -355 36 -297 48
rect -355 -36 -343 36
rect -309 -36 -297 36
rect -355 -48 -297 -36
rect 297 36 355 48
rect 297 -36 309 36
rect 343 -36 355 36
rect 297 -48 355 -36
<< ndiffc >>
rect -343 -36 -309 36
rect 309 -36 343 36
<< psubdiff >>
rect -457 188 -361 222
rect 361 188 457 222
rect -457 126 -423 188
rect 423 126 457 188
rect -457 -188 -423 -126
rect 423 -188 457 -126
rect -457 -222 -361 -188
rect 361 -222 457 -188
<< psubdiffcont >>
rect -361 188 361 222
rect -457 -126 -423 126
rect 423 -126 457 126
rect -361 -222 361 -188
<< poly >>
rect -297 120 297 136
rect -297 86 -281 120
rect 281 86 297 120
rect -297 48 297 86
rect -297 -86 297 -48
rect -297 -120 -281 -86
rect 281 -120 297 -86
rect -297 -136 297 -120
<< polycont >>
rect -281 86 281 120
rect -281 -120 281 -86
<< locali >>
rect -457 188 -361 222
rect 361 188 457 222
rect -457 126 -423 188
rect 423 126 457 188
rect -297 86 -281 120
rect 281 86 297 120
rect -343 36 -309 52
rect -343 -52 -309 -36
rect 309 36 343 52
rect 309 -52 343 -36
rect -297 -120 -281 -86
rect 281 -120 297 -86
rect -457 -188 -423 -126
rect 423 -188 457 -126
rect -457 -222 -361 -188
rect 361 -222 457 -188
<< viali >>
rect -281 86 281 120
rect -343 -36 -309 36
rect 309 -36 343 36
rect -281 -120 281 -86
<< metal1 >>
rect -293 120 293 126
rect -293 86 -281 120
rect 281 86 293 120
rect -293 80 293 86
rect -349 36 -303 48
rect -349 -36 -343 36
rect -309 -36 -303 36
rect -349 -48 -303 -36
rect 303 36 349 48
rect 303 -36 309 36
rect 343 -36 349 36
rect 303 -48 349 -36
rect -293 -86 293 -80
rect -293 -120 -281 -86
rect 281 -120 293 -86
rect -293 -126 293 -120
<< properties >>
string FIXED_BBOX -440 -205 440 205
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.48 l 2.97 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
