magic
tech sky130A
magscale 1 2
timestamp 1706224144
<< error_p >>
rect -29 123 29 129
rect -29 89 -17 123
rect -29 83 29 89
rect -29 -89 29 -83
rect -29 -123 -17 -89
rect -29 -129 29 -123
<< nwell >>
rect -215 -261 215 261
<< pmos >>
rect -19 -42 19 42
<< pdiff >>
rect -77 30 -19 42
rect -77 -30 -65 30
rect -31 -30 -19 30
rect -77 -42 -19 -30
rect 19 30 77 42
rect 19 -30 31 30
rect 65 -30 77 30
rect 19 -42 77 -30
<< pdiffc >>
rect -65 -30 -31 30
rect 31 -30 65 30
<< nsubdiff >>
rect 145 129 179 191
rect 145 -191 179 -129
<< nsubdiffcont >>
rect 145 -129 179 129
<< poly >>
rect -33 123 33 139
rect -33 89 -17 123
rect 17 89 33 123
rect -33 73 33 89
rect -19 42 19 73
rect -19 -73 19 -42
rect -33 -89 33 -73
rect -33 -123 -17 -89
rect 17 -123 33 -89
rect -33 -139 33 -123
<< polycont >>
rect -17 89 17 123
rect -17 -123 17 -89
<< locali >>
rect 145 129 179 191
rect -33 89 -17 123
rect 17 89 33 123
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect -33 -123 -17 -89
rect 17 -123 33 -89
rect 145 -191 179 -129
<< viali >>
rect -17 89 17 123
rect -65 -30 -31 30
rect 31 -30 65 30
rect -17 -123 17 -89
<< metal1 >>
rect -29 123 29 129
rect -29 89 -17 123
rect 17 89 29 123
rect -29 83 29 89
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect -29 -89 29 -83
rect -29 -123 -17 -89
rect 17 -123 29 -89
rect -29 -129 29 -123
<< properties >>
string FIXED_BBOX -162 -208 162 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.193 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
