magic
tech sky130A
timestamp 1703731503
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
rect 0 -1400 100 -1300
rect 0 -1600 100 -1500
rect 0 -1800 100 -1700
rect 0 -2000 100 -1900
rect 0 -2200 100 -2100
rect 0 -2400 100 -2300
rect 0 -2600 100 -2500
rect 0 -2800 100 -2700
rect 0 -3000 100 -2900
rect 0 -3200 100 -3100
rect 0 -3400 100 -3300
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 Vp
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 Vin
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 V1
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 V2
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 V3
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 V4
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 128 0 0 0 V5
port 6 nsew
flabel metal1 0 -1400 100 -1300 0 FreeSans 128 0 0 0 V6
port 7 nsew
flabel metal1 0 -1600 100 -1500 0 FreeSans 128 0 0 0 V7
port 8 nsew
flabel metal1 0 -1800 100 -1700 0 FreeSans 128 0 0 0 V8
port 9 nsew
flabel metal1 0 -2000 100 -1900 0 FreeSans 128 0 0 0 V9
port 10 nsew
flabel metal1 0 -2200 100 -2100 0 FreeSans 128 0 0 0 V10
port 11 nsew
flabel metal1 0 -2400 100 -2300 0 FreeSans 128 0 0 0 V11
port 12 nsew
flabel metal1 0 -2600 100 -2500 0 FreeSans 128 0 0 0 V12
port 13 nsew
flabel metal1 0 -2800 100 -2700 0 FreeSans 128 0 0 0 V13
port 14 nsew
flabel metal1 0 -3000 100 -2900 0 FreeSans 128 0 0 0 V14
port 15 nsew
flabel metal1 0 -3200 100 -3100 0 FreeSans 128 0 0 0 V15
port 16 nsew
flabel metal1 0 -3400 100 -3300 0 FreeSans 128 0 0 0 Vn
port 17 nsew
<< end >>
