magic
tech sky130A
magscale 1 2
timestamp 1705440138
<< checkpaint >>
rect 13096 9618 17512 10758
rect 6417 8812 17512 9618
rect 6417 6586 28808 8812
rect 5239 4922 28808 6586
rect 5239 4548 34599 4922
rect 4698 4500 34599 4548
rect -1260 3840 34599 4500
rect 35267 3840 56721 10534
rect -1260 -660 56721 3840
rect 4636 -2490 28808 -660
rect 6218 -3719 28808 -2490
rect 7354 -9982 28808 -3719
rect 35267 -8260 56721 -660
<< locali >>
rect 7822 1386 7862 1388
rect 7800 1354 7862 1386
rect 7822 1296 7862 1354
<< viali >>
rect 7822 1258 7862 1296
<< metal1 >>
rect 7027 5155 7085 5395
rect 6663 4143 7083 4201
rect 6663 2795 6721 4143
rect 7018 3232 7078 3238
rect 7078 3168 7312 3228
rect 7018 3158 7078 3164
rect 6394 1152 6454 2306
rect 9990 1926 9996 1978
rect 10057 1948 10063 1978
rect 10057 1926 10064 1948
rect 9990 1886 10064 1926
rect 9990 1884 10062 1886
rect 7811 1302 7873 1308
rect 7810 1296 7874 1302
rect 7810 1258 7822 1296
rect 7862 1258 7874 1296
rect 7810 1252 7874 1258
rect 8715 1287 8753 1405
rect 9090 1294 9142 1300
rect 6394 1092 6526 1152
rect 7811 1133 7873 1252
rect 8715 1249 9090 1287
rect 9090 1236 9142 1242
rect 9806 1172 9858 1176
rect 8888 1170 9864 1172
rect 6466 710 6526 1092
rect 7167 1071 7963 1133
rect 8888 1110 9806 1170
rect 9858 1110 9864 1170
rect 8888 1108 9864 1110
rect 8888 1072 8952 1108
rect 9806 1104 9858 1108
rect 7080 600 7678 660
rect 7618 222 7678 600
rect 7901 599 7963 1071
rect 9728 983 9773 1046
rect 10687 1014 10738 1035
rect 9936 986 9988 992
rect 9728 938 9936 983
rect 9728 868 9773 938
rect 9936 928 9988 934
rect 10682 986 10738 1014
rect 10682 934 10686 986
rect 10682 928 10738 934
rect 12471 534 12477 586
rect 12534 534 12540 586
rect 9516 404 9752 440
rect 7612 162 7618 222
rect 7678 162 7684 222
rect 6703 67 6741 93
rect 6703 45 8429 67
rect 6703 7 8454 45
rect 9042 -67 9270 -65
rect 9042 -119 9211 -67
rect 9274 -119 9280 -67
rect 9042 -121 9270 -119
rect 9516 -418 9552 404
rect 12482 351 12529 534
rect 8924 -454 9552 -418
rect 6406 -630 6412 -570
rect 6472 -630 6542 -570
rect 6620 -807 6654 -741
rect 8924 -1160 8960 -454
rect 9642 -663 9891 -653
rect 9642 -717 9653 -663
rect 9705 -717 9891 -663
rect 9642 -727 9891 -717
rect 7614 -1196 9746 -1160
rect 9710 -1852 9746 -1196
rect 12240 -1240 12246 -1188
rect 12302 -1190 12308 -1188
rect 12302 -1238 12398 -1190
rect 12302 -1240 12308 -1238
rect 9710 -1888 9960 -1852
<< via1 >>
rect 7018 3164 7078 3232
rect 9996 1926 10057 1978
rect 9090 1242 9142 1294
rect 9806 1110 9858 1170
rect 9936 934 9988 986
rect 10686 934 10738 986
rect 12477 534 12534 586
rect 7618 162 7678 222
rect 9211 -119 9274 -67
rect 6412 -630 6472 -570
rect 9653 -717 9705 -663
rect 12246 -1240 12302 -1188
<< metal2 >>
rect 6770 5361 8254 5429
rect 6770 3232 6838 5361
rect 6770 3164 7018 3232
rect 7078 3164 7084 3232
rect 9996 2165 10057 2168
rect 9962 2109 9971 2165
rect 10081 2109 10090 2165
rect 9996 1978 10057 2109
rect 9996 1920 10057 1926
rect 9084 1242 9090 1294
rect 9142 1284 9148 1294
rect 9142 1252 10102 1284
rect 9142 1242 9148 1252
rect 9867 1195 9923 1204
rect 9800 1110 9806 1170
rect 9858 1110 9867 1170
rect 9923 1110 9925 1170
rect 9867 1076 9923 1085
rect 9930 934 9936 986
rect 9988 976 9994 986
rect 10070 976 10102 1252
rect 10680 976 10686 986
rect 9988 944 10686 976
rect 9988 934 9994 944
rect 10680 934 10686 944
rect 10738 934 10744 986
rect 12477 653 12533 662
rect 12533 591 12534 651
rect 12477 586 12534 591
rect 12477 528 12534 534
rect 7618 222 7678 228
rect 7618 156 7678 162
rect 7624 -94 7672 156
rect 9211 -67 9274 -61
rect 6418 -142 7672 -94
rect 7961 -93 8017 -84
rect 6418 -564 6466 -142
rect 7798 -148 7961 -100
rect 7961 -164 8017 -155
rect 9202 -167 9211 -111
rect 9274 -119 9282 -111
rect 9273 -167 9282 -119
rect 9211 -170 9274 -167
rect 6412 -570 6472 -564
rect 6412 -636 6472 -630
rect 9595 -659 9651 -650
rect 9651 -717 9653 -663
rect 9705 -717 9711 -663
rect 9595 -730 9651 -721
rect 12246 -1184 12302 -1182
rect 12154 -1188 12302 -1184
rect 12154 -1240 12246 -1188
rect 12246 -1246 12302 -1240
<< via2 >>
rect 9971 2109 10081 2165
rect 9867 1085 9923 1195
rect 12477 591 12533 653
rect 7961 -155 8017 -93
rect 9211 -119 9273 -111
rect 9211 -167 9273 -119
rect 9595 -721 9651 -659
<< metal3 >>
rect 9966 2165 10086 2170
rect 9966 2109 9971 2165
rect 10081 2109 10086 2165
rect 9966 1968 10086 2109
rect 9862 1195 10290 1200
rect 9862 1085 9867 1195
rect 9923 1085 10290 1195
rect 9862 1080 10290 1085
rect 9726 653 12538 658
rect 9726 591 12477 653
rect 12533 591 12538 653
rect 9726 586 12538 591
rect 9726 104 9798 586
rect 8878 32 9798 104
rect 8878 -88 8950 32
rect 7954 -93 8950 -88
rect 7954 -155 7961 -93
rect 8017 -155 8950 -93
rect 7954 -160 8950 -155
rect 9206 -111 9278 -106
rect 9206 -167 9211 -111
rect 9273 -167 9278 -111
rect 9206 -654 9278 -167
rect 9206 -659 9656 -654
rect 9206 -721 9595 -659
rect 9651 -721 9656 -659
rect 9206 -726 9656 -721
<< metal4 >>
rect 12436 5330 12492 5360
use therm  therm_0
timestamp 1705440138
transform 1 0 37473 0 1 600
box -946 -7600 17988 8674
use Analog  x1
timestamp 1705195269
transform 1 0 18064 0 1 7400
box -12168 -9924 -170 2098
use therm  x2
timestamp 1705440138
transform 1 0 9560 0 1 -1122
box -946 -7600 17988 8674
use th02  x16
timestamp 1705440134
transform 1 0 0 0 1 2560
box 0 -1960 4395 680
use th03  x17
timestamp 1705440134
transform 1 0 4395 0 1 1800
box 0 -1200 1840 706
use th04  x18
timestamp 1705440135
transform 1 0 6235 0 1 1900
box 0 -1300 1216 476
use th05  x19
timestamp 1705440135
transform 1 0 7451 0 1 1800
box 0 -1200 2064 258
use th06  x20
timestamp 1705440135
transform 1 0 9515 0 1 1800
box 0 -1200 1542 200
use th07  x21
timestamp 1705440135
transform 1 0 11057 0 1 1890
box 0 -1290 1462 200
use th08  x22
timestamp 1705440135
transform 1 0 12519 0 1 1992
box 0 -1392 1396 200
use th09  x23
timestamp 1705440135
transform 1 0 13915 0 1 2098
box 0 -1498 1918 398
use th10  x24
timestamp 1705440135
transform 1 0 15833 0 1 1800
box 0 -1200 1590 790
use th11  x25
timestamp 1705440136
transform 1 0 17423 0 1 1800
box 0 -1200 1584 1464
use th12  x26
timestamp 1705440136
transform 1 0 19007 0 1 1800
box 0 -1200 1662 716
use th13  x27
timestamp 1705440136
transform 1 0 20669 0 1 1800
box 0 -1200 2062 556
use th14  x28
timestamp 1705440136
transform 1 0 22731 0 1 1800
box 0 -1200 4172 772
use th15  x29
timestamp 1705440136
transform 1 0 26903 0 1 1800
box 0 -1200 6436 1862
use preamp  x30
timestamp 1705440136
transform 1 0 33339 0 1 1800
box 0 -1200 1470 780
use th01  x31
timestamp 1705440137
transform 1 0 34809 0 1 1800
box 0 -1200 2664 200
<< end >>
