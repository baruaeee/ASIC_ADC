magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_s >>
rect 6497 1926 6531 1944
rect 6497 1890 6567 1926
rect 6514 1856 6585 1890
rect 3028 999 3063 1033
rect 6181 1016 6215 1034
rect 3029 980 3063 999
rect 3048 583 3063 980
rect 3082 946 3117 980
rect 3082 583 3116 946
rect 3082 549 3097 583
rect 6145 530 6215 1016
rect 6327 613 6385 619
rect 6327 579 6339 613
rect 6327 573 6385 579
rect 6145 494 6198 530
rect 6514 477 6584 1856
rect 6696 1788 6754 1794
rect 6696 1754 6708 1788
rect 6696 1748 6754 1754
rect 6866 839 6900 857
rect 8358 850 8393 857
rect 8358 839 8392 850
rect 6866 803 6936 839
rect 6883 769 6954 803
rect 6696 560 6754 566
rect 6696 526 6708 560
rect 6696 520 6754 526
rect 6514 441 6567 477
rect 6883 424 6953 769
rect 6883 388 6936 424
rect 8322 371 8392 839
rect 8504 782 8562 788
rect 8504 748 8516 782
rect 8504 742 8562 748
rect 8504 454 8562 460
rect 8504 420 8516 454
rect 8504 414 8562 420
rect 8322 335 8375 371
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_Y3KFQV  XM4
timestamp 1703732895
transform 1 0 1523 0 1 808
box -1576 -261 1576 261
use sky130_fd_pr__pfet_01v8_Y3KFQV  XM5
timestamp 1703732895
transform 1 0 4622 0 1 755
box -1576 -261 1576 261
use sky130_fd_pr__nfet_01v8_NLLP5F  XM6
timestamp 1703732895
transform 1 0 6356 0 1 2031
box -211 -1590 211 1590
use sky130_fd_pr__pfet_01v8_UJPVTG  XM8
timestamp 1703732895
transform 1 0 6725 0 1 1157
box -211 -769 211 769
use sky130_fd_pr__nfet_01v8_ZFMUVB  XM11
timestamp 1703732895
transform 1 0 7629 0 1 587
box -746 -252 746 252
use sky130_fd_pr__pfet_01v8_XGS3BL  XM12
timestamp 1703732895
transform 1 0 8533 0 1 601
box -211 -319 211 319
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
