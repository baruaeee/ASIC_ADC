* NGSPICE file created from th01.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_3QB9EZ a_n296_n139# a_n354_n42# a_296_n42# w_n492_n261#
+ VSUBS
X0 a_296_n42# a_n296_n139# a_n354_n42# w_n492_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.96
C0 a_n296_n139# w_n492_n261# 1.04f
C1 a_n296_n139# a_296_n42# 0.0218f
C2 a_296_n42# w_n492_n261# 0.0498f
C3 a_n296_n139# a_n354_n42# 0.0218f
C4 a_n354_n42# w_n492_n261# 0.0498f
C5 a_296_n42# a_n354_n42# 0.00943f
C6 a_296_n42# VSUBS 0.0352f
C7 a_n354_n42# VSUBS 0.0352f
C8 a_n296_n139# VSUBS 0.797f
C9 w_n492_n261# VSUBS 2.19f
.ends

.subckt sky130_fd_pr__nfet_01v8_J2SMPG a_n33_n398# a_15_n310# a_n175_n484# a_n73_n310#
X0 a_15_n310# a_n33_n398# a_n73_n310# a_n175_n484# sky130_fd_pr__nfet_01v8 ad=0.899 pd=6.78 as=0.899 ps=6.78 w=3.1 l=0.15
C0 a_n73_n310# a_n33_n398# 0.0365f
C1 a_n73_n310# a_15_n310# 0.496f
C2 a_15_n310# a_n33_n398# 0.0365f
C3 a_15_n310# a_n175_n484# 0.345f
C4 a_n73_n310# a_n175_n484# 0.345f
C5 a_n33_n398# a_n175_n484# 0.349f
.ends

.subckt sky130_fd_pr__nfet_01v8_G45C34 a_297_n48# a_n297_n136# a_n457_n222# a_n355_n48#
X0 a_297_n48# a_n297_n136# a_n355_n48# a_n457_n222# sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.54 as=0.139 ps=1.54 w=0.48 l=2.97
C0 a_n355_n48# a_n297_n136# 0.0239f
C1 a_n355_n48# a_297_n48# 0.0107f
C2 a_297_n48# a_n297_n136# 0.0239f
C3 a_297_n48# a_n457_n222# 0.0929f
C4 a_n355_n48# a_n457_n222# 0.0929f
C5 a_n297_n136# a_n457_n222# 1.8f
.ends

.subckt sky130_fd_pr__pfet_01v8_XA2NHL a_15_n310# w_n211_n529# a_n73_n310# a_n33_n407#
+ VSUBS
X0 a_15_n310# a_n33_n407# a_n73_n310# w_n211_n529# sky130_fd_pr__pfet_01v8 ad=0.899 pd=6.78 as=0.899 ps=6.78 w=3.1 l=0.15
C0 a_n33_n407# w_n211_n529# 0.241f
C1 a_n33_n407# a_15_n310# 0.0346f
C2 a_15_n310# w_n211_n529# 0.21f
C3 a_n33_n407# a_n73_n310# 0.0346f
C4 a_n73_n310# w_n211_n529# 0.21f
C5 a_15_n310# a_n73_n310# 0.496f
C6 a_15_n310# VSUBS 0.135f
C7 a_n73_n310# VSUBS 0.135f
C8 a_n33_n407# VSUBS 0.121f
C9 w_n211_n529# VSUBS 1.97f
.ends

.subckt th01 Vp Vin Vout Vn
XXM2 Vin Vp m1_931_n929# Vp Vn sky130_fd_pr__pfet_01v8_3QB9EZ
XXM3 Vin m1_931_n929# Vn Vn sky130_fd_pr__nfet_01v8_J2SMPG
XXM4 Vn m1_931_n929# Vn Vout sky130_fd_pr__nfet_01v8_G45C34
XXM5 Vp Vp Vout m1_931_n929# Vn sky130_fd_pr__pfet_01v8_XA2NHL
C0 Vin Vp 0.391f
C1 Vin Vout 5.64e-20
C2 Vin Vn 0.0908f
C3 Vin m1_931_n929# 0.206f
C4 Vp Vout 0.0877f
C5 Vp Vn 0.338f
C6 Vout Vn 0.0892f
C7 Vp m1_931_n929# 0.324f
C8 Vout m1_931_n929# 0.202f
C9 Vn m1_931_n929# 0.205f
C10 m1_931_n929# 0 2.11f
C11 Vp 0 4.01f
C12 Vout 0 0.316f
C13 Vn 0 0.164f
C14 Vin 0 1.03f
.ends

