* NGSPICE file created from th02.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_D7Y3TR a_n63_n101# a_n33_n75# a_n249_n145# a_63_n75#
+ a_n125_n75#
X0 a_63_n75# a_n63_n101# a_n33_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.233 pd=2.12 as=0.124 ps=1.08 w=0.75 l=0.15
X1 a_n33_n75# a_n63_n101# a_n125_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.08 as=0.233 ps=2.12 w=0.75 l=0.15
C0 a_n33_n75# a_n63_n101# 0.0186f
C1 a_63_n75# a_n63_n101# 0.0104f
C2 a_n33_n75# a_n125_n75# 0.113f
C3 a_n33_n75# a_63_n75# 0.113f
C4 a_n63_n101# a_n125_n75# 0.00451f
C5 a_63_n75# a_n249_n145# 0.0963f
C6 a_n33_n75# a_n249_n145# 0.0361f
C7 a_n125_n75# a_n249_n145# 0.105f
C8 a_n63_n101# a_n249_n145# 0.294f
.ends

.subckt sky130_fd_pr__pfet_01v8_2ZD99F w_n349_n261# a_n153_n139# a_n211_n42# a_153_n42#
+ VSUBS
X0 a_153_n42# a_n153_n139# a_n211_n42# w_n349_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.53
C0 a_n211_n42# w_n349_n261# 0.0224f
C1 a_153_n42# w_n349_n261# 0.0224f
C2 a_n211_n42# a_n153_n139# 0.0177f
C3 a_153_n42# a_n153_n139# 0.0177f
C4 a_n211_n42# a_153_n42# 0.0169f
C5 w_n349_n261# a_n153_n139# 0.476f
C6 a_153_n42# VSUBS 0.0518f
C7 a_n211_n42# VSUBS 0.0518f
C8 a_n153_n139# VSUBS 0.506f
C9 w_n349_n261# VSUBS 1.25f
.ends

.subckt sky130_fd_pr__nfet_01v8_2BW22M a_154_n42# a_n154_n130# a_n314_n182# a_n212_n42#
X0 a_154_n42# a_n154_n130# a_n212_n42# a_n314_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.54
C0 a_154_n42# a_n154_n130# 0.0178f
C1 a_154_n42# a_n212_n42# 0.0169f
C2 a_n154_n130# a_n212_n42# 0.0178f
C3 a_154_n42# a_n314_n182# 0.0737f
C4 a_n212_n42# a_n314_n182# 0.0816f
C5 a_n154_n130# a_n314_n182# 0.924f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJP3BL a_15_n150# w_n211_n369# a_n73_n150# a_n33_n247#
+ VSUBS
X0 a_15_n150# a_n33_n247# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.15
C0 a_n73_n150# w_n211_n369# 0.0292f
C1 a_15_n150# w_n211_n369# 0.0292f
C2 a_n73_n150# a_n33_n247# 0.0267f
C3 a_15_n150# a_n33_n247# 0.0267f
C4 a_n73_n150# a_15_n150# 0.242f
C5 w_n211_n369# a_n33_n247# 0.19f
C6 a_15_n150# VSUBS 0.126f
C7 a_n73_n150# VSUBS 0.126f
C8 a_n33_n247# VSUBS 0.146f
C9 w_n211_n369# VSUBS 1.02f
.ends

.subckt sky130_fd_pr__nfet_01v8_LH5FDA a_n150_n130# a_276_n182# a_n208_n42# a_150_n42#
X0 a_150_n42# a_n150_n130# a_n208_n42# a_276_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.5
C0 a_150_n42# a_n150_n130# 0.0176f
C1 a_150_n42# a_n208_n42# 0.0172f
C2 a_n150_n130# a_n208_n42# 0.0176f
C3 a_150_n42# a_276_n182# 0.0815f
C4 a_n208_n42# a_276_n182# 0.0736f
C5 a_n150_n130# a_276_n182# 0.904f
.ends

.subckt th02 Vp Vin V02 Vn
XXM0 Vin Vn Vn m1_983_133# m1_983_133# sky130_fd_pr__nfet_01v8_D7Y3TR
XXM1 Vp Vin m1_571_144# m1_983_133# Vn sky130_fd_pr__pfet_01v8_2ZD99F
XXM2 m1_571_144# Vp Vn Vp sky130_fd_pr__nfet_01v8_2BW22M
XXM3 V02 Vp Vp m1_983_133# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_983_133# Vn V02 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 Vn Vin 0.0263f
C1 m1_983_133# Vin 0.279f
C2 Vp Vn 0.0244f
C3 Vp m1_983_133# 0.346f
C4 m1_571_144# Vin 0.332f
C5 Vp m1_571_144# 0.176f
C6 V02 Vn 0.00239f
C7 V02 m1_983_133# 0.155f
C8 V02 m1_571_144# 0.011f
C9 Vp Vin 0.251f
C10 Vn m1_983_133# 0.216f
C11 V02 Vin 0.00845f
C12 Vn m1_571_144# 0.00115f
C13 m1_571_144# m1_983_133# 0.0183f
C14 Vp V02 0.0906f
C15 Vn 0 0.261f
C16 V02 0 0.354f
C17 Vp 0 3.18f
C18 m1_571_144# 0 0.258f
C19 m1_983_133# 0 1.45f
C20 Vin 0 0.899f
.ends

