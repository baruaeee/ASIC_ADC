magic
tech sky130A
magscale 1 2
timestamp 1702941824
<< checkpaint >>
rect 1294 2099 4236 2180
rect 671 -925 4236 2099
rect 1294 -978 4236 -925
<< error_s >>
rect 1562 1109 1615 1110
rect 1544 1075 1615 1109
rect 1545 1074 1615 1075
rect 1562 1040 1633 1074
rect 552 999 587 1033
rect 1229 1016 1263 1034
rect 553 980 587 999
rect 572 583 587 980
rect 606 946 641 980
rect 606 583 640 946
rect 606 549 621 583
rect 1193 530 1263 1016
rect 1375 1007 1433 1013
rect 1375 973 1387 1007
rect 1375 967 1433 973
rect 1375 613 1433 619
rect 1375 579 1387 613
rect 1375 573 1433 579
rect 1193 494 1246 530
rect 1562 477 1632 1040
rect 1744 972 1802 978
rect 1744 938 1756 972
rect 1744 932 1802 938
rect 1744 560 1802 566
rect 1744 526 1756 560
rect 1744 520 1802 526
rect 1562 441 1615 477
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_X47ZMQ  XM1
timestamp 0
transform 1 0 1773 0 1 749
box -211 -361 211 361
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 0
transform 1 0 2765 0 1 601
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_2YSB4L  XM3
timestamp 0
transform 1 0 2269 0 1 587
box -338 -252 338 252
use sky130_fd_pr__pfet_01v8_WXD9AX  XM7
timestamp 0
transform 1 0 285 0 1 808
box -338 -261 338 261
use sky130_fd_pr__pfet_01v8_WXD9AX  XM9
timestamp 0
transform 1 0 908 0 1 755
box -338 -261 338 261
use sky130_fd_pr__nfet_01v8_Q8HSKG  XM10
timestamp 0
transform 1 0 1404 0 1 793
box -211 -352 211 352
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
