VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
  MACRO oaTaper STRING ;
END PROPERTYDEFINITIONS

MACRO pre_therm
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN pre_therm 0 0 ;
  SIZE 10.785 BY 12.42 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y15
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.32 11.005 8.975 11.695 ;
        RECT 8.715 9.025 8.975 11.695 ;
      LAYER met2 ;
        RECT 8.2 13.335 8.7 13.835 ;
        RECT 8.32 11.35 8.58 13.835 ;
      LAYER via ;
        RECT 8.375 11.435 8.525 11.585 ;
    END
  END Y15
  PIN Y14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 10.455 7.3 10.775 7.56 ;
        RECT 10.455 4.84 10.685 7.56 ;
        RECT 10.025 4.84 10.685 5.53 ;
      LAYER met2 ;
        RECT 11.465 7.18 11.965 7.68 ;
        RECT 10.455 7.3 11.965 7.56 ;
      LAYER via ;
        RECT 10.54 7.355 10.69 7.505 ;
    END
  END Y14
  PIN Y13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.815 5.46 9.135 5.72 ;
        RECT 8.9 4.815 9.13 7.56 ;
        RECT 8.535 4.815 9.13 5.505 ;
      LAYER met2 ;
        RECT 11.465 5.34 11.965 5.84 ;
        RECT 8.815 5.46 11.965 5.72 ;
      LAYER via ;
        RECT 8.9 5.515 9.05 5.665 ;
    END
  END Y13
  PIN Y12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.28 6.97 7.77 7.66 ;
        RECT 7.51 4.76 7.77 7.66 ;
        RECT 7.145 4.765 7.77 5.455 ;
        RECT 7.45 4.76 7.77 5.455 ;
      LAYER met2 ;
        RECT 11.465 4.64 11.965 5.14 ;
        RECT 7.45 4.76 11.965 5.02 ;
      LAYER via ;
        RECT 7.535 4.815 7.685 4.965 ;
    END
  END Y12
  PIN Y11
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.41 10.98 7.225 11.67 ;
        RECT 6.965 9.025 7.225 11.67 ;
      LAYER met2 ;
        RECT 6.29 13.335 6.79 13.835 ;
        RECT 6.41 11.35 6.67 13.835 ;
      LAYER via ;
        RECT 6.465 11.435 6.615 11.585 ;
    END
  END Y11
  PIN Y10
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.735 11.025 5.435 11.715 ;
        RECT 5.175 8.97 5.435 11.715 ;
        RECT 4.685 8.97 5.435 9.66 ;
      LAYER met2 ;
        RECT 4.615 13.335 5.115 13.835 ;
        RECT 4.735 11.395 4.995 13.835 ;
      LAYER via ;
        RECT 4.79 11.48 4.94 11.63 ;
    END
  END Y10
  PIN Y09
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.46 5.83 6.39 6.09 ;
        RECT 5.46 5.83 5.79 6.46 ;
        RECT 5.53 4.89 5.76 6.46 ;
        RECT 5.495 5.83 5.755 6.78 ;
      LAYER met2 ;
        RECT 3.19 7.38 5.755 7.64 ;
        RECT 5.495 6.46 5.755 7.64 ;
        RECT 3.715 13.335 4.215 13.835 ;
        RECT 3.835 12.875 4.095 13.835 ;
        RECT 3.19 12.875 4.095 13.135 ;
        RECT 3.19 7.38 3.45 13.135 ;
      LAYER via ;
        RECT 5.55 6.545 5.7 6.695 ;
    END
  END Y09
  PIN Y08
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.13 4.765 4.46 6.525 ;
        RECT 4.13 4.765 4.39 6.845 ;
        RECT 3.81 4.765 4.46 5.455 ;
      LAYER met2 ;
        RECT 2.73 6.92 4.39 7.18 ;
        RECT 4.13 6.525 4.39 7.18 ;
        RECT 2.73 13.335 3.23 13.835 ;
        RECT 2.73 6.92 2.99 13.835 ;
      LAYER via ;
        RECT 4.185 6.61 4.335 6.76 ;
    END
  END Y08
  PIN Y07
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.27 6.995 2.97 7.685 ;
        RECT 2.74 4.88 2.97 7.685 ;
        RECT 2.17 4.88 2.97 5.21 ;
      LAYER met2 ;
        RECT 0.37 13.02 2.53 13.34 ;
        RECT 2.27 7.365 2.53 13.34 ;
        RECT 0.37 13.02 0.87 13.84 ;
      LAYER via ;
        RECT 2.325 7.45 2.475 7.6 ;
    END
  END Y07
  PIN Y06
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.74 6.9 1.44 7.59 ;
        RECT 1.21 4.83 1.44 7.59 ;
        RECT 0.795 4.83 1.44 5.16 ;
      LAYER met2 ;
        RECT -1.18 7.33 1.06 7.59 ;
        RECT -1.18 7.21 -0.68 7.71 ;
      LAYER via ;
        RECT 0.825 7.385 0.975 7.535 ;
    END
  END Y06
  PIN Y05
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 9.94 2.825 10.71 3.515 ;
        RECT 10.48 0.615 10.71 3.515 ;
        RECT 10.145 0.615 10.71 1.305 ;
      LAYER met2 ;
        RECT 11.465 0.495 11.965 0.995 ;
        RECT 10.39 0.615 11.965 0.875 ;
      LAYER via ;
        RECT 10.475 0.67 10.625 0.82 ;
    END
  END Y05
  PIN Y04
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.495 2.615 9.375 3.305 ;
        RECT 9.145 0.725 9.375 3.305 ;
        RECT 8.81 0.725 9.375 1.415 ;
      LAYER met2 ;
        RECT 8.69 -1.265 9.19 -0.765 ;
        RECT 8.81 -1.265 9.07 1.045 ;
      LAYER via ;
        RECT 8.865 0.81 9.015 0.96 ;
    END
  END Y04
  PIN Y03
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.98 3.07 7.765 3.695 ;
        RECT 7.535 0.615 7.765 3.695 ;
        RECT 7.035 0.615 7.765 1.305 ;
        RECT 6.98 3.045 7.21 3.695 ;
      LAYER met2 ;
        RECT 6.915 -1.265 7.415 -0.765 ;
        RECT 7.035 -1.265 7.295 0.935 ;
      LAYER via ;
        RECT 7.09 0.7 7.24 0.85 ;
    END
  END Y03
  PIN Y02
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.87 2.9 4.615 3.59 ;
        RECT 4.385 0.685 4.615 3.59 ;
        RECT 3.885 0.685 4.615 1.015 ;
      LAYER met2 ;
        RECT 3.765 -1.265 4.265 -0.765 ;
        RECT 3.885 -1.265 4.145 1.005 ;
      LAYER via ;
        RECT 3.94 0.77 4.09 0.92 ;
    END
  END Y02
  PIN Y01
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.58 2.86 3.1 3.55 ;
        RECT 2.875 0.525 3.1 3.55 ;
        RECT 2.6 0.525 3.1 0.855 ;
      LAYER met2 ;
        RECT 2.48 -1.265 2.98 -0.765 ;
        RECT 2.6 -1.265 2.86 0.845 ;
      LAYER via ;
        RECT 2.655 0.61 2.805 0.76 ;
    END
  END Y01
  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
        RECT 9.275 -0.165 10.005 0.165 ;
        RECT 9.05 8.115 9.78 8.445 ;
        RECT 9.275 -0.165 9.605 8.445 ;
      LAYER met1 ;
        RECT 0 -0.2 10.785 0.2 ;
        RECT 3.26 8.08 10.785 8.48 ;
      LAYER met2 ;
        RECT 9.3 -0.185 9.98 0.185 ;
        RECT 9.075 8.095 9.755 8.465 ;
      LAYER via ;
        RECT 9.175 8.205 9.325 8.355 ;
        RECT 9.4 -0.075 9.55 0.075 ;
        RECT 9.495 8.205 9.645 8.355 ;
        RECT 9.72 -0.075 9.87 0.075 ;
      LAYER via2 ;
        RECT 9.115 8.18 9.315 8.38 ;
        RECT 9.34 -0.1 9.54 0.1 ;
        RECT 9.515 8.18 9.715 8.38 ;
        RECT 9.74 -0.1 9.94 0.1 ;
    END
  END VSS
  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 10.055 12.255 10.785 12.585 ;
        RECT 10.455 3.975 10.785 12.585 ;
        RECT 10.055 3.975 10.785 4.305 ;
      LAYER met3 ;
        RECT 10.06 3.95 10.78 4.33 ;
        RECT 10.05 3.975 10.78 4.305 ;
        RECT 10.06 12.23 10.78 12.61 ;
        RECT 10.05 12.255 10.78 12.585 ;
      LAYER met1 ;
        RECT 9.405 3.9 10.785 4.38 ;
        RECT -0.125 3.94 10.785 4.34 ;
        RECT 6.585 3.9 9.345 4.34 ;
        RECT 7.9 3.9 9.28 4.38 ;
        RECT 7.765 3.9 9.28 4.345 ;
        RECT 6.27 3.94 7.65 4.38 ;
        RECT 1.63 3.94 6.02 4.38 ;
        RECT 3.26 3.9 4.64 4.38 ;
        RECT 1.63 3.9 3.01 4.38 ;
        RECT -0.125 3.9 1.38 4.38 ;
        RECT -0.125 0.47 0.245 1.52 ;
        RECT -0.125 0.47 0.075 4.38 ;
        RECT 4.08 12.22 10.785 12.62 ;
        RECT 4.08 12.22 5.46 12.66 ;
      LAYER met2 ;
        RECT 10.075 3.955 10.755 4.325 ;
        RECT 10.075 12.235 10.755 12.605 ;
      LAYER via ;
        RECT 10.23 12.345 10.38 12.495 ;
        RECT 10.23 4.065 10.38 4.215 ;
        RECT 10.55 12.345 10.7 12.495 ;
        RECT 10.55 4.065 10.7 4.215 ;
      LAYER via2 ;
        RECT 10.115 12.32 10.315 12.52 ;
        RECT 10.115 4.04 10.315 4.24 ;
        RECT 10.515 12.32 10.715 12.52 ;
        RECT 10.515 4.04 10.715 4.24 ;
      LAYER via3 ;
        RECT 10.12 12.32 10.32 12.52 ;
        RECT 10.12 4.04 10.32 4.24 ;
        RECT 10.52 12.32 10.72 12.52 ;
        RECT 10.52 4.04 10.72 4.24 ;
    END
  END VDD
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.1 0.805 5.655 1.175 ;
        RECT 4.79 6.02 5.16 6.39 ;
        RECT 4.79 5.825 5.05 6.39 ;
        RECT 3.23 6.35 3.6 6.72 ;
        RECT 1.88 5.775 2.25 6.145 ;
        RECT 0.37 5.775 0.74 6.145 ;
        RECT 0.23 1.855 0.6 2.705 ;
        RECT -0.095 10.615 0.345 11.995 ;
        RECT -0.68 10.615 0.345 10.875 ;
        RECT -0.68 6.145 -0.42 10.875 ;
      LAYER met2 ;
        RECT 4.345 0.855 5.36 1.175 ;
        RECT -1.18 5.885 5.05 6.145 ;
        RECT 0.69 5.825 5.05 6.145 ;
        RECT -0.68 2.445 4.605 2.705 ;
        RECT 4.345 0.855 4.605 2.705 ;
        RECT 3.23 5.825 3.49 6.67 ;
        RECT -0.68 2.445 -0.42 6.465 ;
        RECT -1.18 5.765 -0.42 6.265 ;
      LAYER via ;
        RECT -0.625 6.23 -0.475 6.38 ;
        RECT 0.315 2.5 0.465 2.65 ;
        RECT 0.455 5.94 0.605 6.09 ;
        RECT 1.935 5.91 2.085 6.06 ;
        RECT 3.285 6.435 3.435 6.585 ;
        RECT 4.845 5.91 4.995 6.06 ;
        RECT 5.155 0.94 5.305 1.09 ;
    END
  END IN
  OBS
    LAYER mcon ;
      RECT 10.485 7.28 10.655 7.45 ;
      RECT 10.24 -0.085 10.41 0.085 ;
      RECT 10.24 4.055 10.41 4.225 ;
      RECT 10.24 8.195 10.41 8.365 ;
      RECT 10.175 0.695 10.345 0.865 ;
      RECT 10.175 1.055 10.345 1.225 ;
      RECT 10.055 4.92 10.225 5.09 ;
      RECT 10.055 5.28 10.225 5.45 ;
      RECT 9.97 2.905 10.14 3.075 ;
      RECT 9.97 3.265 10.14 3.435 ;
      RECT 9.84 6.45 10.01 6.62 ;
      RECT 9.83 1.725 10 1.895 ;
      RECT 9.78 -0.085 9.95 0.085 ;
      RECT 9.78 4.055 9.95 4.225 ;
      RECT 9.78 8.195 9.95 8.365 ;
      RECT 8.93 7.28 9.1 7.45 ;
      RECT 8.84 0.805 9.01 0.975 ;
      RECT 8.84 1.165 9.01 1.335 ;
      RECT 8.8 8.195 8.97 8.365 ;
      RECT 8.745 9.105 8.915 9.275 ;
      RECT 8.735 -0.085 8.905 0.085 ;
      RECT 8.735 4.055 8.905 4.225 ;
      RECT 8.565 4.895 8.735 5.065 ;
      RECT 8.565 5.255 8.735 5.425 ;
      RECT 8.525 2.695 8.695 2.865 ;
      RECT 8.525 3.055 8.695 3.225 ;
      RECT 8.39 0.945 8.56 1.115 ;
      RECT 8.36 12.335 8.53 12.505 ;
      RECT 8.35 11.085 8.52 11.255 ;
      RECT 8.35 11.445 8.52 11.615 ;
      RECT 8.345 6.405 8.515 6.575 ;
      RECT 8.34 8.195 8.51 8.365 ;
      RECT 8.275 -0.085 8.445 0.085 ;
      RECT 8.275 4.055 8.445 4.225 ;
      RECT 8.14 9.96 8.31 10.13 ;
      RECT 7.9 8.195 8.07 8.365 ;
      RECT 7.9 12.335 8.07 12.505 ;
      RECT 7.465 4.055 7.635 4.225 ;
      RECT 7.42 8.195 7.59 8.365 ;
      RECT 7.31 7.05 7.48 7.22 ;
      RECT 7.31 7.41 7.48 7.58 ;
      RECT 7.175 4.865 7.345 5.035 ;
      RECT 7.175 5.225 7.345 5.395 ;
      RECT 7.105 -0.085 7.275 0.085 ;
      RECT 7.105 4.055 7.275 4.225 ;
      RECT 7.065 0.695 7.235 0.865 ;
      RECT 7.065 1.055 7.235 1.225 ;
      RECT 7.01 3.105 7.18 3.275 ;
      RECT 7.01 3.465 7.18 3.635 ;
      RECT 6.995 9.105 7.165 9.275 ;
      RECT 6.97 8.195 7.14 8.365 ;
      RECT 6.965 6.01 7.135 6.18 ;
      RECT 6.695 1.785 6.865 1.955 ;
      RECT 6.645 -0.085 6.815 0.085 ;
      RECT 6.645 4.055 6.815 4.225 ;
      RECT 6.61 8.195 6.78 8.365 ;
      RECT 6.61 12.335 6.78 12.505 ;
      RECT 6.44 11.06 6.61 11.23 ;
      RECT 6.44 11.42 6.61 11.59 ;
      RECT 6.17 9.96 6.34 10.13 ;
      RECT 6.15 8.195 6.32 8.365 ;
      RECT 6.15 12.335 6.32 12.505 ;
      RECT 5.935 4.055 6.105 4.225 ;
      RECT 5.79 8.195 5.96 8.365 ;
      RECT 5.56 4.97 5.73 5.14 ;
      RECT 5.54 6.26 5.71 6.43 ;
      RECT 5.475 -0.085 5.645 0.085 ;
      RECT 5.475 4.055 5.645 4.225 ;
      RECT 5.365 0.905 5.535 1.075 ;
      RECT 5.33 8.195 5.5 8.365 ;
      RECT 5.28 1.705 5.45 1.875 ;
      RECT 5.28 2.065 5.45 2.235 ;
      RECT 5.015 -0.085 5.185 0.085 ;
      RECT 5.015 4.055 5.185 4.225 ;
      RECT 4.915 8.195 5.085 8.365 ;
      RECT 4.915 12.335 5.085 12.505 ;
      RECT 4.89 6.12 5.06 6.29 ;
      RECT 4.765 11.105 4.935 11.275 ;
      RECT 4.765 11.465 4.935 11.635 ;
      RECT 4.715 9.05 4.885 9.22 ;
      RECT 4.715 9.41 4.885 9.58 ;
      RECT 4.495 10.055 4.665 10.225 ;
      RECT 4.455 8.195 4.625 8.365 ;
      RECT 4.455 12.335 4.625 12.505 ;
      RECT 4.21 6.325 4.38 6.495 ;
      RECT 4.095 -0.085 4.265 0.085 ;
      RECT 4.095 4.055 4.265 4.225 ;
      RECT 4.095 8.195 4.265 8.365 ;
      RECT 3.915 0.765 4.085 0.935 ;
      RECT 3.9 2.98 4.07 3.15 ;
      RECT 3.9 3.34 4.07 3.51 ;
      RECT 3.84 4.845 4.01 5.015 ;
      RECT 3.84 5.205 4.01 5.375 ;
      RECT 3.635 -0.085 3.805 0.085 ;
      RECT 3.635 1.545 3.805 1.715 ;
      RECT 3.635 4.055 3.805 4.225 ;
      RECT 3.635 8.195 3.805 8.365 ;
      RECT 3.33 6.45 3.5 6.62 ;
      RECT 2.63 0.61 2.8 0.78 ;
      RECT 2.61 2.94 2.78 3.11 ;
      RECT 2.61 3.3 2.78 3.47 ;
      RECT 2.465 -0.085 2.635 0.085 ;
      RECT 2.465 4.055 2.635 4.225 ;
      RECT 2.465 8.195 2.635 8.365 ;
      RECT 2.3 7.075 2.47 7.245 ;
      RECT 2.3 7.435 2.47 7.605 ;
      RECT 2.2 4.96 2.37 5.13 ;
      RECT 2.12 1.545 2.29 1.715 ;
      RECT 2.005 -0.085 2.175 0.085 ;
      RECT 2.005 4.055 2.175 4.225 ;
      RECT 2.005 8.195 2.175 8.365 ;
      RECT 1.98 5.875 2.15 6.045 ;
      RECT 1.265 10.885 1.435 11.055 ;
      RECT 1.015 3.485 1.185 3.655 ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.835 8.195 1.005 8.365 ;
      RECT 0.825 4.91 0.995 5.08 ;
      RECT 0.77 6.98 0.94 7.15 ;
      RECT 0.77 7.34 0.94 7.51 ;
      RECT 0.525 9.405 0.695 9.575 ;
      RECT 0.525 9.765 0.695 9.935 ;
      RECT 0.485 0.55 0.655 0.72 ;
      RECT 0.485 0.91 0.655 1.08 ;
      RECT 0.485 1.27 0.655 1.44 ;
      RECT 0.47 5.875 0.64 6.045 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
      RECT 0.375 8.195 0.545 8.365 ;
      RECT 0.33 2.05 0.5 2.22 ;
      RECT 0.305 8.78 0.475 8.95 ;
      RECT 0.06 10.99 0.23 11.16 ;
      RECT 0.06 11.45 0.23 11.62 ;
      RECT 0.045 0.55 0.215 0.72 ;
      RECT 0.045 0.91 0.215 1.08 ;
      RECT 0.045 1.27 0.215 1.44 ;
    LAYER met1 ;
      RECT 9.73 1.625 9.99 2.005 ;
      RECT 9.73 1.625 10.1 1.995 ;
      RECT 5.255 1.57 5.48 2.47 ;
      RECT 6.595 1.685 6.965 2.325 ;
      RECT 5.25 1.645 5.48 2.295 ;
      RECT 5.25 1.685 6.965 2.005 ;
      RECT 6.07 9.86 6.33 10.275 ;
      RECT 6.07 9.86 6.44 10.23 ;
      RECT 1.185 9.325 1.515 11.085 ;
      RECT 1.185 9.955 4.765 10.325 ;
      RECT 0.495 9.325 1.515 10.015 ;
      RECT 0.275 8.08 0.505 9.01 ;
      RECT 0 8.08 3.01 8.48 ;
      RECT 0.955 0.47 1.245 3.685 ;
      RECT 2.02 1.35 2.39 2.2 ;
      RECT 0.955 1.35 2.39 1.67 ;
      RECT 0.455 0.47 1.245 1.52 ;
      RECT 9.74 6.35 10.11 6.72 ;
      RECT 8.29 0.845 8.66 1.215 ;
      RECT 8.245 6.305 8.615 6.675 ;
      RECT 8.04 9.86 8.41 10.23 ;
      RECT 6.865 5.91 7.235 6.28 ;
      RECT 3.535 1.35 3.905 2.2 ;
    LAYER via ;
      RECT 9.825 6.405 9.975 6.555 ;
      RECT 9.785 1.77 9.935 1.92 ;
      RECT 8.345 0.98 8.495 1.13 ;
      RECT 8.3 6.39 8.45 6.54 ;
      RECT 8.095 9.995 8.245 10.145 ;
      RECT 6.92 6.045 7.07 6.195 ;
      RECT 6.76 1.77 6.91 1.92 ;
      RECT 6.125 10.04 6.275 10.19 ;
      RECT 4.56 10.04 4.71 10.19 ;
      RECT 3.59 1.965 3.74 2.115 ;
      RECT 2.185 1.965 2.335 2.115 ;
    LAYER met2 ;
      RECT 4.505 9.955 6.415 10.275 ;
      RECT 6.155 5.96 6.415 10.275 ;
      RECT 4.505 9.955 8.3 10.23 ;
      RECT 8.04 9.91 8.3 10.23 ;
      RECT 8.245 5.96 8.505 6.625 ;
      RECT 8.245 6.35 10.06 6.61 ;
      RECT 6.155 5.96 8.505 6.28 ;
      RECT 6.705 1.685 9.99 2.005 ;
      RECT 8.29 0.895 8.55 2.005 ;
      RECT 2.13 1.88 3.795 2.2 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END pre_therm

END LIBRARY
