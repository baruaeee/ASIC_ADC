magic
tech sky130A
magscale 1 2
timestamp 1706270854
<< psubdiff >>
rect 1182 -1008 1216 -946
rect 1182 -1041 1254 -1008
rect 1183 -1042 1254 -1041
<< nsubdiff >>
rect 947 22 1005 56
<< locali >>
rect 979 22 1006 56
rect 815 -367 877 -333
rect 843 -589 877 -367
rect 843 -623 1216 -589
rect 1182 -681 1216 -623
rect 1182 -802 1334 -740
rect 1182 -1008 1216 -957
rect 1182 -1039 1254 -1008
rect 1183 -1042 1254 -1039
rect 1440 -1042 1461 -1008
<< viali >>
rect 945 22 979 56
rect 1461 -1042 1495 -1008
<< metal1 >>
rect 924 161 1024 196
rect 587 127 1024 161
rect 587 89 621 127
rect 924 96 1024 127
rect 378 56 430 62
rect 543 55 657 89
rect 944 68 978 96
rect 939 56 985 68
rect 378 -2 430 4
rect 529 -42 657 -3
rect 738 -6 792 56
rect 939 22 945 56
rect 979 22 985 56
rect 939 10 985 22
rect 563 -95 602 -42
rect 563 -134 864 -95
rect 825 -223 864 -134
rect 944 -141 978 10
rect 944 -194 1057 -141
rect 1283 -151 1317 -133
rect 1283 -185 1517 -151
rect 1283 -197 1317 -185
rect 825 -259 934 -223
rect 1115 -259 1227 -257
rect 825 -262 1227 -259
rect 417 -291 716 -290
rect 417 -325 849 -291
rect 895 -296 1227 -262
rect 895 -298 1189 -296
rect 417 -369 451 -325
rect 815 -371 849 -325
rect 509 -396 755 -378
rect 509 -412 595 -396
rect 589 -448 595 -412
rect 647 -412 755 -396
rect 647 -448 653 -412
rect 1150 -468 1189 -298
rect 1483 -344 1517 -185
rect 1472 -444 1572 -344
rect 1150 -507 1385 -468
rect 280 -668 380 -576
rect 1346 -633 1385 -507
rect 280 -676 301 -668
rect 295 -720 301 -676
rect 353 -676 380 -668
rect 353 -720 359 -676
rect 1387 -754 1421 -701
rect 1525 -754 1559 -444
rect 1387 -788 1559 -754
rect 430 -804 464 -796
rect 394 -856 400 -804
rect 452 -856 464 -804
rect 1068 -798 1102 -796
rect 1068 -804 1144 -798
rect 1068 -856 1092 -804
rect 1387 -833 1421 -788
rect 1092 -862 1144 -856
rect 1292 -906 1344 -905
rect 492 -932 1040 -906
rect 492 -940 696 -932
rect 694 -966 696 -940
rect 748 -940 1040 -932
rect 1292 -911 1378 -906
rect 748 -966 756 -940
rect 1344 -940 1378 -911
rect 1292 -969 1344 -963
rect 696 -990 748 -984
rect 1470 -996 1570 -972
rect 1455 -1008 1570 -996
rect 1455 -1042 1461 -1008
rect 1495 -1042 1570 -1008
rect 1455 -1054 1570 -1042
rect 1470 -1072 1570 -1054
<< via1 >>
rect 378 4 430 56
rect 595 -448 647 -396
rect 301 -720 353 -668
rect 400 -856 452 -804
rect 1092 -856 1144 -804
rect 696 -984 748 -932
rect 1292 -963 1344 -911
<< metal2 >>
rect 372 47 378 56
rect 310 13 378 47
rect 310 -662 344 13
rect 372 4 378 13
rect 430 4 436 56
rect 595 -396 647 -390
rect 595 -454 647 -448
rect 604 -611 638 -454
rect 409 -645 638 -611
rect 301 -668 353 -662
rect 301 -726 353 -720
rect 310 -941 344 -726
rect 409 -798 443 -645
rect 400 -804 452 -798
rect 1086 -856 1092 -804
rect 1144 -813 1150 -804
rect 1144 -856 1159 -813
rect 400 -862 452 -856
rect 1125 -920 1159 -856
rect 1286 -920 1292 -911
rect 690 -941 696 -932
rect 310 -975 696 -941
rect 690 -984 696 -975
rect 748 -984 754 -932
rect 1125 -954 1292 -920
rect 1286 -963 1292 -954
rect 1344 -963 1350 -911
use sky130_fd_pr__pfet_01v8_P28Q2U  XM0
timestamp 1706270542
transform 0 -1 632 1 0 -351
box -211 -354 211 354
use sky130_fd_pr__nfet_01v8_ZMY3VB  XM1
timestamp 1706270542
transform -1 0 766 0 1 -826
box -486 -252 486 252
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 1706239161
transform 0 -1 597 1 0 25
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_WV9GCW  XM3
timestamp 1706270542
transform 1 0 1170 0 1 -169
box -296 -261 296 261
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1706270542
transform -1 0 1361 0 -1 -768
box -211 -310 211 310
<< labels >>
flabel metal1 1472 -444 1572 -344 0 FreeSans 256 0 0 0 V12
port 1 nsew
flabel metal1 280 -676 380 -576 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 924 96 1024 196 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 1470 -1072 1570 -972 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
