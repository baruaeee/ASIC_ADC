magic
tech sky130A
magscale 1 2
timestamp 1706529083
<< metal1 >>
rect 1535 6285 1541 6337
rect 1593 6285 1599 6337
rect 1710 4885 1762 4891
rect 1710 4826 1762 4832
rect 4140 2414 4388 2462
<< via1 >>
rect 1541 6285 1593 6337
rect 1710 4832 1762 4885
<< metal2 >>
rect 1434 7053 5555 7106
rect 1434 4885 1487 7053
rect 1543 6950 5278 6997
rect 1543 6343 1590 6950
rect 5231 6651 5278 6950
rect 5502 6793 5555 7053
rect 5502 6740 7595 6793
rect 1541 6337 1593 6343
rect 1541 6279 1593 6285
rect 1434 4832 1710 4885
rect 1762 4832 1768 4885
use therm  therm_0
timestamp 1706527770
transform 1 0 4297 0 1 72
box -111 1962 7123 6724
use Analog  x1
timestamp 1706529083
transform 1 0 0 0 1 7400
box 1538 -6946 5443 -6
<< end >>
