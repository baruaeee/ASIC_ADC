* NGSPICE file created from th01.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_E9WT88 w_n828_n261# a_n632_n139# a_632_n42# a_n690_n42#
+ VSUBS
X0 a_632_n42# a_n632_n139# a_n690_n42# w_n828_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=6.32
C0 a_n632_n139# a_632_n42# 0.0246f
C1 a_632_n42# w_n828_n261# 0.0498f
C2 a_n632_n139# w_n828_n261# 2.08f
C3 a_632_n42# a_n690_n42# 0.0046f
C4 a_n632_n139# a_n690_n42# 0.0246f
C5 a_n690_n42# w_n828_n261# 0.0498f
C6 a_632_n42# VSUBS 0.0373f
C7 a_n690_n42# VSUBS 0.0373f
C8 a_n632_n139# VSUBS 1.65f
C9 w_n828_n261# VSUBS 3.56f
.ends

.subckt sky130_fd_pr__nfet_01v8_JBS6VA a_n73_n632# a_n175_n806# a_15_n632# a_n33_n720#
X0 a_15_n632# a_n33_n720# a_n73_n632# a_n175_n806# sky130_fd_pr__nfet_01v8 ad=1.83 pd=13.2 as=1.83 ps=13.2 w=6.32 l=0.15
C0 a_n73_n632# a_15_n632# 1.01f
C1 a_n73_n632# a_n33_n720# 0.0502f
C2 a_n33_n720# a_15_n632# 0.0502f
C3 a_15_n632# a_n175_n806# 0.671f
C4 a_n73_n632# a_n175_n806# 0.671f
C5 a_n33_n720# a_n175_n806# 0.352f
.ends

.subckt sky130_fd_pr__nfet_01v8_43TXAA a_n658_n42# a_n760_n216# a_n600_n130# a_600_n42#
X0 a_600_n42# a_n600_n130# a_n658_n42# a_n760_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=6
C0 a_n600_n130# a_600_n42# 0.0244f
C1 a_n658_n42# a_n600_n130# 0.0244f
C2 a_n658_n42# a_600_n42# 0.00484f
C3 a_600_n42# a_n760_n216# 0.0875f
C4 a_n658_n42# a_n760_n216# 0.0875f
C5 a_n600_n130# a_n760_n216# 3.46f
.ends

.subckt sky130_fd_pr__pfet_01v8_MGA5QL w_n214_n819# a_n33_n697# a_n76_n600# a_18_n600#
+ VSUBS
X0 a_18_n600# a_n33_n697# a_n76_n600# w_n214_n819# sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.6 as=1.74 ps=12.6 w=6 l=0.18
C0 a_18_n600# a_n76_n600# 0.896f
C1 a_n33_n697# a_n76_n600# 0.0466f
C2 w_n214_n819# a_18_n600# 0.388f
C3 a_n33_n697# w_n214_n819# 0.239f
C4 w_n214_n819# a_n76_n600# 0.388f
C5 a_n33_n697# a_18_n600# 0.0466f
C6 a_18_n600# VSUBS 0.255f
C7 a_n76_n600# VSUBS 0.255f
C8 a_n33_n697# VSUBS 0.125f
C9 w_n214_n819# VSUBS 3.01f
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_FM7VE8 a_n35_n1932# a_n165_n2062# a_n35_1500#
X0 a_n35_1500# a_n35_n1932# a_n165_n2062# sky130_fd_pr__res_xhigh_po_0p35 l=15
C0 a_n35_n1932# a_n165_n2062# 0.598f
C1 a_n35_1500# a_n165_n2062# 0.598f
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_7RFGLT a_n165_n1062# a_n35_500# a_n35_n932#
X0 a_n35_500# a_n35_n932# a_n165_n1062# sky130_fd_pr__res_xhigh_po_0p35 l=5
C0 a_n35_500# a_n35_n932# 0.00382f
C1 a_n35_n932# a_n165_n1062# 0.593f
C2 a_n35_500# a_n165_n1062# 0.593f
.ends

.subckt sky130_fd_pr__nfet_01v8_69TQ3K a_n260_n274# a_100_n100# a_n158_n100# a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n260_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_n100_n188# a_100_n100# 0.0268f
C1 a_n158_n100# a_n100_n188# 0.0268f
C2 a_n158_n100# a_100_n100# 0.0556f
C3 a_100_n100# a_n260_n274# 0.146f
C4 a_n158_n100# a_n260_n274# 0.146f
C5 a_n100_n188# a_n260_n274# 0.724f
.ends

.subckt sky130_fd_pr__pfet_01v8_3HMWVM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
+ VSUBS
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_100_n100# a_n158_n100# 0.0556f
C1 a_n100_n197# a_n158_n100# 0.0268f
C2 w_n296_n319# a_100_n100# 0.0852f
C3 a_n100_n197# w_n296_n319# 0.434f
C4 w_n296_n319# a_n158_n100# 0.0852f
C5 a_n100_n197# a_100_n100# 0.0268f
C6 a_100_n100# VSUBS 0.0607f
C7 a_n158_n100# VSUBS 0.0607f
C8 a_n100_n197# VSUBS 0.311f
C9 w_n296_n319# VSUBS 1.65f
.ends

.subckt sky130_fd_pr__nfet_01v8_PSFW3M a_n88_n100# a_n33_n188# a_n190_n274# a_30_n100#
X0 a_30_n100# a_n33_n188# a_n88_n100# a_n190_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n33_n188# a_30_n100# 0.0111f
C1 a_n88_n100# a_n33_n188# 0.0111f
C2 a_n88_n100# a_30_n100# 0.121f
C3 a_30_n100# a_n190_n274# 0.139f
C4 a_n88_n100# a_n190_n274# 0.139f
C5 a_n33_n188# a_n190_n274# 0.346f
.ends

.subckt op-amp Vp vin Vout m1_2069_183# m1_155_757# m1_924_890# Vn
XXR1 Vout Vn m1_109_n237# sky130_fd_pr__res_xhigh_po_0p35_FM7VE8
XXR2 Vn m1_109_n237# Vn sky130_fd_pr__res_xhigh_po_0p35_7RFGLT
XXR3 Vp Vn m1_n55_181# sky130_fd_pr__res_xhigh_po_0p35_FM7VE8
XXM1 Vn Vn m1_2069_183# m1_1581_69# sky130_fd_pr__nfet_01v8_69TQ3K
XXM2 m1_924_890# m1_109_n237# m1_1581_69# m1_924_890# Vn sky130_fd_pr__pfet_01v8_3HMWVM
XXM3 Vn m1_1581_69# Vn m1_1581_69# sky130_fd_pr__nfet_01v8_69TQ3K
XXM4 m1_924_890# vin m1_924_890# m1_2069_183# Vn sky130_fd_pr__pfet_01v8_3HMWVM
XXM5 Vp m1_155_757# m1_924_890# Vp Vn sky130_fd_pr__pfet_01v8_3HMWVM
XXM6 m1_2069_183# Vp Vn Vout sky130_fd_pr__nfet_01v8_PSFW3M
XXM7 Vp m1_155_757# Vout Vp Vn sky130_fd_pr__pfet_01v8_3HMWVM
XXM9 Vp m1_155_757# m1_155_757# Vp Vn sky130_fd_pr__pfet_01v8_3HMWVM
XXM8 Vn Vout Vn m1_2069_183# sky130_fd_pr__nfet_01v8_69TQ3K
XXM10 Vn m1_155_757# Vn m1_n55_181# sky130_fd_pr__nfet_01v8_69TQ3K
XXM11 Vn Vn m1_n55_181# m1_n55_181# sky130_fd_pr__nfet_01v8_69TQ3K
C0 m1_1581_69# m1_109_n237# 0.118f
C1 Vp m1_924_890# 0.844f
C2 m1_1581_69# m1_n55_181# 0.00446f
C3 m1_1581_69# m1_2069_183# 0.271f
C4 Vp Vout 0.217f
C5 Vp m1_155_757# 0.801f
C6 Vp vin 0.108f
C7 Vp m1_109_n237# 0.0163f
C8 Vout m1_924_890# 0.00373f
C9 Vp m1_n55_181# 0.489f
C10 Vp m1_2069_183# 0.164f
C11 m1_924_890# m1_155_757# 0.429f
C12 m1_924_890# vin 0.243f
C13 Vout m1_155_757# 0.0585f
C14 m1_924_890# m1_109_n237# 0.238f
C15 Vout vin 0.00109f
C16 m1_924_890# m1_n55_181# 8.44e-20
C17 m1_924_890# m1_2069_183# 0.114f
C18 Vout m1_109_n237# 7.8e-20
C19 m1_155_757# vin 0.0746f
C20 m1_1581_69# Vn 0.486f
C21 m1_109_n237# m1_155_757# 0.158f
C22 Vout m1_2069_183# 0.242f
C23 m1_109_n237# vin 0.0127f
C24 m1_155_757# m1_n55_181# 0.334f
C25 m1_155_757# m1_2069_183# 0.123f
C26 vin m1_2069_183# 0.186f
C27 m1_109_n237# m1_n55_181# 0.0477f
C28 m1_109_n237# m1_2069_183# 3.07e-19
C29 Vp Vn 0.969f
C30 m1_924_890# Vn 0.424f
C31 Vp m1_1581_69# 0.00755f
C32 Vout Vn 0.784f
C33 Vn m1_155_757# 0.264f
C34 Vn vin 0.0177f
C35 Vn m1_109_n237# 1.03f
C36 m1_1581_69# m1_924_890# 0.129f
C37 Vn m1_n55_181# 0.537f
C38 Vn m1_2069_183# 0.454f
C39 Vout m1_1581_69# 0.0035f
C40 m1_1581_69# m1_155_757# 0.0687f
C41 m1_1581_69# vin 0.0119f
C42 Vp 0 5.89f
C43 Vn 0 -0.792f
C44 m1_n55_181# 0 2.29f
C45 m1_155_757# 0 1.31f
C46 Vout 0 3.44f
C47 m1_2069_183# 0 1.05f
C48 m1_924_890# 0 2.64f
C49 vin 0 0.256f
C50 m1_1581_69# 0 1.4f
C51 m1_109_n237# 0 1.8f
.ends

.subckt th01 Vp Vin Vout Vn
XXM4 Vp Vin m1_3566_n290# Vp Vn sky130_fd_pr__pfet_01v8_E9WT88
XXM5 Vn Vn m1_3566_n290# Vin sky130_fd_pr__nfet_01v8_JBS6VA
XXM6 Vn Vn m1_3566_n290# Vout sky130_fd_pr__nfet_01v8_43TXAA
XXM7 Vp m1_3566_n290# Vout Vp Vn sky130_fd_pr__pfet_01v8_MGA5QL
Xop-amp_0 Vp op-amp_0/vin Vin op-amp_0/m1_2069_183# op-amp_0/m1_155_757# op-amp_0/m1_924_890#
+ Vn op-amp
C0 op-amp_0/m1_155_757# op-amp_0/m1_2069_183# 7.59e-19
C1 Vout Vn 0.0886f
C2 op-amp_0/m1_2069_183# m1_3566_n290# 8.06e-20
C3 op-amp_0/vin Vin 4.42e-22
C4 Vp Vin 0.682f
C5 Vout Vp 0.13f
C6 Vin op-amp_0/m1_155_757# 0.00409f
C7 Vp Vn 0.429f
C8 Vin m1_3566_n290# 0.195f
C9 Vin op-amp_0/m1_924_890# 3.01e-19
C10 Vout m1_3566_n290# 0.378f
C11 Vp op-amp_0/vin 4.69e-20
C12 Vn op-amp_0/m1_155_757# -0.00372f
C13 Vn m1_3566_n290# 0.173f
C14 Vp op-amp_0/m1_155_757# 0.0762f
C15 Vp m1_3566_n290# 0.325f
C16 Vin op-amp_0/m1_2069_183# -0.00107f
C17 Vp op-amp_0/m1_924_890# 2.09e-20
C18 Vn op-amp_0/m1_2069_183# 0.023f
C19 Vout Vin 1.06e-19
C20 Vp op-amp_0/m1_2069_183# -0.00114f
C21 Vin Vn 0.323f
C22 Vp 0 12.4f
C23 Vn 0 0.174f
C24 op-amp_0/m1_n55_181# 0 2.29f
C25 op-amp_0/m1_155_757# 0 1.31f
C26 Vin 0 4.93f
C27 op-amp_0/m1_2069_183# 0 1.05f
C28 op-amp_0/m1_924_890# 0 2.64f
C29 op-amp_0/vin 0 0.256f
C30 op-amp_0/m1_1581_69# 0 1.4f
C31 op-amp_0/m1_109_n237# 0 1.8f
C32 m1_3566_n290# 0 4.14f
C33 Vout 0 0.535f
.ends

