magic
tech sky130A
magscale 1 2
timestamp 1704305861
<< nwell >>
rect -746 -261 746 261
<< pmos >>
rect -550 -42 550 42
<< pdiff >>
rect -608 30 -550 42
rect -608 -30 -596 30
rect -562 -30 -550 30
rect -608 -42 -550 -30
rect 550 30 608 42
rect 550 -30 562 30
rect 596 -30 608 30
rect 550 -42 608 -30
<< pdiffc >>
rect -596 -30 -562 30
rect 562 -30 596 30
<< nsubdiff >>
rect -710 191 -614 225
rect 614 191 710 225
rect -710 129 -676 191
rect 676 129 710 191
rect -710 -191 -676 -129
rect 676 -191 710 -129
rect -710 -225 -614 -191
rect 614 -225 710 -191
<< nsubdiffcont >>
rect -614 191 614 225
rect -710 -129 -676 129
rect 676 -129 710 129
rect -614 -225 614 -191
<< poly >>
rect -550 123 550 139
rect -550 89 -534 123
rect 534 89 550 123
rect -550 42 550 89
rect -550 -89 550 -42
rect -550 -123 -534 -89
rect 534 -123 550 -89
rect -550 -139 550 -123
<< polycont >>
rect -534 89 534 123
rect -534 -123 534 -89
<< locali >>
rect -710 191 -614 225
rect 614 191 710 225
rect -710 129 -676 191
rect 676 129 710 191
rect -550 89 -534 123
rect 534 89 550 123
rect -596 30 -562 46
rect -596 -46 -562 -30
rect 562 30 596 46
rect 562 -46 596 -30
rect -550 -123 -534 -89
rect 534 -123 550 -89
rect -710 -191 -676 -129
rect 676 -191 710 -129
rect -710 -225 -614 -191
rect 614 -225 710 -191
<< viali >>
rect -534 89 534 123
rect -596 -30 -562 30
rect 562 -30 596 30
rect -534 -123 534 -89
<< metal1 >>
rect -546 123 546 129
rect -546 89 -534 123
rect 534 89 546 123
rect -546 83 546 89
rect -602 30 -556 42
rect -602 -30 -596 30
rect -562 -30 -556 30
rect -602 -42 -556 -30
rect 556 30 602 42
rect 556 -30 562 30
rect 596 -30 602 30
rect 556 -42 602 -30
rect -546 -89 546 -83
rect -546 -123 -534 -89
rect 534 -123 546 -89
rect -546 -129 546 -123
<< properties >>
string FIXED_BBOX -693 -208 693 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 5.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
