magic
tech sky130A
timestamp 1703732895
<< pwell >>
rect -373 -126 373 126
<< nmos >>
rect -275 -21 275 21
<< ndiff >>
rect -304 15 -275 21
rect -304 -15 -298 15
rect -281 -15 -275 15
rect -304 -21 -275 -15
rect 275 15 304 21
rect 275 -15 281 15
rect 298 -15 304 15
rect 275 -21 304 -15
<< ndiffc >>
rect -298 -15 -281 15
rect 281 -15 298 15
<< psubdiff >>
rect -355 91 -307 108
rect 307 91 355 108
rect -355 60 -338 91
rect 338 60 355 91
rect -355 -91 -338 -60
rect 338 -91 355 -60
rect -355 -108 -307 -91
rect 307 -108 355 -91
<< psubdiffcont >>
rect -307 91 307 108
rect -355 -60 -338 60
rect 338 -60 355 60
rect -307 -108 307 -91
<< poly >>
rect -275 57 275 65
rect -275 40 -267 57
rect 267 40 275 57
rect -275 21 275 40
rect -275 -40 275 -21
rect -275 -57 -267 -40
rect 267 -57 275 -40
rect -275 -65 275 -57
<< polycont >>
rect -267 40 267 57
rect -267 -57 267 -40
<< locali >>
rect -355 91 -307 108
rect 307 91 355 108
rect -355 60 -338 91
rect 338 60 355 91
rect -275 40 -267 57
rect 267 40 275 57
rect -298 15 -281 23
rect -298 -23 -281 -15
rect 281 15 298 23
rect 281 -23 298 -15
rect -275 -57 -267 -40
rect 267 -57 275 -40
rect -355 -91 -338 -60
rect 338 -91 355 -60
rect -355 -108 -307 -91
rect 307 -108 355 -91
<< viali >>
rect -267 40 267 57
rect -298 -15 -281 15
rect 281 -15 298 15
rect -267 -57 267 -40
<< metal1 >>
rect -273 57 273 60
rect -273 40 -267 57
rect 267 40 273 57
rect -273 37 273 40
rect -301 15 -278 21
rect -301 -15 -298 15
rect -281 -15 -278 15
rect -301 -21 -278 -15
rect 278 15 301 21
rect 278 -15 281 15
rect 298 -15 301 15
rect 278 -21 301 -15
rect -273 -40 273 -37
rect -273 -57 -267 -40
rect 267 -57 273 -40
rect -273 -60 273 -57
<< properties >>
string FIXED_BBOX -346 -99 346 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 5.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
