magic
tech sky130A
magscale 1 2
timestamp 1703731503
<< error_p >>
rect 666 5637 707 5669
rect 1072 5589 1113 5621
rect 1570 5541 1611 5573
rect 1884 5493 1925 5525
rect 2382 5445 2423 5477
rect 2696 5397 2733 5429
rect 3010 5349 3051 5381
rect 3324 5301 3365 5333
rect 3822 5253 3863 5285
rect 4634 5157 4675 5189
rect 5040 5109 5081 5141
rect 5354 5061 5391 5093
rect 5760 5013 5789 5045
rect 6350 4965 6391 4997
rect 6664 4917 6701 4949
rect 7162 4869 7203 4901
rect 8158 4773 8199 4805
rect 9744 4629 9773 4661
rect 10242 4581 10283 4613
rect 11330 4485 11371 4517
rect 11920 4437 11961 4469
rect 13874 4293 13913 4325
rect 14778 4197 14819 4229
rect 17722 4200 17912 4220
rect 15184 4149 15213 4181
rect 17750 4172 17940 4192
rect 15498 4101 15539 4133
rect 15996 4053 16037 4085
rect 16716 3957 16753 3989
rect 17712 3861 17725 3893
rect 17684 3600 17740 3628
rect 17712 3572 17740 3600
rect 314 2685 355 2717
rect 720 2637 761 2669
rect 1218 2589 1259 2621
rect 1532 2541 1573 2573
rect 2030 2493 2071 2525
rect 2344 2445 2381 2477
rect 2658 2397 2699 2429
rect 2972 2349 3013 2381
rect 3470 2301 3511 2333
rect 4282 2205 4323 2237
rect 4688 2157 4729 2189
rect 5002 2109 5039 2141
rect 5408 2061 5437 2093
rect 5998 2013 6039 2045
rect 6312 1965 6349 1997
rect 6810 1917 6851 1949
rect 7806 1821 7847 1853
rect 9392 1677 9421 1709
rect 9890 1629 9931 1661
rect 10978 1533 11019 1565
rect 11568 1485 11609 1517
rect 13522 1341 13561 1373
rect 14426 1245 14467 1277
rect 14832 1197 14861 1229
rect 15146 1149 15187 1181
rect 15644 1101 15685 1133
rect 16364 1005 16401 1037
rect 17360 909 17373 941
use analog_therm  x1
timestamp 1703731503
transform 1 0 76 0 1 4872
box -76 -4272 17988 2728
<< end >>
