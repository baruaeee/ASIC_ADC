magic
tech sky130A
magscale 1 2
timestamp 1704880472
<< pwell >>
rect 560 -160 594 -114
rect 880 -176 930 -100
<< locali >>
rect 494 392 638 456
rect 672 -334 834 -188
rect 1268 -418 1344 -268
<< metal1 >>
rect 922 681 1122 754
rect 576 647 1167 681
rect 576 453 610 647
rect 922 554 1167 647
rect 1113 525 1167 554
rect 576 391 641 453
rect 855 397 993 447
rect 560 297 827 331
rect 560 218 594 297
rect 452 18 652 218
rect 943 169 993 397
rect 1113 391 1205 525
rect 1368 390 1438 524
rect 1227 281 1341 331
rect 1227 169 1277 281
rect 1402 192 1438 390
rect 943 123 1277 169
rect 732 119 1277 123
rect 732 73 993 119
rect 560 -107 594 18
rect 732 -84 782 73
rect 1148 -94 1184 119
rect 1352 52 1552 192
rect 1304 -8 1552 52
rect 1304 -12 1380 -8
rect 1304 -34 1352 -12
rect 1268 -70 1352 -34
rect 559 -141 621 -107
rect 560 -159 621 -141
rect 560 -160 594 -159
rect 880 -176 930 -100
rect 755 -215 837 -189
rect 755 -221 843 -215
rect 755 -239 851 -221
rect 1148 -238 1218 -94
rect 755 -250 875 -239
rect 1148 -240 1182 -238
rect 755 -302 1058 -250
rect 1265 -302 1343 -269
rect 755 -336 1343 -302
rect 755 -372 1058 -336
rect 858 -450 1058 -372
use sky130_fd_pr__pfet_01v8_9DPZTU  XM2
timestamp 1704877912
transform 1 0 747 0 1 421
box -291 -261 291 261
use sky130_fd_pr__nfet_01v8_586EUA  XM3
timestamp 1704877912
transform 0 -1 755 1 0 -137
box -235 -305 235 305
use sky130_fd_pr__nfet_01v8_PJBF84  XM4
timestamp 1704877912
transform 0 -1 1304 1 0 -168
box -284 -258 284 258
use sky130_fd_pr__pfet_01v8_RVEGTV  XM5
timestamp 1704877912
transform 1 0 1287 0 1 457
box -265 -297 265 297
<< labels >>
flabel metal1 452 18 652 218 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 1352 -8 1552 192 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 858 -450 1058 -250 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 922 554 1122 754 0 FreeSans 256 0 0 0 Vp
port 0 nsew
<< end >>
