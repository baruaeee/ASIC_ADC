magic
tech sky130A
magscale 1 2
timestamp 1706574286
<< viali >>
rect 1777 6273 1811 6307
rect 1961 6273 1995 6307
rect 2237 6273 2271 6307
rect 3249 6273 3283 6307
rect 3801 6273 3835 6307
rect 3433 6205 3467 6239
rect 2145 6137 2179 6171
rect 1501 6069 1535 6103
rect 2421 6069 2455 6103
rect 3065 6069 3099 6103
rect 3985 6069 4019 6103
rect 2605 5865 2639 5899
rect 2329 5797 2363 5831
rect 2513 5729 2547 5763
rect 3893 5729 3927 5763
rect 1409 5661 1443 5695
rect 1777 5661 1811 5695
rect 2421 5661 2455 5695
rect 3065 5661 3099 5695
rect 3341 5661 3375 5695
rect 3985 5661 4019 5695
rect 1961 5593 1995 5627
rect 2789 5593 2823 5627
rect 5181 5593 5215 5627
rect 1593 5525 1627 5559
rect 2053 5525 2087 5559
rect 2145 5525 2179 5559
rect 2697 5525 2731 5559
rect 2881 5525 2915 5559
rect 3249 5525 3283 5559
rect 4353 5525 4387 5559
rect 5457 5525 5491 5559
rect 2237 5321 2271 5355
rect 2513 5321 2547 5355
rect 3249 5321 3283 5355
rect 1777 5253 1811 5287
rect 1869 5253 1903 5287
rect 2605 5253 2639 5287
rect 3701 5253 3735 5287
rect 1501 5185 1535 5219
rect 1659 5185 1693 5219
rect 1961 5185 1995 5219
rect 2145 5185 2179 5219
rect 3893 5185 3927 5219
rect 4041 5185 4075 5219
rect 4169 5185 4203 5219
rect 4261 5185 4295 5219
rect 4358 5185 4392 5219
rect 4629 5185 4663 5219
rect 4813 5185 4847 5219
rect 4905 5185 4939 5219
rect 4997 5185 5031 5219
rect 5181 5185 5215 5219
rect 2396 5117 2430 5151
rect 2881 5117 2915 5151
rect 3157 5117 3191 5151
rect 3709 5049 3743 5083
rect 2973 4981 3007 5015
rect 4537 4981 4571 5015
rect 2053 4777 2087 4811
rect 2237 4777 2271 4811
rect 3249 4777 3283 4811
rect 3617 4777 3651 4811
rect 4537 4777 4571 4811
rect 5457 4777 5491 4811
rect 1593 4709 1627 4743
rect 1685 4709 1719 4743
rect 1409 4573 1443 4607
rect 2329 4573 2363 4607
rect 2513 4573 2547 4607
rect 2605 4573 2639 4607
rect 2789 4573 2823 4607
rect 2881 4573 2915 4607
rect 2973 4573 3007 4607
rect 3157 4573 3191 4607
rect 3525 4573 3559 4607
rect 3617 4573 3651 4607
rect 3801 4573 3835 4607
rect 3959 4573 3993 4607
rect 4261 4573 4295 4607
rect 4445 4573 4479 4607
rect 4537 4573 4571 4607
rect 4629 4573 4663 4607
rect 4077 4505 4111 4539
rect 4169 4505 4203 4539
rect 5181 4505 5215 4539
rect 2053 4437 2087 4471
rect 3065 4437 3099 4471
rect 4905 4437 4939 4471
rect 2973 4233 3007 4267
rect 3433 4233 3467 4267
rect 4353 4233 4387 4267
rect 5181 4233 5215 4267
rect 2881 4165 2915 4199
rect 3709 4165 3743 4199
rect 1409 4097 1443 4131
rect 3065 4097 3099 4131
rect 3617 4097 3651 4131
rect 3801 4097 3835 4131
rect 4261 4097 4295 4131
rect 4997 4097 5031 4131
rect 1685 4029 1719 4063
rect 2697 3961 2731 3995
rect 3985 3961 4019 3995
rect 3249 3893 3283 3927
rect 2053 3689 2087 3723
rect 2237 3689 2271 3723
rect 3617 3689 3651 3723
rect 4537 3689 4571 3723
rect 4721 3689 4755 3723
rect 3249 3621 3283 3655
rect 1869 3553 1903 3587
rect 3985 3553 4019 3587
rect 1685 3485 1719 3519
rect 2053 3485 2087 3519
rect 2605 3485 2639 3519
rect 2973 3485 3007 3519
rect 3065 3485 3099 3519
rect 3525 3485 3559 3519
rect 3617 3485 3651 3519
rect 4077 3485 4111 3519
rect 4445 3485 4479 3519
rect 1777 3417 1811 3451
rect 2697 3417 2731 3451
rect 2789 3417 2823 3451
rect 4353 3417 4387 3451
rect 4689 3417 4723 3451
rect 4905 3417 4939 3451
rect 1593 3349 1627 3383
rect 2421 3349 2455 3383
rect 3801 3349 3835 3383
rect 2145 3145 2179 3179
rect 4445 3145 4479 3179
rect 1777 3077 1811 3111
rect 3065 3077 3099 3111
rect 4169 3077 4203 3111
rect 1961 3009 1995 3043
rect 2513 3009 2547 3043
rect 3525 3009 3559 3043
rect 4813 3009 4847 3043
rect 2421 2941 2455 2975
rect 2881 2941 2915 2975
rect 3341 2941 3375 2975
rect 4721 2941 4755 2975
rect 3801 2873 3835 2907
rect 4353 2873 4387 2907
rect 1501 2805 1535 2839
rect 3525 2805 3559 2839
rect 3709 2805 3743 2839
rect 4169 2805 4203 2839
rect 2237 2601 2271 2635
rect 2881 2601 2915 2635
rect 3525 2601 3559 2635
rect 3985 2601 4019 2635
rect 4813 2601 4847 2635
rect 4997 2601 5031 2635
rect 5273 2601 5307 2635
rect 1593 2533 1627 2567
rect 1409 2397 1443 2431
rect 2053 2397 2087 2431
rect 2697 2397 2731 2431
rect 3341 2397 3375 2431
rect 4169 2397 4203 2431
rect 4629 2397 4663 2431
rect 5181 2397 5215 2431
rect 5457 2397 5491 2431
<< metal1 >>
rect 1104 6554 5888 6576
rect 1104 6502 3410 6554
rect 3462 6502 3474 6554
rect 3526 6502 3538 6554
rect 3590 6502 3602 6554
rect 3654 6502 3666 6554
rect 3718 6502 5888 6554
rect 1104 6480 5888 6502
rect 864 6372 1064 6458
rect 3234 6400 3240 6452
rect 3292 6400 3298 6452
rect 3252 6372 3280 6400
rect 864 6344 1992 6372
rect 3252 6344 3832 6372
rect 864 6338 1064 6344
rect 798 6236 998 6284
rect 1762 6264 1768 6316
rect 1820 6264 1826 6316
rect 1964 6313 1992 6344
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6304 3295 6307
rect 3326 6304 3332 6316
rect 3283 6276 3332 6304
rect 3283 6273 3295 6276
rect 3237 6267 3295 6273
rect 2240 6236 2268 6267
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 3804 6313 3832 6344
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 798 6208 2268 6236
rect 798 6164 998 6208
rect 3142 6196 3148 6248
rect 3200 6236 3206 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3200 6208 3433 6236
rect 3200 6196 3206 6208
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3421 6199 3479 6205
rect 2133 6171 2191 6177
rect 2133 6137 2145 6171
rect 2179 6168 2191 6171
rect 3878 6168 3884 6180
rect 2179 6140 3884 6168
rect 2179 6137 2191 6140
rect 2133 6131 2191 6137
rect 3878 6128 3884 6140
rect 3936 6128 3942 6180
rect 1486 6060 1492 6112
rect 1544 6060 1550 6112
rect 2406 6060 2412 6112
rect 2464 6060 2470 6112
rect 3053 6103 3111 6109
rect 3053 6069 3065 6103
rect 3099 6100 3111 6103
rect 3234 6100 3240 6112
rect 3099 6072 3240 6100
rect 3099 6069 3111 6072
rect 3053 6063 3111 6069
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 3973 6103 4031 6109
rect 3973 6100 3985 6103
rect 3844 6072 3985 6100
rect 3844 6060 3850 6072
rect 3973 6069 3985 6072
rect 4019 6100 4031 6103
rect 4614 6100 4620 6112
rect 4019 6072 4620 6100
rect 4019 6069 4031 6072
rect 3973 6063 4031 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 1104 6010 5888 6032
rect 1104 5958 2750 6010
rect 2802 5958 2814 6010
rect 2866 5958 2878 6010
rect 2930 5958 2942 6010
rect 2994 5958 3006 6010
rect 3058 5958 5888 6010
rect 1104 5936 5888 5958
rect 1670 5856 1676 5908
rect 1728 5896 1734 5908
rect 2222 5896 2228 5908
rect 1728 5868 2228 5896
rect 1728 5856 1734 5868
rect 2222 5856 2228 5868
rect 2280 5896 2286 5908
rect 2593 5899 2651 5905
rect 2593 5896 2605 5899
rect 2280 5868 2605 5896
rect 2280 5856 2286 5868
rect 2593 5865 2605 5868
rect 2639 5865 2651 5899
rect 2593 5859 2651 5865
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 3142 5896 3148 5908
rect 3016 5868 3148 5896
rect 3016 5856 3022 5868
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 2317 5831 2375 5837
rect 2317 5797 2329 5831
rect 2363 5828 2375 5831
rect 3050 5828 3056 5840
rect 2363 5800 3056 5828
rect 2363 5797 2375 5800
rect 2317 5791 2375 5797
rect 3050 5788 3056 5800
rect 3108 5788 3114 5840
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 2501 5763 2559 5769
rect 2501 5760 2513 5763
rect 1912 5732 2513 5760
rect 1912 5720 1918 5732
rect 2501 5729 2513 5732
rect 2547 5729 2559 5763
rect 2501 5723 2559 5729
rect 3878 5720 3884 5772
rect 3936 5720 3942 5772
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5692 1823 5695
rect 2038 5692 2044 5704
rect 1811 5664 2044 5692
rect 1811 5661 1823 5664
rect 1765 5655 1823 5661
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 1780 5556 1808 5655
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2130 5652 2136 5704
rect 2188 5692 2194 5704
rect 2406 5702 2412 5704
rect 2399 5692 2412 5702
rect 2188 5664 2412 5692
rect 2188 5652 2194 5664
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 2700 5664 3065 5692
rect 1949 5627 2007 5633
rect 1949 5593 1961 5627
rect 1995 5624 2007 5627
rect 2148 5624 2176 5652
rect 2700 5624 2728 5664
rect 3053 5661 3065 5664
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 3329 5695 3387 5701
rect 3329 5661 3341 5695
rect 3375 5661 3387 5695
rect 3329 5655 3387 5661
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 4019 5664 4200 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 1995 5596 2176 5624
rect 2516 5596 2728 5624
rect 1995 5593 2007 5596
rect 1949 5587 2007 5593
rect 1627 5528 1808 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 1854 5516 1860 5568
rect 1912 5556 1918 5568
rect 2041 5559 2099 5565
rect 2041 5556 2053 5559
rect 1912 5528 2053 5556
rect 1912 5516 1918 5528
rect 2041 5525 2053 5528
rect 2087 5525 2099 5559
rect 2041 5519 2099 5525
rect 2133 5559 2191 5565
rect 2133 5525 2145 5559
rect 2179 5556 2191 5559
rect 2222 5556 2228 5568
rect 2179 5528 2228 5556
rect 2179 5525 2191 5528
rect 2133 5519 2191 5525
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 2314 5516 2320 5568
rect 2372 5556 2378 5568
rect 2516 5556 2544 5596
rect 2774 5584 2780 5636
rect 2832 5584 2838 5636
rect 3344 5624 3372 5655
rect 4062 5624 4068 5636
rect 3344 5596 4068 5624
rect 4062 5584 4068 5596
rect 4120 5584 4126 5636
rect 2372 5528 2544 5556
rect 2372 5516 2378 5528
rect 2590 5516 2596 5568
rect 2648 5556 2654 5568
rect 2685 5559 2743 5565
rect 2685 5556 2697 5559
rect 2648 5528 2697 5556
rect 2648 5516 2654 5528
rect 2685 5525 2697 5528
rect 2731 5525 2743 5559
rect 2685 5519 2743 5525
rect 2869 5559 2927 5565
rect 2869 5525 2881 5559
rect 2915 5556 2927 5559
rect 3142 5556 3148 5568
rect 2915 5528 3148 5556
rect 2915 5525 2927 5528
rect 2869 5519 2927 5525
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 3970 5556 3976 5568
rect 3283 5528 3976 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 3970 5516 3976 5528
rect 4028 5556 4034 5568
rect 4172 5556 4200 5664
rect 5166 5584 5172 5636
rect 5224 5584 5230 5636
rect 4028 5528 4200 5556
rect 4341 5559 4399 5565
rect 4028 5516 4034 5528
rect 4341 5525 4353 5559
rect 4387 5556 4399 5559
rect 4522 5556 4528 5568
rect 4387 5528 4528 5556
rect 4387 5525 4399 5528
rect 4341 5519 4399 5525
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 5442 5516 5448 5568
rect 5500 5516 5506 5568
rect 1104 5466 5888 5488
rect 1104 5414 3410 5466
rect 3462 5414 3474 5466
rect 3526 5414 3538 5466
rect 3590 5414 3602 5466
rect 3654 5414 3666 5466
rect 3718 5414 5888 5466
rect 1104 5392 5888 5414
rect 1670 5352 1676 5364
rect 1504 5324 1676 5352
rect 1504 5225 1532 5324
rect 1670 5312 1676 5324
rect 1728 5312 1734 5364
rect 2038 5352 2044 5364
rect 1780 5324 2044 5352
rect 1780 5293 1808 5324
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 2225 5355 2283 5361
rect 2225 5321 2237 5355
rect 2271 5352 2283 5355
rect 2314 5352 2320 5364
rect 2271 5324 2320 5352
rect 2271 5321 2283 5324
rect 2225 5315 2283 5321
rect 2314 5312 2320 5324
rect 2372 5312 2378 5364
rect 2501 5355 2559 5361
rect 2501 5321 2513 5355
rect 2547 5352 2559 5355
rect 2866 5352 2872 5364
rect 2547 5324 2872 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 3234 5312 3240 5364
rect 3292 5312 3298 5364
rect 3878 5352 3884 5364
rect 3620 5324 3884 5352
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5253 1823 5287
rect 1765 5247 1823 5253
rect 1857 5287 1915 5293
rect 1857 5253 1869 5287
rect 1903 5284 1915 5287
rect 2406 5284 2412 5296
rect 1903 5256 2412 5284
rect 1903 5253 1915 5256
rect 1857 5247 1915 5253
rect 2406 5244 2412 5256
rect 2464 5244 2470 5296
rect 2593 5287 2651 5293
rect 2593 5253 2605 5287
rect 2639 5284 2651 5287
rect 2958 5284 2964 5296
rect 2639 5256 2964 5284
rect 2639 5253 2651 5256
rect 2593 5247 2651 5253
rect 2958 5244 2964 5256
rect 3016 5284 3022 5296
rect 3510 5284 3516 5296
rect 3016 5256 3516 5284
rect 3016 5244 3022 5256
rect 3510 5244 3516 5256
rect 3568 5244 3574 5296
rect 3620 5284 3648 5324
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 4120 5324 4568 5352
rect 4120 5312 4126 5324
rect 3689 5287 3747 5293
rect 3689 5284 3701 5287
rect 3620 5256 3701 5284
rect 3689 5253 3701 5256
rect 3735 5253 3747 5287
rect 4540 5284 4568 5324
rect 3689 5247 3747 5253
rect 4080 5256 4476 5284
rect 4540 5256 5212 5284
rect 1489 5219 1547 5225
rect 1489 5185 1501 5219
rect 1535 5185 1547 5219
rect 1489 5179 1547 5185
rect 1647 5219 1705 5225
rect 1647 5185 1659 5219
rect 1693 5216 1705 5219
rect 1693 5188 1900 5216
rect 1693 5185 1705 5188
rect 1647 5179 1705 5185
rect 1872 5080 1900 5188
rect 1946 5176 1952 5228
rect 2004 5176 2010 5228
rect 4080 5225 4108 5256
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 3881 5219 3939 5225
rect 3881 5216 3893 5219
rect 2179 5188 3893 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 3881 5185 3893 5188
rect 3927 5185 3939 5219
rect 3881 5179 3939 5185
rect 4029 5219 4108 5225
rect 4029 5185 4041 5219
rect 4075 5188 4108 5219
rect 4075 5185 4087 5188
rect 4029 5179 4087 5185
rect 4154 5176 4160 5228
rect 4212 5176 4218 5228
rect 4246 5176 4252 5228
rect 4304 5176 4310 5228
rect 4338 5176 4344 5228
rect 4396 5225 4402 5228
rect 4396 5179 4404 5225
rect 4448 5216 4476 5256
rect 4522 5216 4528 5228
rect 4448 5188 4528 5216
rect 4396 5176 4402 5179
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 4614 5176 4620 5228
rect 4672 5176 4678 5228
rect 4798 5176 4804 5228
rect 4856 5176 4862 5228
rect 4890 5176 4896 5228
rect 4948 5176 4954 5228
rect 5184 5225 5212 5256
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 2222 5108 2228 5160
rect 2280 5148 2286 5160
rect 2384 5151 2442 5157
rect 2384 5148 2396 5151
rect 2280 5120 2396 5148
rect 2280 5108 2286 5120
rect 2384 5117 2396 5120
rect 2430 5117 2442 5151
rect 2384 5111 2442 5117
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 2869 5151 2927 5157
rect 2869 5148 2881 5151
rect 2832 5120 2881 5148
rect 2832 5108 2838 5120
rect 2869 5117 2881 5120
rect 2915 5117 2927 5151
rect 2869 5111 2927 5117
rect 2884 5080 2912 5111
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 3145 5151 3203 5157
rect 3145 5148 3157 5151
rect 3108 5120 3157 5148
rect 3108 5108 3114 5120
rect 3145 5117 3157 5120
rect 3191 5148 3203 5151
rect 5000 5148 5028 5179
rect 3191 5120 5028 5148
rect 3191 5117 3203 5120
rect 3145 5111 3203 5117
rect 3326 5080 3332 5092
rect 1872 5052 2360 5080
rect 2884 5052 3332 5080
rect 2332 5024 2360 5052
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 3697 5083 3755 5089
rect 3697 5049 3709 5083
rect 3743 5080 3755 5083
rect 3970 5080 3976 5092
rect 3743 5052 3976 5080
rect 3743 5049 3755 5052
rect 3697 5043 3755 5049
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 5166 5040 5172 5092
rect 5224 5040 5230 5092
rect 2314 4972 2320 5024
rect 2372 4972 2378 5024
rect 2961 5015 3019 5021
rect 2961 4981 2973 5015
rect 3007 5012 3019 5015
rect 4154 5012 4160 5024
rect 3007 4984 4160 5012
rect 3007 4981 3019 4984
rect 2961 4975 3019 4981
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 4525 5015 4583 5021
rect 4525 4981 4537 5015
rect 4571 5012 4583 5015
rect 5184 5012 5212 5040
rect 4571 4984 5212 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 1104 4922 5888 4944
rect 1104 4870 2750 4922
rect 2802 4870 2814 4922
rect 2866 4870 2878 4922
rect 2930 4870 2942 4922
rect 2994 4870 3006 4922
rect 3058 4870 5888 4922
rect 1104 4848 5888 4870
rect 1946 4768 1952 4820
rect 2004 4768 2010 4820
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4808 2099 4811
rect 2130 4808 2136 4820
rect 2087 4780 2136 4808
rect 2087 4777 2099 4780
rect 2041 4771 2099 4777
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 2222 4768 2228 4820
rect 2280 4768 2286 4820
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 3237 4811 3295 4817
rect 3237 4777 3249 4811
rect 3283 4808 3295 4811
rect 3326 4808 3332 4820
rect 3283 4780 3332 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 1673 4743 1731 4749
rect 1673 4740 1685 4743
rect 1627 4712 1685 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 1673 4709 1685 4712
rect 1719 4740 1731 4743
rect 1854 4740 1860 4752
rect 1719 4712 1860 4740
rect 1719 4709 1731 4712
rect 1673 4703 1731 4709
rect 1854 4700 1860 4712
rect 1912 4700 1918 4752
rect 1964 4740 1992 4768
rect 3050 4740 3056 4752
rect 1964 4712 3056 4740
rect 844 4604 1044 4668
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 844 4576 1409 4604
rect 844 4548 1044 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 1762 4564 1768 4616
rect 1820 4604 1826 4616
rect 2516 4613 2544 4712
rect 3050 4700 3056 4712
rect 3108 4700 3114 4752
rect 3160 4672 3188 4768
rect 2792 4644 3188 4672
rect 2317 4607 2375 4613
rect 2317 4604 2329 4607
rect 1820 4576 2329 4604
rect 1820 4564 1826 4576
rect 2317 4573 2329 4576
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4573 2559 4607
rect 2501 4567 2559 4573
rect 2590 4564 2596 4616
rect 2648 4564 2654 4616
rect 2792 4613 2820 4644
rect 3068 4616 3096 4644
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 2884 4536 2912 4567
rect 2958 4564 2964 4616
rect 3016 4564 3022 4616
rect 3050 4564 3056 4616
rect 3108 4564 3114 4616
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4604 3203 4607
rect 3252 4604 3280 4771
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 3602 4768 3608 4820
rect 3660 4768 3666 4820
rect 4154 4808 4160 4820
rect 3704 4780 4160 4808
rect 3704 4672 3732 4780
rect 4154 4768 4160 4780
rect 4212 4808 4218 4820
rect 4525 4811 4583 4817
rect 4525 4808 4537 4811
rect 4212 4780 4537 4808
rect 4212 4768 4218 4780
rect 4525 4777 4537 4780
rect 4571 4777 4583 4811
rect 4525 4771 4583 4777
rect 5442 4768 5448 4820
rect 5500 4768 5506 4820
rect 3191 4576 3280 4604
rect 3436 4644 3732 4672
rect 3191 4573 3203 4576
rect 3145 4567 3203 4573
rect 3436 4536 3464 4644
rect 4154 4632 4160 4684
rect 4212 4632 4218 4684
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4604 3663 4607
rect 3694 4604 3700 4616
rect 3651 4576 3700 4604
rect 3651 4573 3663 4576
rect 3605 4567 3663 4573
rect 2884 4508 3464 4536
rect 3528 4536 3556 4567
rect 3694 4564 3700 4576
rect 3752 4564 3758 4616
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 3970 4613 3976 4616
rect 3947 4607 3976 4613
rect 3947 4573 3959 4607
rect 3947 4567 3976 4573
rect 3970 4564 3976 4567
rect 4028 4564 4034 4616
rect 4172 4604 4200 4632
rect 4080 4576 4200 4604
rect 3804 4536 3832 4564
rect 4080 4545 4108 4576
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 4479 4576 4537 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4614 4564 4620 4616
rect 4672 4564 4678 4616
rect 3528 4508 3832 4536
rect 4065 4539 4123 4545
rect 4065 4505 4077 4539
rect 4111 4505 4123 4539
rect 4065 4499 4123 4505
rect 2038 4428 2044 4480
rect 2096 4428 2102 4480
rect 2314 4428 2320 4480
rect 2372 4468 2378 4480
rect 3053 4471 3111 4477
rect 3053 4468 3065 4471
rect 2372 4440 3065 4468
rect 2372 4428 2378 4440
rect 3053 4437 3065 4440
rect 3099 4468 3111 4471
rect 4080 4468 4108 4499
rect 4154 4496 4160 4548
rect 4212 4536 4218 4548
rect 4798 4536 4804 4548
rect 4212 4508 4804 4536
rect 4212 4496 4218 4508
rect 4798 4496 4804 4508
rect 4856 4496 4862 4548
rect 5166 4496 5172 4548
rect 5224 4496 5230 4548
rect 4706 4468 4712 4480
rect 3099 4440 4712 4468
rect 3099 4437 3111 4440
rect 3053 4431 3111 4437
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 4890 4428 4896 4480
rect 4948 4428 4954 4480
rect 1104 4378 5888 4400
rect 1104 4326 3410 4378
rect 3462 4326 3474 4378
rect 3526 4326 3538 4378
rect 3590 4326 3602 4378
rect 3654 4326 3666 4378
rect 3718 4326 5888 4378
rect 1104 4304 5888 4326
rect 2961 4267 3019 4273
rect 2961 4233 2973 4267
rect 3007 4264 3019 4267
rect 3050 4264 3056 4276
rect 3007 4236 3056 4264
rect 3007 4233 3019 4236
rect 2961 4227 3019 4233
rect 3050 4224 3056 4236
rect 3108 4224 3114 4276
rect 3418 4224 3424 4276
rect 3476 4224 3482 4276
rect 3786 4264 3792 4276
rect 3620 4236 3792 4264
rect 2869 4199 2927 4205
rect 2869 4165 2881 4199
rect 2915 4196 2927 4199
rect 3142 4196 3148 4208
rect 2915 4168 3148 4196
rect 2915 4165 2927 4168
rect 2869 4159 2927 4165
rect 3142 4156 3148 4168
rect 3200 4156 3206 4208
rect 3620 4196 3648 4236
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 4341 4267 4399 4273
rect 4341 4264 4353 4267
rect 4304 4236 4353 4264
rect 4304 4224 4310 4236
rect 4341 4233 4353 4236
rect 4387 4233 4399 4267
rect 4341 4227 4399 4233
rect 4890 4224 4896 4276
rect 4948 4224 4954 4276
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 3252 4168 3648 4196
rect 3697 4199 3755 4205
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 2222 4088 2228 4140
rect 2280 4128 2286 4140
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2280 4100 3065 4128
rect 2280 4088 2286 4100
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4060 1731 4063
rect 3252 4060 3280 4168
rect 3697 4165 3709 4199
rect 3743 4196 3755 4199
rect 3743 4168 4016 4196
rect 3743 4165 3755 4168
rect 3697 4159 3755 4165
rect 3988 4140 4016 4168
rect 3510 4128 3516 4140
rect 1719 4032 3280 4060
rect 3344 4100 3516 4128
rect 1719 4029 1731 4032
rect 1673 4023 1731 4029
rect 2406 3952 2412 4004
rect 2464 3992 2470 4004
rect 2685 3995 2743 4001
rect 2685 3992 2697 3995
rect 2464 3964 2697 3992
rect 2464 3952 2470 3964
rect 2685 3961 2697 3964
rect 2731 3961 2743 3995
rect 2685 3955 2743 3961
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3924 3295 3927
rect 3344 3924 3372 4100
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 3602 4088 3608 4140
rect 3660 4088 3666 4140
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4097 3847 4131
rect 3789 4091 3847 4097
rect 3804 4060 3832 4091
rect 3970 4088 3976 4140
rect 4028 4088 4034 4140
rect 4154 4088 4160 4140
rect 4212 4088 4218 4140
rect 4246 4088 4252 4140
rect 4304 4088 4310 4140
rect 4908 4128 4936 4224
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4908 4100 4997 4128
rect 4985 4097 4997 4100
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 4172 4060 4200 4088
rect 3804 4032 4200 4060
rect 3510 3952 3516 4004
rect 3568 3992 3574 4004
rect 3973 3995 4031 4001
rect 3973 3992 3985 3995
rect 3568 3964 3985 3992
rect 3568 3952 3574 3964
rect 3973 3961 3985 3964
rect 4019 3992 4031 3995
rect 4019 3964 4936 3992
rect 4019 3961 4031 3964
rect 3973 3955 4031 3961
rect 4908 3936 4936 3964
rect 3283 3896 3372 3924
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 4614 3924 4620 3936
rect 3844 3896 4620 3924
rect 3844 3884 3850 3896
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4890 3884 4896 3936
rect 4948 3884 4954 3936
rect 1104 3834 5888 3856
rect 1104 3782 2750 3834
rect 2802 3782 2814 3834
rect 2866 3782 2878 3834
rect 2930 3782 2942 3834
rect 2994 3782 3006 3834
rect 3058 3782 5888 3834
rect 1104 3760 5888 3782
rect 2041 3723 2099 3729
rect 2041 3689 2053 3723
rect 2087 3720 2099 3723
rect 2130 3720 2136 3732
rect 2087 3692 2136 3720
rect 2087 3689 2099 3692
rect 2041 3683 2099 3689
rect 2130 3680 2136 3692
rect 2188 3680 2194 3732
rect 2225 3723 2283 3729
rect 2225 3689 2237 3723
rect 2271 3720 2283 3723
rect 2498 3720 2504 3732
rect 2271 3692 2504 3720
rect 2271 3689 2283 3692
rect 2225 3683 2283 3689
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 3605 3723 3663 3729
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 3970 3720 3976 3732
rect 3651 3692 3976 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 4246 3680 4252 3732
rect 4304 3680 4310 3732
rect 4338 3680 4344 3732
rect 4396 3680 4402 3732
rect 4525 3723 4583 3729
rect 4525 3689 4537 3723
rect 4571 3720 4583 3723
rect 4614 3720 4620 3732
rect 4571 3692 4620 3720
rect 4571 3689 4583 3692
rect 4525 3683 4583 3689
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 4706 3680 4712 3732
rect 4764 3680 4770 3732
rect 2958 3612 2964 3664
rect 3016 3652 3022 3664
rect 3237 3655 3295 3661
rect 3237 3652 3249 3655
rect 3016 3624 3249 3652
rect 3016 3612 3022 3624
rect 3237 3621 3249 3624
rect 3283 3652 3295 3655
rect 4264 3652 4292 3680
rect 3283 3624 4292 3652
rect 3283 3621 3295 3624
rect 3237 3615 3295 3621
rect 1854 3544 1860 3596
rect 1912 3544 1918 3596
rect 3878 3584 3884 3596
rect 1964 3556 3884 3584
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 1964 3516 1992 3556
rect 3878 3544 3884 3556
rect 3936 3584 3942 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 3936 3556 3985 3584
rect 3936 3544 3942 3556
rect 3973 3553 3985 3556
rect 4019 3553 4031 3587
rect 3973 3547 4031 3553
rect 1719 3488 1992 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 2038 3476 2044 3528
rect 2096 3476 2102 3528
rect 2593 3519 2651 3525
rect 2593 3516 2605 3519
rect 2148 3488 2605 3516
rect 1762 3408 1768 3460
rect 1820 3408 1826 3460
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 2148 3380 2176 3488
rect 2593 3485 2605 3488
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3485 3019 3519
rect 2961 3479 3019 3485
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 3099 3488 3464 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 2314 3408 2320 3460
rect 2372 3448 2378 3460
rect 2685 3451 2743 3457
rect 2685 3448 2697 3451
rect 2372 3420 2697 3448
rect 2372 3408 2378 3420
rect 2685 3417 2697 3420
rect 2731 3417 2743 3451
rect 2685 3411 2743 3417
rect 2777 3451 2835 3457
rect 2777 3417 2789 3451
rect 2823 3417 2835 3451
rect 2976 3448 3004 3479
rect 3234 3448 3240 3460
rect 2976 3420 3240 3448
rect 2777 3411 2835 3417
rect 1627 3352 2176 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 2406 3340 2412 3392
rect 2464 3340 2470 3392
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 2792 3380 2820 3411
rect 3234 3408 3240 3420
rect 3292 3408 3298 3460
rect 3436 3448 3464 3488
rect 3510 3476 3516 3528
rect 3568 3476 3574 3528
rect 3602 3476 3608 3528
rect 3660 3476 3666 3528
rect 3786 3476 3792 3528
rect 3844 3476 3850 3528
rect 4062 3476 4068 3528
rect 4120 3476 4126 3528
rect 4356 3516 4384 3680
rect 4172 3488 4384 3516
rect 4433 3519 4491 3525
rect 3804 3448 3832 3476
rect 3436 3420 3832 3448
rect 2556 3352 2820 3380
rect 3789 3383 3847 3389
rect 2556 3340 2562 3352
rect 3789 3349 3801 3383
rect 3835 3380 3847 3383
rect 4172 3380 4200 3488
rect 4433 3485 4445 3519
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 4338 3408 4344 3460
rect 4396 3408 4402 3460
rect 4448 3448 4476 3479
rect 4677 3451 4735 3457
rect 4677 3448 4689 3451
rect 4448 3420 4689 3448
rect 4448 3392 4476 3420
rect 4677 3417 4689 3420
rect 4723 3417 4735 3451
rect 4677 3411 4735 3417
rect 4890 3408 4896 3460
rect 4948 3408 4954 3460
rect 3835 3352 4200 3380
rect 3835 3349 3847 3352
rect 3789 3343 3847 3349
rect 4430 3340 4436 3392
rect 4488 3340 4494 3392
rect 1104 3290 5888 3312
rect 1104 3238 3410 3290
rect 3462 3238 3474 3290
rect 3526 3238 3538 3290
rect 3590 3238 3602 3290
rect 3654 3238 3666 3290
rect 3718 3238 5888 3290
rect 1104 3216 5888 3238
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 1728 3148 2145 3176
rect 1728 3136 1734 3148
rect 2133 3145 2145 3148
rect 2179 3145 2191 3179
rect 2133 3139 2191 3145
rect 2406 3136 2412 3188
rect 2464 3136 2470 3188
rect 4062 3176 4068 3188
rect 2976 3148 4068 3176
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3108 1823 3111
rect 2424 3108 2452 3136
rect 1811 3080 2452 3108
rect 1811 3077 1823 3080
rect 784 3040 984 3074
rect 1765 3071 1823 3077
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 784 3012 1961 3040
rect 784 2974 984 3012
rect 1949 3009 1961 3012
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2498 3000 2504 3052
rect 2556 3000 2562 3052
rect 2222 2932 2228 2984
rect 2280 2972 2286 2984
rect 2409 2975 2467 2981
rect 2409 2972 2421 2975
rect 2280 2944 2421 2972
rect 2280 2932 2286 2944
rect 2409 2941 2421 2944
rect 2455 2972 2467 2975
rect 2590 2972 2596 2984
rect 2455 2944 2596 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 2590 2932 2596 2944
rect 2648 2932 2654 2984
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 2976 2972 3004 3148
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4338 3136 4344 3188
rect 4396 3176 4402 3188
rect 4433 3179 4491 3185
rect 4433 3176 4445 3179
rect 4396 3148 4445 3176
rect 4396 3136 4402 3148
rect 4433 3145 4445 3148
rect 4479 3145 4491 3179
rect 4433 3139 4491 3145
rect 3053 3111 3111 3117
rect 3053 3077 3065 3111
rect 3099 3108 3111 3111
rect 3142 3108 3148 3120
rect 3099 3080 3148 3108
rect 3099 3077 3111 3080
rect 3053 3071 3111 3077
rect 3142 3068 3148 3080
rect 3200 3068 3206 3120
rect 3326 3068 3332 3120
rect 3384 3068 3390 3120
rect 3602 3068 3608 3120
rect 3660 3108 3666 3120
rect 4154 3108 4160 3120
rect 3660 3080 4160 3108
rect 3660 3068 3666 3080
rect 4154 3068 4160 3080
rect 4212 3108 4218 3120
rect 4982 3108 4988 3120
rect 4212 3080 4988 3108
rect 4212 3068 4218 3080
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 3344 3040 3372 3068
rect 3513 3043 3571 3049
rect 3513 3040 3525 3043
rect 3344 3012 3525 3040
rect 3513 3009 3525 3012
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 4062 3040 4068 3052
rect 3844 3012 4068 3040
rect 3844 3000 3850 3012
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3040 4859 3043
rect 4890 3040 4896 3052
rect 4847 3012 4896 3040
rect 4847 3009 4859 3012
rect 4801 3003 4859 3009
rect 4890 3000 4896 3012
rect 4948 3040 4954 3052
rect 5258 3040 5264 3052
rect 4948 3012 5264 3040
rect 4948 3000 4954 3012
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 2915 2944 3004 2972
rect 3329 2975 3387 2981
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 3329 2941 3341 2975
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 1488 2836 1494 2860
rect 1482 2808 1494 2836
rect 1546 2808 1552 2860
rect 1489 2805 1501 2808
rect 1535 2805 1547 2808
rect 1489 2799 1547 2805
rect 2958 2796 2964 2848
rect 3016 2836 3022 2848
rect 3344 2836 3372 2935
rect 4246 2932 4252 2984
rect 4304 2972 4310 2984
rect 4709 2975 4767 2981
rect 4709 2972 4721 2975
rect 4304 2944 4721 2972
rect 4304 2932 4310 2944
rect 4709 2941 4721 2944
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 3789 2907 3847 2913
rect 3789 2873 3801 2907
rect 3835 2904 3847 2907
rect 3970 2904 3976 2916
rect 3835 2876 3976 2904
rect 3835 2873 3847 2876
rect 3789 2867 3847 2873
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 4341 2907 4399 2913
rect 4341 2873 4353 2907
rect 4387 2904 4399 2907
rect 4430 2904 4436 2916
rect 4387 2876 4436 2904
rect 4387 2873 4399 2876
rect 4341 2867 4399 2873
rect 4430 2864 4436 2876
rect 4488 2864 4494 2916
rect 3016 2808 3372 2836
rect 3513 2839 3571 2845
rect 3016 2796 3022 2808
rect 3513 2805 3525 2839
rect 3559 2836 3571 2839
rect 3602 2836 3608 2848
rect 3559 2808 3608 2836
rect 3559 2805 3571 2808
rect 3513 2799 3571 2805
rect 3602 2796 3608 2808
rect 3660 2796 3666 2848
rect 3697 2839 3755 2845
rect 3697 2805 3709 2839
rect 3743 2836 3755 2839
rect 3878 2836 3884 2848
rect 3743 2808 3884 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 4157 2839 4215 2845
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 4798 2836 4804 2848
rect 4203 2808 4804 2836
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 1104 2746 5888 2768
rect 1104 2694 2750 2746
rect 2802 2694 2814 2746
rect 2866 2694 2878 2746
rect 2930 2694 2942 2746
rect 2994 2694 3006 2746
rect 3058 2694 5888 2746
rect 1104 2672 5888 2694
rect 2222 2592 2228 2644
rect 2280 2592 2286 2644
rect 2590 2592 2596 2644
rect 2648 2632 2654 2644
rect 2869 2635 2927 2641
rect 2869 2632 2881 2635
rect 2648 2604 2881 2632
rect 2648 2592 2654 2604
rect 2869 2601 2881 2604
rect 2915 2601 2927 2635
rect 2869 2595 2927 2601
rect 3326 2592 3332 2644
rect 3384 2632 3390 2644
rect 3513 2635 3571 2641
rect 3513 2632 3525 2635
rect 3384 2604 3525 2632
rect 3384 2592 3390 2604
rect 3513 2601 3525 2604
rect 3559 2601 3571 2635
rect 3513 2595 3571 2601
rect 3970 2592 3976 2644
rect 4028 2592 4034 2644
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4801 2635 4859 2641
rect 4801 2632 4813 2635
rect 4212 2604 4813 2632
rect 4212 2592 4218 2604
rect 4801 2601 4813 2604
rect 4847 2601 4859 2635
rect 4801 2595 4859 2601
rect 4982 2592 4988 2644
rect 5040 2592 5046 2644
rect 5258 2592 5264 2644
rect 5316 2592 5322 2644
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 3142 2564 3148 2576
rect 1627 2536 3148 2564
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 3142 2524 3148 2536
rect 3200 2524 3206 2576
rect 1394 2388 1400 2440
rect 1452 2388 1458 2440
rect 2038 2388 2044 2440
rect 2096 2388 2102 2440
rect 2682 2388 2688 2440
rect 2740 2388 2746 2440
rect 3326 2388 3332 2440
rect 3384 2388 3390 2440
rect 4154 2388 4160 2440
rect 4212 2388 4218 2440
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 5184 2360 5212 2391
rect 5258 2388 5264 2440
rect 5316 2428 5322 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5316 2400 5457 2428
rect 5316 2388 5322 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 5810 2360 5816 2372
rect 5184 2332 5816 2360
rect 5810 2320 5816 2332
rect 5868 2320 5874 2372
rect 1104 2202 5888 2224
rect 1104 2150 3410 2202
rect 3462 2150 3474 2202
rect 3526 2150 3538 2202
rect 3590 2150 3602 2202
rect 3654 2150 3666 2202
rect 3718 2150 5888 2202
rect 1104 2128 5888 2150
<< via1 >>
rect 3410 6502 3462 6554
rect 3474 6502 3526 6554
rect 3538 6502 3590 6554
rect 3602 6502 3654 6554
rect 3666 6502 3718 6554
rect 3240 6400 3292 6452
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 3332 6264 3384 6316
rect 3148 6196 3200 6248
rect 3884 6128 3936 6180
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 2412 6103 2464 6112
rect 2412 6069 2421 6103
rect 2421 6069 2455 6103
rect 2455 6069 2464 6103
rect 2412 6060 2464 6069
rect 3240 6060 3292 6112
rect 3792 6060 3844 6112
rect 4620 6060 4672 6112
rect 2750 5958 2802 6010
rect 2814 5958 2866 6010
rect 2878 5958 2930 6010
rect 2942 5958 2994 6010
rect 3006 5958 3058 6010
rect 1676 5856 1728 5908
rect 2228 5856 2280 5908
rect 2964 5856 3016 5908
rect 3148 5856 3200 5908
rect 3056 5788 3108 5840
rect 1860 5720 1912 5772
rect 3884 5763 3936 5772
rect 3884 5729 3893 5763
rect 3893 5729 3927 5763
rect 3927 5729 3936 5763
rect 3884 5720 3936 5729
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 2044 5652 2096 5704
rect 2136 5652 2188 5704
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 1860 5516 1912 5568
rect 2228 5516 2280 5568
rect 2320 5516 2372 5568
rect 2780 5627 2832 5636
rect 2780 5593 2789 5627
rect 2789 5593 2823 5627
rect 2823 5593 2832 5627
rect 2780 5584 2832 5593
rect 4068 5584 4120 5636
rect 2596 5516 2648 5568
rect 3148 5516 3200 5568
rect 3976 5516 4028 5568
rect 5172 5627 5224 5636
rect 5172 5593 5181 5627
rect 5181 5593 5215 5627
rect 5215 5593 5224 5627
rect 5172 5584 5224 5593
rect 4528 5516 4580 5568
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 3410 5414 3462 5466
rect 3474 5414 3526 5466
rect 3538 5414 3590 5466
rect 3602 5414 3654 5466
rect 3666 5414 3718 5466
rect 1676 5312 1728 5364
rect 2044 5312 2096 5364
rect 2320 5312 2372 5364
rect 2872 5312 2924 5364
rect 3240 5355 3292 5364
rect 3240 5321 3249 5355
rect 3249 5321 3283 5355
rect 3283 5321 3292 5355
rect 3240 5312 3292 5321
rect 2412 5244 2464 5296
rect 2964 5244 3016 5296
rect 3516 5244 3568 5296
rect 3884 5312 3936 5364
rect 4068 5312 4120 5364
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 4160 5219 4212 5228
rect 4160 5185 4169 5219
rect 4169 5185 4203 5219
rect 4203 5185 4212 5219
rect 4160 5176 4212 5185
rect 4252 5219 4304 5228
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 4252 5176 4304 5185
rect 4344 5219 4396 5228
rect 4344 5185 4358 5219
rect 4358 5185 4392 5219
rect 4392 5185 4396 5219
rect 4344 5176 4396 5185
rect 4528 5176 4580 5228
rect 4620 5219 4672 5228
rect 4620 5185 4629 5219
rect 4629 5185 4663 5219
rect 4663 5185 4672 5219
rect 4620 5176 4672 5185
rect 4804 5219 4856 5228
rect 4804 5185 4813 5219
rect 4813 5185 4847 5219
rect 4847 5185 4856 5219
rect 4804 5176 4856 5185
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 2228 5108 2280 5160
rect 2780 5108 2832 5160
rect 3056 5108 3108 5160
rect 3332 5040 3384 5092
rect 3976 5040 4028 5092
rect 5172 5040 5224 5092
rect 2320 4972 2372 5024
rect 4160 4972 4212 5024
rect 2750 4870 2802 4922
rect 2814 4870 2866 4922
rect 2878 4870 2930 4922
rect 2942 4870 2994 4922
rect 3006 4870 3058 4922
rect 1952 4768 2004 4820
rect 2136 4768 2188 4820
rect 2228 4811 2280 4820
rect 2228 4777 2237 4811
rect 2237 4777 2271 4811
rect 2271 4777 2280 4811
rect 2228 4768 2280 4777
rect 3148 4768 3200 4820
rect 1860 4700 1912 4752
rect 1768 4564 1820 4616
rect 3056 4700 3108 4752
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 2964 4607 3016 4616
rect 2964 4573 2973 4607
rect 2973 4573 3007 4607
rect 3007 4573 3016 4607
rect 2964 4564 3016 4573
rect 3056 4564 3108 4616
rect 3332 4768 3384 4820
rect 3608 4811 3660 4820
rect 3608 4777 3617 4811
rect 3617 4777 3651 4811
rect 3651 4777 3660 4811
rect 3608 4768 3660 4777
rect 4160 4768 4212 4820
rect 5448 4811 5500 4820
rect 5448 4777 5457 4811
rect 5457 4777 5491 4811
rect 5491 4777 5500 4811
rect 5448 4768 5500 4777
rect 4160 4632 4212 4684
rect 3700 4564 3752 4616
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 3976 4607 4028 4616
rect 3976 4573 3993 4607
rect 3993 4573 4028 4607
rect 3976 4564 4028 4573
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 2044 4471 2096 4480
rect 2044 4437 2053 4471
rect 2053 4437 2087 4471
rect 2087 4437 2096 4471
rect 2044 4428 2096 4437
rect 2320 4428 2372 4480
rect 4160 4539 4212 4548
rect 4160 4505 4169 4539
rect 4169 4505 4203 4539
rect 4203 4505 4212 4539
rect 4160 4496 4212 4505
rect 4804 4496 4856 4548
rect 5172 4539 5224 4548
rect 5172 4505 5181 4539
rect 5181 4505 5215 4539
rect 5215 4505 5224 4539
rect 5172 4496 5224 4505
rect 4712 4428 4764 4480
rect 4896 4471 4948 4480
rect 4896 4437 4905 4471
rect 4905 4437 4939 4471
rect 4939 4437 4948 4471
rect 4896 4428 4948 4437
rect 3410 4326 3462 4378
rect 3474 4326 3526 4378
rect 3538 4326 3590 4378
rect 3602 4326 3654 4378
rect 3666 4326 3718 4378
rect 3056 4224 3108 4276
rect 3424 4267 3476 4276
rect 3424 4233 3433 4267
rect 3433 4233 3467 4267
rect 3467 4233 3476 4267
rect 3424 4224 3476 4233
rect 3148 4156 3200 4208
rect 3792 4224 3844 4276
rect 4252 4224 4304 4276
rect 4896 4224 4948 4276
rect 5172 4267 5224 4276
rect 5172 4233 5181 4267
rect 5181 4233 5215 4267
rect 5215 4233 5224 4267
rect 5172 4224 5224 4233
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 2228 4088 2280 4140
rect 2412 3952 2464 4004
rect 3516 4088 3568 4140
rect 3608 4131 3660 4140
rect 3608 4097 3617 4131
rect 3617 4097 3651 4131
rect 3651 4097 3660 4131
rect 3608 4088 3660 4097
rect 3976 4088 4028 4140
rect 4160 4088 4212 4140
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 3516 3952 3568 4004
rect 3792 3884 3844 3936
rect 4620 3884 4672 3936
rect 4896 3884 4948 3936
rect 2750 3782 2802 3834
rect 2814 3782 2866 3834
rect 2878 3782 2930 3834
rect 2942 3782 2994 3834
rect 3006 3782 3058 3834
rect 2136 3680 2188 3732
rect 2504 3680 2556 3732
rect 3976 3680 4028 3732
rect 4252 3680 4304 3732
rect 4344 3680 4396 3732
rect 4620 3680 4672 3732
rect 4712 3723 4764 3732
rect 4712 3689 4721 3723
rect 4721 3689 4755 3723
rect 4755 3689 4764 3723
rect 4712 3680 4764 3689
rect 2964 3612 3016 3664
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 3884 3544 3936 3596
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 1768 3451 1820 3460
rect 1768 3417 1777 3451
rect 1777 3417 1811 3451
rect 1811 3417 1820 3451
rect 1768 3408 1820 3417
rect 2320 3408 2372 3460
rect 2412 3383 2464 3392
rect 2412 3349 2421 3383
rect 2421 3349 2455 3383
rect 2455 3349 2464 3383
rect 2412 3340 2464 3349
rect 2504 3340 2556 3392
rect 3240 3408 3292 3460
rect 3516 3519 3568 3528
rect 3516 3485 3525 3519
rect 3525 3485 3559 3519
rect 3559 3485 3568 3519
rect 3516 3476 3568 3485
rect 3608 3519 3660 3528
rect 3608 3485 3617 3519
rect 3617 3485 3651 3519
rect 3651 3485 3660 3519
rect 3608 3476 3660 3485
rect 3792 3476 3844 3528
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 4344 3451 4396 3460
rect 4344 3417 4353 3451
rect 4353 3417 4387 3451
rect 4387 3417 4396 3451
rect 4344 3408 4396 3417
rect 4896 3451 4948 3460
rect 4896 3417 4905 3451
rect 4905 3417 4939 3451
rect 4939 3417 4948 3451
rect 4896 3408 4948 3417
rect 4436 3340 4488 3392
rect 3410 3238 3462 3290
rect 3474 3238 3526 3290
rect 3538 3238 3590 3290
rect 3602 3238 3654 3290
rect 3666 3238 3718 3290
rect 1676 3136 1728 3188
rect 2412 3136 2464 3188
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 2228 2932 2280 2984
rect 2596 2932 2648 2984
rect 4068 3136 4120 3188
rect 4344 3136 4396 3188
rect 3148 3068 3200 3120
rect 3332 3068 3384 3120
rect 3608 3068 3660 3120
rect 4160 3111 4212 3120
rect 4160 3077 4169 3111
rect 4169 3077 4203 3111
rect 4203 3077 4212 3111
rect 4160 3068 4212 3077
rect 4988 3068 5040 3120
rect 3792 3000 3844 3052
rect 4068 3000 4120 3052
rect 4896 3000 4948 3052
rect 5264 3000 5316 3052
rect 1494 2839 1546 2860
rect 1494 2808 1501 2839
rect 1501 2808 1535 2839
rect 1535 2808 1546 2839
rect 2964 2796 3016 2848
rect 4252 2932 4304 2984
rect 3976 2864 4028 2916
rect 4436 2864 4488 2916
rect 3608 2796 3660 2848
rect 3884 2796 3936 2848
rect 4804 2796 4856 2848
rect 2750 2694 2802 2746
rect 2814 2694 2866 2746
rect 2878 2694 2930 2746
rect 2942 2694 2994 2746
rect 3006 2694 3058 2746
rect 2228 2635 2280 2644
rect 2228 2601 2237 2635
rect 2237 2601 2271 2635
rect 2271 2601 2280 2635
rect 2228 2592 2280 2601
rect 2596 2592 2648 2644
rect 3332 2592 3384 2644
rect 3976 2635 4028 2644
rect 3976 2601 3985 2635
rect 3985 2601 4019 2635
rect 4019 2601 4028 2635
rect 3976 2592 4028 2601
rect 4160 2592 4212 2644
rect 4988 2635 5040 2644
rect 4988 2601 4997 2635
rect 4997 2601 5031 2635
rect 5031 2601 5040 2635
rect 4988 2592 5040 2601
rect 5264 2635 5316 2644
rect 5264 2601 5273 2635
rect 5273 2601 5307 2635
rect 5307 2601 5316 2635
rect 5264 2592 5316 2601
rect 3148 2524 3200 2576
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5264 2388 5316 2440
rect 5816 2320 5868 2372
rect 3410 2150 3462 2202
rect 3474 2150 3526 2202
rect 3538 2150 3590 2202
rect 3602 2150 3654 2202
rect 3666 2150 3718 2202
<< metal2 >>
rect 1436 6670 1636 6790
rect 3240 6690 3296 6890
rect 1502 6118 1530 6670
rect 3252 6458 3280 6690
rect 3410 6556 3718 6565
rect 3410 6554 3416 6556
rect 3472 6554 3496 6556
rect 3552 6554 3576 6556
rect 3632 6554 3656 6556
rect 3712 6554 3718 6556
rect 3472 6502 3474 6554
rect 3654 6502 3656 6554
rect 3410 6500 3416 6502
rect 3472 6500 3496 6502
rect 3552 6500 3576 6502
rect 3632 6500 3656 6502
rect 3712 6500 3718 6502
rect 3410 6491 3718 6500
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 774 5688 974 5740
rect 1400 5704 1452 5710
rect 774 5660 1400 5688
rect 774 5620 974 5660
rect 1400 5646 1452 5652
rect 1688 5370 1716 5850
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1398 4176 1454 4185
rect 1398 4111 1400 4120
rect 1452 4111 1454 4120
rect 1400 4082 1452 4088
rect 1688 3482 1716 5306
rect 1780 4622 1808 6258
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1872 5574 1900 5714
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1872 4758 1900 5510
rect 2056 5370 2084 5646
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1964 4826 1992 5170
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1860 4752 1912 4758
rect 1860 4694 1912 4700
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1872 3602 1900 4694
rect 2056 4486 2084 5306
rect 2148 4826 2176 5646
rect 2240 5574 2268 5850
rect 2424 5710 2452 6054
rect 2750 6012 3058 6021
rect 2750 6010 2756 6012
rect 2812 6010 2836 6012
rect 2892 6010 2916 6012
rect 2972 6010 2996 6012
rect 3052 6010 3058 6012
rect 2812 5958 2814 6010
rect 2994 5958 2996 6010
rect 2750 5956 2756 5958
rect 2812 5956 2836 5958
rect 2892 5956 2916 5958
rect 2972 5956 2996 5958
rect 3052 5956 3058 5958
rect 2750 5947 3058 5956
rect 3160 5914 3188 6190
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2332 5370 2360 5510
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 2240 4826 2268 5102
rect 2332 5030 2360 5306
rect 2412 5296 2464 5302
rect 2608 5250 2636 5510
rect 2464 5244 2636 5250
rect 2412 5238 2636 5244
rect 2424 5222 2636 5238
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 2056 3534 2084 4422
rect 2148 3738 2176 4762
rect 2608 4622 2636 5222
rect 2792 5166 2820 5578
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2884 5273 2912 5306
rect 2976 5302 3004 5850
rect 3056 5840 3108 5846
rect 3056 5782 3108 5788
rect 2964 5296 3016 5302
rect 2870 5264 2926 5273
rect 2964 5238 3016 5244
rect 2870 5199 2926 5208
rect 3068 5166 3096 5782
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 2750 4924 3058 4933
rect 2750 4922 2756 4924
rect 2812 4922 2836 4924
rect 2892 4922 2916 4924
rect 2972 4922 2996 4924
rect 3052 4922 3058 4924
rect 2812 4870 2814 4922
rect 2994 4870 2996 4922
rect 2750 4868 2756 4870
rect 2812 4868 2836 4870
rect 2892 4868 2916 4870
rect 2972 4868 2996 4870
rect 3052 4868 3058 4870
rect 2750 4859 3058 4868
rect 3160 4826 3188 5510
rect 3252 5370 3280 6054
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3056 4752 3108 4758
rect 3252 4706 3280 5306
rect 3344 5273 3372 6258
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3410 5468 3718 5477
rect 3410 5466 3416 5468
rect 3472 5466 3496 5468
rect 3552 5466 3576 5468
rect 3632 5466 3656 5468
rect 3712 5466 3718 5468
rect 3472 5414 3474 5466
rect 3654 5414 3656 5466
rect 3410 5412 3416 5414
rect 3472 5412 3496 5414
rect 3552 5412 3576 5414
rect 3632 5412 3656 5414
rect 3712 5412 3718 5414
rect 3410 5403 3718 5412
rect 3804 5352 3832 6054
rect 3896 5778 3924 6122
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3896 5370 3924 5714
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3620 5324 3832 5352
rect 3884 5364 3936 5370
rect 3516 5296 3568 5302
rect 3330 5264 3386 5273
rect 3386 5222 3464 5250
rect 3516 5238 3568 5244
rect 3330 5199 3386 5208
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3344 4826 3372 5034
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3108 4700 3280 4706
rect 3056 4694 3280 4700
rect 3068 4678 3280 4694
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 3056 4616 3108 4622
rect 3108 4576 3280 4604
rect 3056 4558 3108 4564
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 2044 3528 2096 3534
rect 1688 3466 1808 3482
rect 2044 3470 2096 3476
rect 1688 3460 1820 3466
rect 1688 3454 1768 3460
rect 1688 3194 1716 3454
rect 1768 3402 1820 3408
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 2240 2990 2268 4082
rect 2332 3466 2360 4422
rect 2976 4026 3004 4558
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 3068 4049 3096 4218
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 2412 4004 2464 4010
rect 2412 3946 2464 3952
rect 2516 3998 3004 4026
rect 3054 4040 3110 4049
rect 2424 3482 2452 3946
rect 2516 3738 2544 3998
rect 3054 3975 3110 3984
rect 2750 3836 3058 3845
rect 2750 3834 2756 3836
rect 2812 3834 2836 3836
rect 2892 3834 2916 3836
rect 2972 3834 2996 3836
rect 3052 3834 3058 3836
rect 2812 3782 2814 3834
rect 2994 3782 2996 3834
rect 2750 3780 2756 3782
rect 2812 3780 2836 3782
rect 2892 3780 2916 3782
rect 2972 3780 2996 3782
rect 3052 3780 3058 3782
rect 2750 3771 3058 3780
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 2320 3460 2372 3466
rect 2424 3454 2544 3482
rect 2320 3402 2372 3408
rect 2516 3398 2544 3454
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2424 3194 2452 3334
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2516 3058 2544 3334
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 1494 2860 1546 2866
rect 1483 2804 1492 2860
rect 1548 2804 1557 2860
rect 1494 2802 1546 2804
rect 2516 2774 2544 2994
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2240 2746 2544 2774
rect 2240 2650 2268 2746
rect 2608 2650 2636 2926
rect 2976 2854 3004 3606
rect 3160 3126 3188 4150
rect 3252 3466 3280 4576
rect 3436 4468 3464 5222
rect 3528 4593 3556 5238
rect 3620 4826 3648 5324
rect 3884 5306 3936 5312
rect 3896 4978 3924 5306
rect 3988 5098 4016 5510
rect 4080 5370 4108 5578
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4080 5250 4108 5306
rect 4080 5234 4200 5250
rect 4540 5234 4568 5510
rect 4632 5234 4660 6054
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 4894 5264 4950 5273
rect 4080 5228 4212 5234
rect 4080 5222 4160 5228
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3712 4950 3924 4978
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3712 4622 3740 4950
rect 3988 4842 4016 5034
rect 3804 4814 4016 4842
rect 3804 4622 3832 4814
rect 3700 4616 3752 4622
rect 3514 4584 3570 4593
rect 3700 4558 3752 4564
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3976 4616 4028 4622
rect 4080 4604 4108 5222
rect 4160 5170 4212 5176
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4804 5228 4856 5234
rect 4894 5199 4896 5208
rect 4804 5170 4856 5176
rect 4948 5199 4950 5208
rect 4896 5170 4948 5176
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4172 4826 4200 4966
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4264 4706 4292 5170
rect 4172 4690 4292 4706
rect 4160 4684 4292 4690
rect 4212 4678 4292 4684
rect 4160 4626 4212 4632
rect 4028 4576 4108 4604
rect 4252 4616 4304 4622
rect 4158 4584 4214 4593
rect 3976 4558 4028 4564
rect 3514 4519 3570 4528
rect 3344 4440 3464 4468
rect 3344 4264 3372 4440
rect 3410 4380 3718 4389
rect 3410 4378 3416 4380
rect 3472 4378 3496 4380
rect 3552 4378 3576 4380
rect 3632 4378 3656 4380
rect 3712 4378 3718 4380
rect 3472 4326 3474 4378
rect 3654 4326 3656 4378
rect 3410 4324 3416 4326
rect 3472 4324 3496 4326
rect 3552 4324 3576 4326
rect 3632 4324 3656 4326
rect 3712 4324 3718 4326
rect 3410 4315 3718 4324
rect 3804 4282 3832 4558
rect 4252 4558 4304 4564
rect 4158 4519 4160 4528
rect 4212 4519 4214 4528
rect 4160 4490 4212 4496
rect 4172 4298 4200 4490
rect 3424 4276 3476 4282
rect 3344 4236 3424 4264
rect 3424 4218 3476 4224
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 4080 4270 4200 4298
rect 4264 4282 4292 4558
rect 4252 4276 4304 4282
rect 4080 4185 4108 4270
rect 4252 4218 4304 4224
rect 3514 4176 3570 4185
rect 4066 4176 4122 4185
rect 3514 4111 3516 4120
rect 3568 4111 3570 4120
rect 3608 4140 3660 4146
rect 3516 4082 3568 4088
rect 3608 4082 3660 4088
rect 3976 4140 4028 4146
rect 4066 4111 4122 4120
rect 4160 4140 4212 4146
rect 3976 4082 4028 4088
rect 4160 4082 4212 4088
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 3330 4040 3386 4049
rect 3330 3975 3386 3984
rect 3516 4004 3568 4010
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 3344 3126 3372 3975
rect 3516 3946 3568 3952
rect 3528 3534 3556 3946
rect 3620 3534 3648 4082
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3534 3832 3878
rect 3988 3738 4016 4082
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3620 3380 3648 3470
rect 3620 3352 3832 3380
rect 3410 3292 3718 3301
rect 3410 3290 3416 3292
rect 3472 3290 3496 3292
rect 3552 3290 3576 3292
rect 3632 3290 3656 3292
rect 3712 3290 3718 3292
rect 3472 3238 3474 3290
rect 3654 3238 3656 3290
rect 3410 3236 3416 3238
rect 3472 3236 3496 3238
rect 3552 3236 3576 3238
rect 3632 3236 3656 3238
rect 3712 3236 3718 3238
rect 3410 3227 3718 3236
rect 3148 3120 3200 3126
rect 3148 3062 3200 3068
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 3608 3120 3660 3126
rect 3608 3062 3660 3068
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2750 2748 3058 2757
rect 2750 2746 2756 2748
rect 2812 2746 2836 2748
rect 2892 2746 2916 2748
rect 2972 2746 2996 2748
rect 3052 2746 3058 2748
rect 2812 2694 2814 2746
rect 2994 2694 2996 2746
rect 2750 2692 2756 2694
rect 2812 2692 2836 2694
rect 2892 2692 2916 2694
rect 2972 2692 2996 2694
rect 3052 2692 3058 2694
rect 2750 2683 3058 2692
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 3160 2582 3188 3062
rect 3344 2650 3372 3062
rect 3620 2854 3648 3062
rect 3804 3058 3832 3352
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3896 2854 3924 3538
rect 3988 2922 4016 3674
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4080 3194 4108 3470
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4172 3126 4200 4082
rect 4264 3738 4292 4082
rect 4356 3738 4384 5170
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4632 3942 4660 4558
rect 4816 4554 4844 5170
rect 5184 5098 5212 5578
rect 5448 5568 5500 5574
rect 5446 5536 5448 5545
rect 5500 5536 5502 5545
rect 5446 5471 5502 5480
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5446 4856 5502 4865
rect 5446 4791 5448 4800
rect 5500 4791 5502 4800
rect 5448 4762 5500 4768
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4632 3738 4660 3878
rect 4724 3738 4752 4422
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4356 3194 4384 3402
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3988 2650 4016 2858
rect 4080 2774 4108 2994
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 4264 2774 4292 2926
rect 4448 2922 4476 3334
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4816 2854 4844 4490
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4908 4282 4936 4422
rect 5184 4282 5212 4490
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3466 4936 3878
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4908 3058 4936 3402
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4080 2746 4292 2774
rect 4172 2650 4200 2746
rect 5000 2650 5028 3062
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5276 2650 5304 2994
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 5184 2502 5304 2530
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 1412 1972 1440 2382
rect 2056 1998 2084 2382
rect 2700 2004 2728 2382
rect 1400 1772 1456 1972
rect 2040 1798 2096 1998
rect 2684 1804 2740 2004
rect 3344 2002 3372 2382
rect 3410 2204 3718 2213
rect 3410 2202 3416 2204
rect 3472 2202 3496 2204
rect 3552 2202 3576 2204
rect 3632 2202 3656 2204
rect 3712 2202 3718 2204
rect 3472 2150 3474 2202
rect 3654 2150 3656 2202
rect 3410 2148 3416 2150
rect 3472 2148 3496 2150
rect 3552 2148 3576 2150
rect 3632 2148 3656 2150
rect 3712 2148 3718 2150
rect 3410 2139 3718 2148
rect 4172 2010 4200 2382
rect 4632 2014 4660 2382
rect 3324 1802 3380 2002
rect 4158 1810 4214 2010
rect 4616 1814 4672 2014
rect 5184 2006 5212 2502
rect 5276 2446 5304 2502
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5828 2018 5856 2314
rect 5166 1806 5222 2006
rect 5808 1818 5864 2018
<< via2 >>
rect 3416 6554 3472 6556
rect 3496 6554 3552 6556
rect 3576 6554 3632 6556
rect 3656 6554 3712 6556
rect 3416 6502 3462 6554
rect 3462 6502 3472 6554
rect 3496 6502 3526 6554
rect 3526 6502 3538 6554
rect 3538 6502 3552 6554
rect 3576 6502 3590 6554
rect 3590 6502 3602 6554
rect 3602 6502 3632 6554
rect 3656 6502 3666 6554
rect 3666 6502 3712 6554
rect 3416 6500 3472 6502
rect 3496 6500 3552 6502
rect 3576 6500 3632 6502
rect 3656 6500 3712 6502
rect 1398 4140 1454 4176
rect 1398 4120 1400 4140
rect 1400 4120 1452 4140
rect 1452 4120 1454 4140
rect 2756 6010 2812 6012
rect 2836 6010 2892 6012
rect 2916 6010 2972 6012
rect 2996 6010 3052 6012
rect 2756 5958 2802 6010
rect 2802 5958 2812 6010
rect 2836 5958 2866 6010
rect 2866 5958 2878 6010
rect 2878 5958 2892 6010
rect 2916 5958 2930 6010
rect 2930 5958 2942 6010
rect 2942 5958 2972 6010
rect 2996 5958 3006 6010
rect 3006 5958 3052 6010
rect 2756 5956 2812 5958
rect 2836 5956 2892 5958
rect 2916 5956 2972 5958
rect 2996 5956 3052 5958
rect 2870 5208 2926 5264
rect 2756 4922 2812 4924
rect 2836 4922 2892 4924
rect 2916 4922 2972 4924
rect 2996 4922 3052 4924
rect 2756 4870 2802 4922
rect 2802 4870 2812 4922
rect 2836 4870 2866 4922
rect 2866 4870 2878 4922
rect 2878 4870 2892 4922
rect 2916 4870 2930 4922
rect 2930 4870 2942 4922
rect 2942 4870 2972 4922
rect 2996 4870 3006 4922
rect 3006 4870 3052 4922
rect 2756 4868 2812 4870
rect 2836 4868 2892 4870
rect 2916 4868 2972 4870
rect 2996 4868 3052 4870
rect 3416 5466 3472 5468
rect 3496 5466 3552 5468
rect 3576 5466 3632 5468
rect 3656 5466 3712 5468
rect 3416 5414 3462 5466
rect 3462 5414 3472 5466
rect 3496 5414 3526 5466
rect 3526 5414 3538 5466
rect 3538 5414 3552 5466
rect 3576 5414 3590 5466
rect 3590 5414 3602 5466
rect 3602 5414 3632 5466
rect 3656 5414 3666 5466
rect 3666 5414 3712 5466
rect 3416 5412 3472 5414
rect 3496 5412 3552 5414
rect 3576 5412 3632 5414
rect 3656 5412 3712 5414
rect 3330 5208 3386 5264
rect 3054 3984 3110 4040
rect 2756 3834 2812 3836
rect 2836 3834 2892 3836
rect 2916 3834 2972 3836
rect 2996 3834 3052 3836
rect 2756 3782 2802 3834
rect 2802 3782 2812 3834
rect 2836 3782 2866 3834
rect 2866 3782 2878 3834
rect 2878 3782 2892 3834
rect 2916 3782 2930 3834
rect 2930 3782 2942 3834
rect 2942 3782 2972 3834
rect 2996 3782 3006 3834
rect 3006 3782 3052 3834
rect 2756 3780 2812 3782
rect 2836 3780 2892 3782
rect 2916 3780 2972 3782
rect 2996 3780 3052 3782
rect 1492 2808 1494 2860
rect 1494 2808 1546 2860
rect 1546 2808 1548 2860
rect 1492 2804 1548 2808
rect 3514 4528 3570 4584
rect 4894 5228 4950 5264
rect 4894 5208 4896 5228
rect 4896 5208 4948 5228
rect 4948 5208 4950 5228
rect 3416 4378 3472 4380
rect 3496 4378 3552 4380
rect 3576 4378 3632 4380
rect 3656 4378 3712 4380
rect 3416 4326 3462 4378
rect 3462 4326 3472 4378
rect 3496 4326 3526 4378
rect 3526 4326 3538 4378
rect 3538 4326 3552 4378
rect 3576 4326 3590 4378
rect 3590 4326 3602 4378
rect 3602 4326 3632 4378
rect 3656 4326 3666 4378
rect 3666 4326 3712 4378
rect 3416 4324 3472 4326
rect 3496 4324 3552 4326
rect 3576 4324 3632 4326
rect 3656 4324 3712 4326
rect 4158 4548 4214 4584
rect 4158 4528 4160 4548
rect 4160 4528 4212 4548
rect 4212 4528 4214 4548
rect 3514 4140 3570 4176
rect 3514 4120 3516 4140
rect 3516 4120 3568 4140
rect 3568 4120 3570 4140
rect 4066 4120 4122 4176
rect 3330 3984 3386 4040
rect 3416 3290 3472 3292
rect 3496 3290 3552 3292
rect 3576 3290 3632 3292
rect 3656 3290 3712 3292
rect 3416 3238 3462 3290
rect 3462 3238 3472 3290
rect 3496 3238 3526 3290
rect 3526 3238 3538 3290
rect 3538 3238 3552 3290
rect 3576 3238 3590 3290
rect 3590 3238 3602 3290
rect 3602 3238 3632 3290
rect 3656 3238 3666 3290
rect 3666 3238 3712 3290
rect 3416 3236 3472 3238
rect 3496 3236 3552 3238
rect 3576 3236 3632 3238
rect 3656 3236 3712 3238
rect 2756 2746 2812 2748
rect 2836 2746 2892 2748
rect 2916 2746 2972 2748
rect 2996 2746 3052 2748
rect 2756 2694 2802 2746
rect 2802 2694 2812 2746
rect 2836 2694 2866 2746
rect 2866 2694 2878 2746
rect 2878 2694 2892 2746
rect 2916 2694 2930 2746
rect 2930 2694 2942 2746
rect 2942 2694 2972 2746
rect 2996 2694 3006 2746
rect 3006 2694 3052 2746
rect 2756 2692 2812 2694
rect 2836 2692 2892 2694
rect 2916 2692 2972 2694
rect 2996 2692 3052 2694
rect 5446 5516 5448 5536
rect 5448 5516 5500 5536
rect 5500 5516 5502 5536
rect 5446 5480 5502 5516
rect 5446 4820 5502 4856
rect 5446 4800 5448 4820
rect 5448 4800 5500 4820
rect 5500 4800 5502 4820
rect 3416 2202 3472 2204
rect 3496 2202 3552 2204
rect 3576 2202 3632 2204
rect 3656 2202 3712 2204
rect 3416 2150 3462 2202
rect 3462 2150 3472 2202
rect 3496 2150 3526 2202
rect 3526 2150 3538 2202
rect 3538 2150 3552 2202
rect 3576 2150 3590 2202
rect 3590 2150 3602 2202
rect 3602 2150 3632 2202
rect 3656 2150 3666 2202
rect 3666 2150 3712 2202
rect 3416 2148 3472 2150
rect 3496 2148 3552 2150
rect 3576 2148 3632 2150
rect 3656 2148 3712 2150
<< metal3 >>
rect 3406 6560 3722 6561
rect 3406 6496 3412 6560
rect 3476 6496 3492 6560
rect 3556 6496 3572 6560
rect 3636 6496 3652 6560
rect 3716 6496 3722 6560
rect 3406 6495 3722 6496
rect 2746 6016 3062 6017
rect 2746 5952 2752 6016
rect 2816 5952 2832 6016
rect 2896 5952 2912 6016
rect 2976 5952 2992 6016
rect 3056 5952 3062 6016
rect 2746 5951 3062 5952
rect 5441 5538 5507 5541
rect 6258 5538 7058 5568
rect 5441 5536 7058 5538
rect 5441 5480 5446 5536
rect 5502 5480 7058 5536
rect 5441 5478 7058 5480
rect 5441 5475 5507 5478
rect 3406 5472 3722 5473
rect 3406 5408 3412 5472
rect 3476 5408 3492 5472
rect 3556 5408 3572 5472
rect 3636 5408 3652 5472
rect 3716 5408 3722 5472
rect 6258 5448 7058 5478
rect 3406 5407 3722 5408
rect 2865 5266 2931 5269
rect 3325 5266 3391 5269
rect 4889 5266 4955 5269
rect 2865 5264 4955 5266
rect 2865 5208 2870 5264
rect 2926 5208 3330 5264
rect 3386 5208 4894 5264
rect 4950 5208 4955 5264
rect 2865 5206 4955 5208
rect 2865 5203 2931 5206
rect 3325 5203 3391 5206
rect 4889 5203 4955 5206
rect 2746 4928 3062 4929
rect 2746 4864 2752 4928
rect 2816 4864 2832 4928
rect 2896 4864 2912 4928
rect 2976 4864 2992 4928
rect 3056 4864 3062 4928
rect 2746 4863 3062 4864
rect 5441 4858 5507 4861
rect 6258 4858 7058 4888
rect 5441 4856 7058 4858
rect 5441 4800 5446 4856
rect 5502 4800 7058 4856
rect 5441 4798 7058 4800
rect 5441 4795 5507 4798
rect 6258 4768 7058 4798
rect 3509 4586 3575 4589
rect 4153 4586 4219 4589
rect 3509 4584 4219 4586
rect 3509 4528 3514 4584
rect 3570 4528 4158 4584
rect 4214 4528 4219 4584
rect 3509 4526 4219 4528
rect 3509 4523 3575 4526
rect 4153 4523 4219 4526
rect 3406 4384 3722 4385
rect 3406 4320 3412 4384
rect 3476 4320 3492 4384
rect 3556 4320 3572 4384
rect 3636 4320 3652 4384
rect 3716 4320 3722 4384
rect 3406 4319 3722 4320
rect 810 4178 1010 4196
rect 1393 4178 1459 4181
rect 810 4176 1459 4178
rect 810 4120 1398 4176
rect 1454 4120 1459 4176
rect 810 4118 1459 4120
rect 810 4096 1010 4118
rect 1393 4115 1459 4118
rect 3509 4178 3575 4181
rect 4061 4178 4127 4181
rect 3509 4176 4127 4178
rect 3509 4120 3514 4176
rect 3570 4120 4066 4176
rect 4122 4120 4127 4176
rect 3509 4118 4127 4120
rect 3509 4115 3575 4118
rect 4061 4115 4127 4118
rect 3049 4042 3115 4045
rect 3325 4042 3391 4045
rect 3049 4040 3391 4042
rect 3049 3984 3054 4040
rect 3110 3984 3330 4040
rect 3386 3984 3391 4040
rect 3049 3982 3391 3984
rect 3049 3979 3115 3982
rect 3325 3979 3391 3982
rect 2746 3840 3062 3841
rect 2746 3776 2752 3840
rect 2816 3776 2832 3840
rect 2896 3776 2912 3840
rect 2976 3776 2992 3840
rect 3056 3776 3062 3840
rect 2746 3775 3062 3776
rect 3406 3296 3722 3297
rect 3406 3232 3412 3296
rect 3476 3232 3492 3296
rect 3556 3232 3572 3296
rect 3636 3232 3652 3296
rect 3716 3232 3722 3296
rect 3406 3231 3722 3232
rect 6056 2924 6856 2962
rect 1490 2865 6856 2924
rect 1487 2864 6856 2865
rect 1487 2860 1553 2864
rect 1487 2804 1492 2860
rect 1548 2804 1553 2860
rect 6056 2842 6856 2864
rect 1487 2799 1553 2804
rect 1490 2798 1550 2799
rect 2746 2752 3062 2753
rect 2746 2688 2752 2752
rect 2816 2688 2832 2752
rect 2896 2688 2912 2752
rect 2976 2688 2992 2752
rect 3056 2688 3062 2752
rect 2746 2687 3062 2688
rect 3406 2208 3722 2209
rect 3406 2144 3412 2208
rect 3476 2144 3492 2208
rect 3556 2144 3572 2208
rect 3636 2144 3652 2208
rect 3716 2144 3722 2208
rect 3406 2143 3722 2144
<< via3 >>
rect 3412 6556 3476 6560
rect 3412 6500 3416 6556
rect 3416 6500 3472 6556
rect 3472 6500 3476 6556
rect 3412 6496 3476 6500
rect 3492 6556 3556 6560
rect 3492 6500 3496 6556
rect 3496 6500 3552 6556
rect 3552 6500 3556 6556
rect 3492 6496 3556 6500
rect 3572 6556 3636 6560
rect 3572 6500 3576 6556
rect 3576 6500 3632 6556
rect 3632 6500 3636 6556
rect 3572 6496 3636 6500
rect 3652 6556 3716 6560
rect 3652 6500 3656 6556
rect 3656 6500 3712 6556
rect 3712 6500 3716 6556
rect 3652 6496 3716 6500
rect 2752 6012 2816 6016
rect 2752 5956 2756 6012
rect 2756 5956 2812 6012
rect 2812 5956 2816 6012
rect 2752 5952 2816 5956
rect 2832 6012 2896 6016
rect 2832 5956 2836 6012
rect 2836 5956 2892 6012
rect 2892 5956 2896 6012
rect 2832 5952 2896 5956
rect 2912 6012 2976 6016
rect 2912 5956 2916 6012
rect 2916 5956 2972 6012
rect 2972 5956 2976 6012
rect 2912 5952 2976 5956
rect 2992 6012 3056 6016
rect 2992 5956 2996 6012
rect 2996 5956 3052 6012
rect 3052 5956 3056 6012
rect 2992 5952 3056 5956
rect 3412 5468 3476 5472
rect 3412 5412 3416 5468
rect 3416 5412 3472 5468
rect 3472 5412 3476 5468
rect 3412 5408 3476 5412
rect 3492 5468 3556 5472
rect 3492 5412 3496 5468
rect 3496 5412 3552 5468
rect 3552 5412 3556 5468
rect 3492 5408 3556 5412
rect 3572 5468 3636 5472
rect 3572 5412 3576 5468
rect 3576 5412 3632 5468
rect 3632 5412 3636 5468
rect 3572 5408 3636 5412
rect 3652 5468 3716 5472
rect 3652 5412 3656 5468
rect 3656 5412 3712 5468
rect 3712 5412 3716 5468
rect 3652 5408 3716 5412
rect 2752 4924 2816 4928
rect 2752 4868 2756 4924
rect 2756 4868 2812 4924
rect 2812 4868 2816 4924
rect 2752 4864 2816 4868
rect 2832 4924 2896 4928
rect 2832 4868 2836 4924
rect 2836 4868 2892 4924
rect 2892 4868 2896 4924
rect 2832 4864 2896 4868
rect 2912 4924 2976 4928
rect 2912 4868 2916 4924
rect 2916 4868 2972 4924
rect 2972 4868 2976 4924
rect 2912 4864 2976 4868
rect 2992 4924 3056 4928
rect 2992 4868 2996 4924
rect 2996 4868 3052 4924
rect 3052 4868 3056 4924
rect 2992 4864 3056 4868
rect 3412 4380 3476 4384
rect 3412 4324 3416 4380
rect 3416 4324 3472 4380
rect 3472 4324 3476 4380
rect 3412 4320 3476 4324
rect 3492 4380 3556 4384
rect 3492 4324 3496 4380
rect 3496 4324 3552 4380
rect 3552 4324 3556 4380
rect 3492 4320 3556 4324
rect 3572 4380 3636 4384
rect 3572 4324 3576 4380
rect 3576 4324 3632 4380
rect 3632 4324 3636 4380
rect 3572 4320 3636 4324
rect 3652 4380 3716 4384
rect 3652 4324 3656 4380
rect 3656 4324 3712 4380
rect 3712 4324 3716 4380
rect 3652 4320 3716 4324
rect 2752 3836 2816 3840
rect 2752 3780 2756 3836
rect 2756 3780 2812 3836
rect 2812 3780 2816 3836
rect 2752 3776 2816 3780
rect 2832 3836 2896 3840
rect 2832 3780 2836 3836
rect 2836 3780 2892 3836
rect 2892 3780 2896 3836
rect 2832 3776 2896 3780
rect 2912 3836 2976 3840
rect 2912 3780 2916 3836
rect 2916 3780 2972 3836
rect 2972 3780 2976 3836
rect 2912 3776 2976 3780
rect 2992 3836 3056 3840
rect 2992 3780 2996 3836
rect 2996 3780 3052 3836
rect 3052 3780 3056 3836
rect 2992 3776 3056 3780
rect 3412 3292 3476 3296
rect 3412 3236 3416 3292
rect 3416 3236 3472 3292
rect 3472 3236 3476 3292
rect 3412 3232 3476 3236
rect 3492 3292 3556 3296
rect 3492 3236 3496 3292
rect 3496 3236 3552 3292
rect 3552 3236 3556 3292
rect 3492 3232 3556 3236
rect 3572 3292 3636 3296
rect 3572 3236 3576 3292
rect 3576 3236 3632 3292
rect 3632 3236 3636 3292
rect 3572 3232 3636 3236
rect 3652 3292 3716 3296
rect 3652 3236 3656 3292
rect 3656 3236 3712 3292
rect 3712 3236 3716 3292
rect 3652 3232 3716 3236
rect 2752 2748 2816 2752
rect 2752 2692 2756 2748
rect 2756 2692 2812 2748
rect 2812 2692 2816 2748
rect 2752 2688 2816 2692
rect 2832 2748 2896 2752
rect 2832 2692 2836 2748
rect 2836 2692 2892 2748
rect 2892 2692 2896 2748
rect 2832 2688 2896 2692
rect 2912 2748 2976 2752
rect 2912 2692 2916 2748
rect 2916 2692 2972 2748
rect 2972 2692 2976 2748
rect 2912 2688 2976 2692
rect 2992 2748 3056 2752
rect 2992 2692 2996 2748
rect 2996 2692 3052 2748
rect 3052 2692 3056 2748
rect 2992 2688 3056 2692
rect 3412 2204 3476 2208
rect 3412 2148 3416 2204
rect 3416 2148 3472 2204
rect 3472 2148 3476 2204
rect 3412 2144 3476 2148
rect 3492 2204 3556 2208
rect 3492 2148 3496 2204
rect 3496 2148 3552 2204
rect 3552 2148 3556 2204
rect 3492 2144 3556 2148
rect 3572 2204 3636 2208
rect 3572 2148 3576 2204
rect 3576 2148 3632 2204
rect 3632 2148 3636 2204
rect 3572 2144 3636 2148
rect 3652 2204 3716 2208
rect 3652 2148 3656 2204
rect 3656 2148 3712 2204
rect 3712 2148 3716 2204
rect 3652 2144 3716 2148
<< metal4 >>
rect 2744 6016 3064 6576
rect 2744 5952 2752 6016
rect 2816 5952 2832 6016
rect 2896 5952 2912 6016
rect 2976 5952 2992 6016
rect 3056 5952 3064 6016
rect 2744 4928 3064 5952
rect 2744 4864 2752 4928
rect 2816 4864 2832 4928
rect 2896 4864 2912 4928
rect 2976 4864 2992 4928
rect 3056 4864 3064 4928
rect 2744 3840 3064 4864
rect 2744 3776 2752 3840
rect 2816 3776 2832 3840
rect 2896 3776 2912 3840
rect 2976 3776 2992 3840
rect 3056 3776 3064 3840
rect 2744 2752 3064 3776
rect 2744 2688 2752 2752
rect 2816 2688 2832 2752
rect 2896 2688 2912 2752
rect 2976 2688 2992 2752
rect 3056 2688 3064 2752
rect 2744 2128 3064 2688
rect 3404 6560 3724 6576
rect 3404 6496 3412 6560
rect 3476 6496 3492 6560
rect 3556 6496 3572 6560
rect 3636 6496 3652 6560
rect 3716 6496 3724 6560
rect 3404 5472 3724 6496
rect 3404 5408 3412 5472
rect 3476 5408 3492 5472
rect 3556 5408 3572 5472
rect 3636 5408 3652 5472
rect 3716 5408 3724 5472
rect 3404 4384 3724 5408
rect 3404 4320 3412 4384
rect 3476 4320 3492 4384
rect 3556 4320 3572 4384
rect 3636 4320 3652 4384
rect 3716 4320 3724 4384
rect 3404 3296 3724 4320
rect 3404 3232 3412 3296
rect 3476 3232 3492 3296
rect 3556 3232 3572 3296
rect 3636 3232 3652 3296
rect 3716 3232 3724 3296
rect 3404 2208 3724 3232
rect 3404 2144 3412 2208
rect 3476 2144 3492 2208
rect 3556 2144 3572 2208
rect 3636 2144 3652 2208
rect 3716 2144 3724 2208
rect 3404 2128 3724 2144
use sky130_fd_sc_hd__or3_1  _26_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform -1 0 3680 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _27_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 1748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _28_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _29_
timestamp 1696625445
transform -1 0 3680 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _30_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _31_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 2300 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 2668 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3772 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _34_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform -1 0 5060 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _35_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _36_
timestamp 1696625445
transform -1 0 4048 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _37_
timestamp 1696625445
transform 1 0 1748 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _38_
timestamp 1696625445
transform 1 0 4600 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _39_
timestamp 1696625445
transform 1 0 3772 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _40_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform -1 0 2852 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _41_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform -1 0 3496 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _42_
timestamp 1696625445
transform 1 0 1656 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _43_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform -1 0 2944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _44_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform -1 0 2208 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _45_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3864 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _46_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform -1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _47_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 2852 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _48_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform -1 0 4968 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _49_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 2392 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _50_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform -1 0 3864 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _51_
timestamp 1696625445
transform 1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _52_
timestamp 1696625445
transform -1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _53_
timestamp 1696625445
transform 1 0 4508 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _54_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform -1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _55_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 2300 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_13
timestamp 1696625445
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_20
timestamp 1696625445
transform 1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_34
timestamp 1696625445
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_41
timestamp 1696625445
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_48
timestamp 1696625445
transform 1 0 5520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_12
timestamp 1696625445
transform 1 0 2208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_20
timestamp 1696625445
transform 1 0 2944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_43 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 5060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1696625445
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_13
timestamp 1696625445
transform 1 0 2300 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_22
timestamp 1696625445
transform 1 0 3128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_42
timestamp 1696625445
transform 1 0 4968 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_48
timestamp 1696625445
transform 1 0 5520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_13
timestamp 1696625445
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_24
timestamp 1696625445
transform 1 0 3312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_32
timestamp 1696625445
transform 1 0 4048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_37
timestamp 1696625445
transform 1 0 4508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_41
timestamp 1696625445
transform 1 0 4876 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_45
timestamp 1696625445
transform 1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_42
timestamp 1696625445
transform 1 0 4968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_3
timestamp 1696625445
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_45
timestamp 1696625445
transform 1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_6
timestamp 1696625445
transform 1 0 1656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_36
timestamp 1696625445
transform 1 0 4416 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_42
timestamp 1696625445
transform 1 0 4968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_15
timestamp 1696625445
transform 1 0 2484 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_26
timestamp 1696625445
transform 1 0 3496 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_44
timestamp 1696625445
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_48
timestamp 1696625445
transform 1 0 5520 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1696625445
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1696625445
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1696625445
transform -1 0 4048 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 1380 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1696625445
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1696625445
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1696625445
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1696625445
transform -1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1696625445
transform -1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1696625445
transform -1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1696625445
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1696625445
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1696625445
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1696625445
transform 1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 5060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1696625445
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1696625445
transform 1 0 5060 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1696625445
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_8
timestamp 1696625445
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1696625445
transform -1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_9
timestamp 1696625445
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1696625445
transform -1 0 5888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_10
timestamp 1696625445
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1696625445
transform -1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_11
timestamp 1696625445
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1696625445
transform -1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_12
timestamp 1696625445
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1696625445
transform -1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_13
timestamp 1696625445
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1696625445
transform -1 0 5888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_14
timestamp 1696625445
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1696625445
transform -1 0 5888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_15
timestamp 1696625445
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1696625445
transform -1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_17
timestamp 1696625445
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_18
timestamp 1696625445
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_19
timestamp 1696625445
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_20
timestamp 1696625445
transform 1 0 3680 0 -1 6528
box -38 -48 130 592
<< labels >>
flabel metal4 s 3404 2128 3724 6576 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2744 2128 3064 6576 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 6258 5448 7058 5568 0 FreeSans 250 0 0 0 b[0]
port 2 nsew signal tristate
flabel metal3 s 6258 4768 7058 4888 0 FreeSans 250 0 0 0 b[2]
port 4 nsew signal tristate
rlabel via1 3496 6528 3496 6528 0 VGND
rlabel metal1 3496 5984 3496 5984 0 VPWR
rlabel metal1 2852 5134 2852 5134 0 _00_
rlabel metal1 2392 3706 2392 3706 0 _01_
rlabel metal2 2346 3944 2346 3944 0 _02_
rlabel metal1 3772 3638 3772 3638 0 _03_
rlabel metal1 1978 3536 1978 3536 0 _04_
rlabel metal1 2944 2958 2944 2958 0 _05_
rlabel metal1 4508 4522 4508 4522 0 _06_
rlabel metal1 4462 3434 4462 3434 0 _07_
rlabel metal1 4416 3162 4416 3162 0 _08_
rlabel metal1 4002 3366 4002 3366 0 _09_
rlabel metal1 2714 5338 2714 5338 0 _10_
rlabel metal1 4094 5134 4094 5134 0 _11_
rlabel via1 4186 5219 4186 5219 0 _12_
rlabel metal1 4076 5202 4076 5202 0 _13_
rlabel metal1 2668 5542 2668 5542 0 _14_
rlabel metal1 1978 4760 1978 4760 0 _15_
rlabel metal2 2254 4964 2254 4964 0 _16_
rlabel metal1 2300 5338 2300 5338 0 _17_
rlabel metal1 3036 5202 3036 5202 0 _18_
rlabel metal1 2392 3502 2392 3502 0 _19_
rlabel metal1 2806 4624 2806 4624 0 _20_
rlabel metal1 4600 3706 4600 3706 0 _21_
rlabel metal1 3588 4998 3588 4998 0 _22_
rlabel metal1 4324 4250 4324 4250 0 _23_
rlabel metal1 4508 4590 4508 4590 0 _24_
rlabel metal1 4968 4114 4968 4114 0 _25_
rlabel via2 5474 5525 5474 5525 0 b[0]
rlabel via2 5474 4811 5474 4811 0 b[2]
rlabel metal1 2392 2550 2392 2550 0 net1
rlabel metal1 4600 3094 4600 3094 0 net10
rlabel metal1 5060 3026 5060 3026 0 net11
rlabel metal1 4508 2618 4508 2618 0 net12
rlabel metal1 3910 2890 3910 2890 0 net13
rlabel metal2 2070 3978 2070 3978 0 net14
rlabel metal1 2116 4794 2116 4794 0 net15
rlabel metal1 4876 4998 4876 4998 0 net16
rlabel metal1 2116 3094 2116 3094 0 net17
rlabel metal2 5198 4386 5198 4386 0 net18
rlabel metal1 2070 4590 2070 4590 0 net19
rlabel metal1 2208 5542 2208 5542 0 net2
rlabel metal1 1978 5542 1978 5542 0 net3
rlabel metal2 4646 5644 4646 5644 0 net4
rlabel metal2 3818 4420 3818 4420 0 net5
rlabel metal2 3910 5950 3910 5950 0 net6
rlabel metal2 2254 2689 2254 2689 0 net7
rlabel metal1 2346 2958 2346 2958 0 net8
rlabel metal1 3450 3026 3450 3026 0 net9
rlabel metal1 866 3468 866 3468 0 p[10]
rlabel metal1 3818 6324 3818 6324 0 p[12]
rlabel metal3 1050 4148 1050 4148 0 p[13]
flabel metal2 s 3240 6690 3296 6890 0 FreeSans 250 90 0 0 p[12]
port 9 nsew signal input
flabel metal1 s 864 6338 1064 6458 0 FreeSans 250 0 0 0 p[14]
port 11 nsew signal input
flabel metal1 s 798 6164 998 6284 0 FreeSans 250 0 0 0 p[9]
port 20 nsew signal input
flabel metal1 s 844 4548 1044 4668 0 FreeSans 250 0 0 0 p[11]
port 8 nsew signal input
flabel metal2 s 774 5620 974 5740 0 FreeSans 250 0 0 0 p[8]
port 19 nsew signal input
flabel metal2 s 1436 6670 1636 6790 0 FreeSans 250 0 0 0 b[3]
port 5 nsew signal tristate
flabel metal3 s 810 4096 1010 4196 0 FreeSans 250 0 0 0 p[13]
port 10 nsew signal input
flabel metal3 s 6056 2842 6856 2962 0 FreeSans 250 0 0 0 b[1]
port 3 nsew signal tristate
flabel metal1 s 784 2974 984 3074 0 FreeSans 250 0 0 0 p[10]
port 7 nsew signal input
flabel metal2 s 1400 1772 1456 1972 0 FreeSans 224 90 0 0 p[0]
port 6 nsew signal input
flabel metal2 s 2040 1798 2096 1998 0 FreeSans 250 90 0 0 p[1]
port 12 nsew signal input
flabel metal2 s 2684 1804 2740 2004 0 FreeSans 250 90 0 0 p[2]
port 13 nsew signal input
flabel metal2 s 3324 1802 3380 2002 0 FreeSans 250 90 0 0 p[3]
port 14 nsew signal input
flabel metal2 s 4158 1810 4214 2010 0 FreeSans 250 90 0 0 p[7]
port 18 nsew signal input
flabel metal2 s 4616 1814 4672 2014 0 FreeSans 250 90 0 0 p[6]
port 17 nsew signal input
flabel metal2 s 5166 1806 5222 2006 0 FreeSans 250 90 0 0 p[5]
port 16 nsew signal input
flabel metal2 s 5808 1818 5864 2018 0 FreeSans 250 90 0 0 p[4]
port 15 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 7058 9202
<< end >>
