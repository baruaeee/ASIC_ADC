magic
tech sky130A
timestamp 1696190656
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 Vin
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 Vout
port 1 nsew
<< end >>
