magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< nwell >>
rect -1576 -261 1576 261
<< pmos >>
rect -1380 -42 1380 42
<< pdiff >>
rect -1438 30 -1380 42
rect -1438 -30 -1426 30
rect -1392 -30 -1380 30
rect -1438 -42 -1380 -30
rect 1380 30 1438 42
rect 1380 -30 1392 30
rect 1426 -30 1438 30
rect 1380 -42 1438 -30
<< pdiffc >>
rect -1426 -30 -1392 30
rect 1392 -30 1426 30
<< nsubdiff >>
rect -1540 191 -1444 225
rect 1444 191 1540 225
rect -1540 129 -1506 191
rect 1506 129 1540 191
rect -1540 -191 -1506 -129
rect 1506 -191 1540 -129
rect -1540 -225 -1444 -191
rect 1444 -225 1540 -191
<< nsubdiffcont >>
rect -1444 191 1444 225
rect -1540 -129 -1506 129
rect 1506 -129 1540 129
rect -1444 -225 1444 -191
<< poly >>
rect -1380 123 1380 139
rect -1380 89 -1364 123
rect 1364 89 1380 123
rect -1380 42 1380 89
rect -1380 -89 1380 -42
rect -1380 -123 -1364 -89
rect 1364 -123 1380 -89
rect -1380 -139 1380 -123
<< polycont >>
rect -1364 89 1364 123
rect -1364 -123 1364 -89
<< locali >>
rect -1540 191 -1444 225
rect 1444 191 1540 225
rect -1540 129 -1506 191
rect 1506 129 1540 191
rect -1380 89 -1364 123
rect 1364 89 1380 123
rect -1426 30 -1392 46
rect -1426 -46 -1392 -30
rect 1392 30 1426 46
rect 1392 -46 1426 -30
rect -1380 -123 -1364 -89
rect 1364 -123 1380 -89
rect -1540 -191 -1506 -129
rect 1506 -191 1540 -129
rect -1540 -225 -1444 -191
rect 1444 -225 1540 -191
<< viali >>
rect -1364 89 1364 123
rect -1426 -30 -1392 30
rect 1392 -30 1426 30
rect -1364 -123 1364 -89
<< metal1 >>
rect -1376 123 1376 129
rect -1376 89 -1364 123
rect 1364 89 1376 123
rect -1376 83 1376 89
rect -1432 30 -1386 42
rect -1432 -30 -1426 30
rect -1392 -30 -1386 30
rect -1432 -42 -1386 -30
rect 1386 30 1432 42
rect 1386 -30 1392 30
rect 1426 -30 1432 30
rect 1386 -42 1432 -30
rect -1376 -89 1376 -83
rect -1376 -123 -1364 -89
rect 1364 -123 1376 -89
rect -1376 -129 1376 -123
<< properties >>
string FIXED_BBOX -1523 -208 1523 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 13.8 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
