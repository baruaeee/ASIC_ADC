magic
tech sky130A
magscale 1 2
timestamp 1706480381
<< pwell >>
rect 744 -972 870 -938
<< locali >>
rect 537 356 540 390
rect 504 336 540 356
rect 1184 -1008 1244 -862
<< viali >>
rect 503 356 537 390
rect 1166 352 1201 387
<< metal1 >>
rect 497 390 543 402
rect 497 356 503 390
rect 537 356 543 390
rect 1152 393 1202 394
rect 1420 393 1520 394
rect 1152 387 1520 393
rect 1152 385 1166 387
rect 497 344 543 356
rect 1151 352 1166 385
rect 1201 352 1520 387
rect 1151 351 1520 352
rect 1152 348 1207 351
rect 1160 346 1207 348
rect 501 -336 535 344
rect 571 144 577 196
rect 629 144 650 196
rect 576 134 650 144
rect 983 181 1018 199
rect 983 146 1104 181
rect 983 133 1018 146
rect 768 50 880 76
rect 768 30 800 50
rect 794 -2 800 30
rect 852 30 880 50
rect 852 -2 858 30
rect 1068 -196 1103 146
rect 1161 96 1195 346
rect 1274 292 1338 298
rect 1420 294 1520 351
rect 1274 244 1340 292
rect 1278 242 1340 244
rect 1245 96 1279 149
rect 1161 61 1279 96
rect 1245 -15 1279 61
rect 1333 95 1367 157
rect 1333 61 1513 95
rect 1333 -47 1367 61
rect 1278 -147 1334 -136
rect 1278 -172 1339 -147
rect 1278 -196 1280 -172
rect 1068 -224 1280 -196
rect 1332 -224 1339 -172
rect 1068 -231 1339 -224
rect 1479 -326 1513 61
rect 500 -445 535 -336
rect 894 -388 910 -336
rect 962 -388 968 -336
rect 1418 -358 1518 -326
rect 894 -394 952 -388
rect 1197 -392 1518 -358
rect 500 -479 779 -445
rect 1197 -501 1231 -392
rect 1418 -426 1518 -392
rect 1179 -535 1243 -501
rect 1099 -650 1133 -587
rect 688 -656 1133 -650
rect 688 -684 886 -656
rect 492 -700 592 -688
rect 492 -704 642 -700
rect 492 -708 646 -704
rect 689 -705 823 -684
rect 880 -708 886 -684
rect 938 -684 1133 -656
rect 1296 -626 1370 -618
rect 1296 -678 1319 -626
rect 1371 -678 1377 -626
rect 1296 -684 1370 -678
rect 938 -708 944 -684
rect 492 -760 582 -708
rect 634 -760 646 -708
rect 492 -764 646 -760
rect 492 -766 642 -764
rect 492 -788 592 -766
rect 691 -798 995 -764
rect 724 -942 730 -890
rect 782 -942 788 -890
rect 961 -944 995 -798
rect 1099 -799 1133 -684
rect 1181 -895 1245 -861
rect 961 -973 1062 -944
rect 1211 -973 1245 -895
rect 961 -1007 1245 -973
rect 962 -1044 1062 -1007
<< via1 >>
rect 577 144 629 196
rect 800 -2 852 50
rect 1280 -224 1332 -172
rect 910 -388 962 -336
rect 886 -708 938 -656
rect 1319 -678 1371 -626
rect 582 -760 634 -708
rect 730 -942 782 -890
<< metal2 >>
rect 577 196 629 202
rect 577 138 629 144
rect 586 -135 620 138
rect 800 50 852 56
rect 800 -8 852 -2
rect 809 -53 843 -8
rect 809 -87 1028 -53
rect 586 -169 953 -135
rect 919 -330 953 -169
rect 910 -336 962 -330
rect 910 -394 962 -388
rect 994 -559 1028 -87
rect 1274 -224 1280 -172
rect 1332 -181 1338 -172
rect 1332 -224 1362 -181
rect 591 -593 1028 -559
rect 591 -702 625 -593
rect 1328 -620 1362 -224
rect 1319 -626 1371 -620
rect 886 -656 938 -650
rect 582 -708 634 -702
rect 1319 -684 1371 -678
rect 886 -714 938 -708
rect 582 -766 634 -760
rect 730 -890 782 -884
rect 895 -938 929 -714
rect 782 -942 929 -938
rect 730 -948 929 -942
rect 739 -972 929 -948
use sky130_fd_pr__nfet_01v8_D7Y3TR  XM0
timestamp 1706211875
transform 0 -1 753 1 0 -781
box -263 -285 263 285
use sky130_fd_pr__pfet_01v8_2ZD99F  XM1
timestamp 1706480381
transform 1 0 819 0 1 165
box -349 -261 349 261
use sky130_fd_pr__nfet_01v8_2BW22M  XM2
timestamp 1706204487
transform 1 0 728 0 1 -364
box -350 -252 350 252
use sky130_fd_pr__pfet_01v8_XJP3BL  XM3
timestamp 1706204487
transform 1 0 1307 0 -1 53
box -211 -369 211 369
use sky130_fd_pr__nfet_01v8_LH5FDA  XM4
timestamp 1706211875
transform 0 -1 1214 -1 0 -698
box -260 -252 346 252
<< labels >>
flabel metal1 1418 -426 1518 -326 0 FreeSans 256 0 0 0 V02
port 2 nsew
flabel metal1 962 -1044 1062 -944 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 492 -788 592 -688 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 1420 294 1520 394 0 FreeSans 256 0 0 0 Vp
port 0 nsew
<< end >>
