magic
tech sky130A
magscale 1 2
timestamp 1704962958
<< nwell >>
rect -492 -261 492 261
<< pmos >>
rect -296 -42 296 42
<< pdiff >>
rect -354 30 -296 42
rect -354 -30 -342 30
rect -308 -30 -296 30
rect -354 -42 -296 -30
rect 296 30 354 42
rect 296 -30 308 30
rect 342 -30 354 30
rect 296 -42 354 -30
<< pdiffc >>
rect -342 -30 -308 30
rect 308 -30 342 30
<< nsubdiff >>
rect -456 191 -360 225
rect 360 191 456 225
rect -456 129 -422 191
rect 422 129 456 191
rect -456 -191 -422 -129
rect 422 -191 456 -129
rect -456 -225 -360 -191
rect 360 -225 456 -191
<< nsubdiffcont >>
rect -360 191 360 225
rect -456 -129 -422 129
rect 422 -129 456 129
rect -360 -225 360 -191
<< poly >>
rect -296 123 296 139
rect -296 89 -280 123
rect 280 89 296 123
rect -296 42 296 89
rect -296 -89 296 -42
rect -296 -123 -280 -89
rect 280 -123 296 -89
rect -296 -139 296 -123
<< polycont >>
rect -280 89 280 123
rect -280 -123 280 -89
<< locali >>
rect -456 191 -360 225
rect 360 191 456 225
rect -456 129 -422 191
rect 422 129 456 191
rect -296 89 -280 123
rect 280 89 296 123
rect -342 30 -308 46
rect -342 -46 -308 -30
rect 308 30 342 46
rect 308 -46 342 -30
rect -296 -123 -280 -89
rect 280 -123 296 -89
rect -456 -191 -422 -129
rect 422 -191 456 -129
rect -456 -225 -360 -191
rect 360 -225 456 -191
<< viali >>
rect -280 89 280 123
rect -342 -30 -308 30
rect 308 -30 342 30
rect -280 -123 280 -89
<< metal1 >>
rect -292 123 292 129
rect -292 89 -280 123
rect 280 89 292 123
rect -292 83 292 89
rect -348 30 -302 42
rect -348 -30 -342 30
rect -308 -30 -302 30
rect -348 -42 -302 -30
rect 302 30 348 42
rect 302 -30 308 30
rect 342 -30 348 30
rect 302 -42 348 -30
rect -292 -89 292 -83
rect -292 -123 -280 -89
rect 280 -123 292 -89
rect -292 -129 292 -123
<< properties >>
string FIXED_BBOX -439 -208 439 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 2.96 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
