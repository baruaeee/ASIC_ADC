magic
tech sky130A
magscale 1 2
timestamp 1706548588
<< nwell >>
rect 9392 560 9464 580
<< metal1 >>
rect 5350 6782 5450 6882
rect 4177 6643 4320 6702
rect 4177 6598 4236 6643
rect 4154 6498 4254 6598
rect 1535 6285 1541 6337
rect 1593 6285 1599 6337
rect 1710 4885 1762 4891
rect 1710 4826 1762 4832
rect 2924 3734 2930 3786
rect 2982 3734 2988 3786
rect 4140 2414 4388 2462
rect 5490 2120 5542 2126
rect 4873 2075 5490 2109
rect 1799 1487 1833 2057
rect 3558 1580 3610 1586
rect 3495 1537 3558 1571
rect 3495 1487 3529 1537
rect 3558 1522 3610 1528
rect 1799 1453 3529 1487
rect 4873 1365 4907 2075
rect 5490 2058 5542 2064
rect 5966 1546 5972 1598
rect 6024 1546 6030 1598
rect 4753 1331 4907 1365
rect 6917 1323 6923 1375
rect 6975 1323 6981 1375
rect 8721 1193 8773 1199
rect 8721 1135 8773 1141
rect 7797 1037 7803 1089
rect 7855 1037 7861 1089
rect 9944 1080 9996 1086
rect 9944 1018 9996 1024
rect 5663 609 5697 687
rect 5802 609 5902 646
rect 5663 575 5902 609
rect 5802 546 5902 575
rect 2659 421 2711 427
rect 2659 363 2711 369
<< via1 >>
rect 1541 6285 1593 6337
rect 1710 4832 1762 4885
rect 2930 3734 2982 3786
rect 3558 1528 3610 1580
rect 5490 2064 5542 2120
rect 5972 1546 6024 1598
rect 6923 1323 6975 1375
rect 8721 1141 8773 1193
rect 7803 1037 7855 1089
rect 9944 1024 9996 1080
rect 2659 369 2711 421
<< metal2 >>
rect 1434 7053 5555 7106
rect 1434 4885 1487 7053
rect 1543 6950 5278 6997
rect 1543 6343 1590 6950
rect 5231 6651 5278 6950
rect 5502 6793 5555 7053
rect 5502 6740 7595 6793
rect 1541 6337 1593 6343
rect 1541 6279 1593 6285
rect 5088 5592 5144 5601
rect 5088 5527 5144 5536
rect 1434 4832 1710 4885
rect 1762 4832 1768 4885
rect 2919 3768 2928 3824
rect 2984 3768 2993 3824
rect 2930 3728 2982 3734
rect 5484 2064 5490 2120
rect 5542 2064 5752 2120
rect 5858 2060 6070 2108
rect 5858 1996 5906 2060
rect 6434 2054 6677 2103
rect 7107 2079 7417 2129
rect 9016 2104 9401 2153
rect 6434 2019 6483 2054
rect 4368 1948 5906 1996
rect 5962 1970 6483 2019
rect 7107 2009 7157 2079
rect 7739 2057 7950 2104
rect 7739 2032 7786 2057
rect 4368 1626 4416 1948
rect 5962 1897 6011 1970
rect 6535 1959 7157 2009
rect 7219 1985 7786 2032
rect 8570 2042 8811 2091
rect 8570 2015 8619 2042
rect 6535 1935 6585 1959
rect 3552 1528 3558 1580
rect 3610 1578 3616 1580
rect 3838 1578 4416 1626
rect 4966 1848 6011 1897
rect 6053 1885 6585 1935
rect 7219 1908 7266 1985
rect 7850 1966 8619 2015
rect 9016 1991 9065 2104
rect 7850 1937 7899 1966
rect 3610 1530 3886 1578
rect 3610 1528 3616 1530
rect 4966 1295 5015 1848
rect 6053 1749 6103 1885
rect 5973 1699 6103 1749
rect 6925 1861 7266 1908
rect 7804 1888 7899 1937
rect 8754 1942 9065 1991
rect 5973 1604 6023 1699
rect 5972 1598 6024 1604
rect 5972 1540 6024 1546
rect 6925 1381 6972 1861
rect 6923 1375 6975 1381
rect 6923 1317 6975 1323
rect 4888 1246 5015 1295
rect 4888 753 4937 1246
rect 7804 1095 7853 1888
rect 8754 1193 8803 1942
rect 8715 1141 8721 1193
rect 8773 1142 8803 1193
rect 8773 1141 8779 1142
rect 7803 1089 7855 1095
rect 10052 1080 10108 2156
rect 7803 1031 7855 1037
rect 9938 1024 9944 1080
rect 9996 1024 10108 1080
rect 4766 704 4937 753
rect 2653 369 2659 421
rect 2711 419 2717 421
rect 4766 419 4815 704
rect 2711 370 4815 419
rect 2711 369 2717 370
<< via2 >>
rect 5088 5536 5144 5592
rect 2928 3786 2984 3824
rect 2928 3768 2930 3786
rect 2930 3768 2982 3786
rect 2982 3768 2984 3786
<< metal3 >>
rect 3526 5626 4550 5686
rect 3526 5092 3586 5626
rect 4490 5594 4550 5626
rect 5083 5594 5149 5597
rect 4490 5592 5149 5594
rect 4490 5536 5088 5592
rect 5144 5536 5149 5592
rect 4490 5534 5149 5536
rect 5083 5531 5149 5534
rect 3210 5032 3586 5092
rect 3210 3956 3270 5032
rect 2926 3896 3270 3956
rect 2926 3829 2986 3896
rect 2923 3824 2989 3829
rect 2923 3768 2928 3824
rect 2984 3768 2989 3824
rect 2923 3763 2989 3768
use therm  therm_0
timestamp 1706543737
transform 1 0 4297 0 1 72
box -111 1962 7123 6724
use Analog  x1
timestamp 1706548588
transform 1 0 0 0 1 7400
box 1538 -7112 10018 -488
<< labels >>
flabel metal1 5350 6782 5450 6882 0 FreeSans 256 180 0 0 Vn
port 17 nsew
flabel metal1 4154 6498 4254 6598 0 FreeSans 256 180 0 0 Vin
port 1 nsew
flabel metal1 5802 546 5902 646 0 FreeSans 256 180 0 0 Vp
port 0 nsew
<< end >>
