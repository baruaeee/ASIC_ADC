magic
tech sky130A
magscale 1 2
timestamp 1704332234
<< locali >>
rect 456 930 592 998
rect 378 736 474 772
rect 378 -20 414 736
rect 940 308 1084 402
rect 1276 132 1356 168
rect 378 -56 490 -20
rect 1320 -434 1356 132
<< viali >>
rect 1320 -470 1356 -434
<< metal1 >>
rect 782 1304 982 1464
rect 505 1266 982 1304
rect 505 1007 543 1266
rect 782 1264 982 1266
rect 584 1042 650 1100
rect 906 1009 944 1264
rect 505 933 587 1007
rect 645 919 734 1007
rect 906 923 1009 1009
rect 1132 930 1421 968
rect 174 838 651 876
rect 696 871 734 919
rect 1022 871 1122 878
rect 174 732 212 838
rect 696 833 1123 871
rect 1383 838 1421 930
rect 160 532 360 732
rect 696 698 734 833
rect 1022 826 1122 833
rect 509 660 734 698
rect 174 261 212 532
rect 509 417 547 660
rect 1083 479 1121 826
rect 1383 638 1584 838
rect 1083 441 1147 479
rect 509 389 565 417
rect 509 303 597 389
rect 717 301 806 393
rect 1383 383 1421 638
rect 1143 345 1421 383
rect 174 223 697 261
rect 552 -224 588 -164
rect 768 -171 806 301
rect 1082 214 1148 276
rect 718 -224 754 -222
rect 1080 -224 1116 -166
rect 552 -260 1116 -224
rect 718 -442 754 -260
rect 1308 -434 1368 -428
rect 1308 -436 1320 -434
rect 1002 -442 1320 -436
rect 718 -470 1320 -442
rect 1356 -470 1368 -434
rect 718 -472 1368 -470
rect 718 -478 1202 -472
rect 1308 -476 1368 -472
rect 1002 -636 1202 -478
use sky130_fd_pr__pfet_01v8_XGAKDL  XM0
timestamp 1704331930
transform 0 -1 835 1 0 -195
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_ZFH27D  XM1
timestamp 1704331930
transform 1 0 660 0 1 348
box -246 -252 246 252
use sky130_fd_pr__pfet_01v8_E7ZT25  XM2
timestamp 1704331930
transform 1 0 617 0 1 964
box -211 -262 211 262
use sky130_fd_pr__pfet_01v8_JM8GTH  XM3
timestamp 1704331930
transform 1 0 1072 0 1 965
box -246 -261 246 261
use sky130_fd_pr__nfet_01v8_L9ESAD  XM4
timestamp 1704331930
transform 1 0 1115 0 1 356
box -211 -260 211 260
<< labels >>
flabel metal1 782 1264 982 1464 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 1384 638 1584 838 0 FreeSans 256 0 0 0 V11
port 1 nsew
flabel metal1 160 532 360 732 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 1002 -636 1202 -436 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
