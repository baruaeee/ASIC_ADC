magic
tech sky130A
magscale 1 2
timestamp 1704877912
<< nwell >>
rect -291 -261 291 261
<< pmos >>
rect -95 -42 95 42
<< pdiff >>
rect -153 30 -95 42
rect -153 -30 -141 30
rect -107 -30 -95 30
rect -153 -42 -95 -30
rect 95 30 153 42
rect 95 -30 107 30
rect 141 -30 153 30
rect 95 -42 153 -30
<< pdiffc >>
rect -141 -30 -107 30
rect 107 -30 141 30
<< nsubdiff >>
rect -255 191 -159 225
rect 159 191 255 225
rect -255 129 -221 191
rect 221 129 255 191
rect -255 -191 -221 -129
rect 221 -191 255 -129
rect -255 -225 -159 -191
rect 159 -225 255 -191
<< nsubdiffcont >>
rect -159 191 159 225
rect -255 -129 -221 129
rect 221 -129 255 129
rect -159 -225 159 -191
<< poly >>
rect -95 123 95 139
rect -95 89 -79 123
rect 79 89 95 123
rect -95 42 95 89
rect -95 -89 95 -42
rect -95 -123 -79 -89
rect 79 -123 95 -89
rect -95 -139 95 -123
<< polycont >>
rect -79 89 79 123
rect -79 -123 79 -89
<< locali >>
rect -255 191 -159 225
rect 159 191 255 225
rect -255 129 -221 191
rect 221 129 255 191
rect -95 89 -79 123
rect 79 89 95 123
rect -141 30 -107 46
rect -141 -46 -107 -30
rect 107 30 141 46
rect 107 -46 141 -30
rect -95 -123 -79 -89
rect 79 -123 95 -89
rect -255 -191 -221 -129
rect 221 -191 255 -129
rect -255 -225 -159 -191
rect 159 -225 255 -191
<< viali >>
rect -79 89 79 123
rect -141 -30 -107 30
rect 107 -30 141 30
rect -79 -123 79 -89
<< metal1 >>
rect -91 123 91 129
rect -91 89 -79 123
rect 79 89 91 123
rect -91 83 91 89
rect -147 30 -101 42
rect -147 -30 -141 30
rect -107 -30 -101 30
rect -147 -42 -101 -30
rect 101 30 147 42
rect 101 -30 107 30
rect 141 -30 147 30
rect 101 -42 147 -30
rect -91 -89 91 -83
rect -91 -123 -79 -89
rect 79 -123 91 -89
rect -91 -129 91 -123
<< properties >>
string FIXED_BBOX -238 -208 238 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.422 l 0.946 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
