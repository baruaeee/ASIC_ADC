.subckt analog_therm b0 Vin b1 b2 b3 Vp Vn
x0 p10 VGND VNB VPB VPWR 1 sky130_fd_sc_hd__clkinv_1
x1 p1 p0 VGND VNB VPB VPWR 2 sky130_fd_sc_hd__nand2_1
x2 p1 p0 p2 VGND VNB VPB VPWR 3 sky130_fd_sc_hd__nand3_1
x3 p1 p0 p3 p2 VGND VNB VPB VPWR 4 sky130_fd_sc_hd__nand4_1
x4 p5 p4 VGND VNB VPB VPWR 5 sky130_fd_sc_hd__nand2_1
x5 p5 p4 p7 p6 VGND VNB VPB VPWR 6 sky130_fd_sc_hd__nand4_1
x6 4 6 VGND VNB VPB VPWR 7 sky130_fd_sc_hd__nor2_1
x7 p8 p9 VGND VNB VPB VPWR 8 sky130_fd_sc_hd__nand2_1
x8 p11 p10 VGND VNB VPB VPWR 9 sky130_fd_sc_hd__nand2_1
x9 4 6 8 9 VGND VNB VPB VPWR 10 sky130_fd_sc_hd__nor4_1
x10 p13 p12 VGND VNB VPB VPWR 11 sky130_fd_sc_hd__and2_0
x11 10 11 VGND VNB VPB VPWR 12 sky130_fd_sc_hd__nand2_1
x12 p14 10 11 VGND VNB VPB VPWR 13 sky130_fd_sc_hd__nand3_1
x13 p7 5 VGND VNB VPB VPWR 14 sky130_fd_sc_hd__nor2_1
x14 p5 p7 p6 VGND VNB VPB VPWR 15 sky130_fd_sc_hd__nor3_1
x15 p6 14 15 p4 VGND VNB VPB VPWR 16 sky130_fd_sc_hd__a22oi_1
x16 p13 p14 VGND VNB VPB VPWR 17 sky130_fd_sc_hd__nor2_1
x17 p13 p12 p14 VGND VNB VPB VPWR 18 sky130_fd_sc_hd__or3_1
x18 p11 p10 VGND VNB VPB VPWR 19 sky130_fd_sc_hd__lpflow_inputiso1p_1
x19 p8 p9 18 19 VGND VNB VPB VPWR 20 sky130_fd_sc_hd__nor4_1
x20 4 20 VGND VNB VPB VPWR 21 sky130_fd_sc_hd__nand2b_1
x21 p9 18 19 p8 VGND VNB VPB VPWR 22 sky130_fd_sc_hd__nor4b_1
x22 p11 8 18 VGND VNB VPB VPWR 23 sky130_fd_sc_hd__nor3_1
x23 p11 1 8 18 VGND VNB VPB VPWR 24 sky130_fd_sc_hd__nor4_1
x24 22 24 7 VGND VNB VPB VPWR 25 sky130_fd_sc_hd__o21ai_0
x25 p1 p2 p0 VGND VNB VPB VPWR 26 sky130_fd_sc_hd__or3b_1
x26 p5 p4 p7 p6 VGND VNB VPB VPWR 27 sky130_fd_sc_hd__or4_1
x27 3 26 27 p3 VGND VNB VPB VPWR 28 sky130_fd_sc_hd__a211oi_1
x28 p12 10 17 20 28 VGND VNB VPB VPWR 29 sky130_fd_sc_hd__a32oi_1
x29 16 21 25 29 13 VGND VNB VPB VPWR b0 sky130_fd_sc_hd__o2111ai_1
x30 4 14 20 VGND VNB VPB VPWR 30 sky130_fd_sc_hd__nand3b_1
x31 7 23 VGND VNB VPB VPWR 31 sky130_fd_sc_hd__nand2_1
x32 p3 2 27 VGND VNB VPB VPWR 32 sky130_fd_sc_hd__nor3_1
x33 20 32 VGND VNB VPB VPWR 33 sky130_fd_sc_hd__nand2_1
x34 12 30 31 33 VGND VNB VPB VPWR b1 sky130_fd_sc_hd__nand4_1
x35 11 17 10 VGND VNB VPB VPWR 34 sky130_fd_sc_hd__o21ai_0
x36 14 15 VGND VNB VPB VPWR 35 sky130_fd_sc_hd__nor2_1
x37 21 35 34 VGND VNB VPB VPWR b2 sky130_fd_sc_hd__o21ai_0
x38 20 22 23 7 VGND VNB VPB VPWR 36 sky130_fd_sc_hd__o31ai_1
x39 34 36 VGND VNB VPB VPWR b3 sky130_fd_sc_hd__nand2_1
x40 Vp Vin p0 p1 p2 p3 p4 p5 p6 p7 p8 p9 p10 p11 p12 p13 p14 Vn Analog
.ends
