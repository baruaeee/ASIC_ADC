magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 150 29 156
rect -29 116 -17 150
rect -29 110 29 116
rect -29 -116 29 -110
rect -29 -150 -17 -116
rect -29 -156 29 -150
<< nwell >>
rect -211 -288 211 288
<< pmos >>
rect -15 -69 15 69
<< pdiff >>
rect -73 57 -15 69
rect -73 -57 -61 57
rect -27 -57 -15 57
rect -73 -69 -15 -57
rect 15 57 73 69
rect 15 -57 27 57
rect 61 -57 73 57
rect 15 -69 73 -57
<< pdiffc >>
rect -61 -57 -27 57
rect 27 -57 61 57
<< nsubdiff >>
rect -175 218 -79 252
rect 79 218 175 252
rect -175 156 -141 218
rect 141 156 175 218
rect -175 -218 -141 -156
rect 141 -218 175 -156
rect -175 -252 -79 -218
rect 79 -252 175 -218
<< nsubdiffcont >>
rect -79 218 79 252
rect -175 -156 -141 156
rect 141 -156 175 156
rect -79 -252 79 -218
<< poly >>
rect -33 150 33 166
rect -33 116 -17 150
rect 17 116 33 150
rect -33 100 33 116
rect -15 69 15 100
rect -15 -100 15 -69
rect -33 -116 33 -100
rect -33 -150 -17 -116
rect 17 -150 33 -116
rect -33 -166 33 -150
<< polycont >>
rect -17 116 17 150
rect -17 -150 17 -116
<< locali >>
rect -175 218 -79 252
rect 79 218 175 252
rect -175 156 -141 218
rect 141 156 175 218
rect -33 116 -17 150
rect 17 116 33 150
rect -61 57 -27 73
rect -61 -73 -27 -57
rect 27 57 61 73
rect 27 -73 61 -57
rect -33 -150 -17 -116
rect 17 -150 33 -116
rect -175 -218 -141 -156
rect 141 -218 175 -156
rect -175 -252 -79 -218
rect 79 -252 175 -218
<< viali >>
rect -17 116 17 150
rect -61 -57 -27 57
rect 27 -57 61 57
rect -17 -150 17 -116
<< metal1 >>
rect -29 150 29 156
rect -29 116 -17 150
rect 17 116 29 150
rect -29 110 29 116
rect -67 57 -21 69
rect -67 -57 -61 57
rect -27 -57 -21 57
rect -67 -69 -21 -57
rect 21 57 67 69
rect 21 -57 27 57
rect 61 -57 67 57
rect 21 -69 67 -57
rect -29 -116 29 -110
rect -29 -150 -17 -116
rect 17 -150 29 -116
rect -29 -156 29 -150
<< properties >>
string FIXED_BBOX -158 -235 158 235
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.69 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
