magic
tech sky130A
magscale 1 2
timestamp 1705440136
<< locali >>
rect 1026 256 1088 347
rect 1250 -98 1312 -26
rect 1224 -556 1458 -494
rect 1628 -808 1778 -748
rect 1016 -902 1112 -840
<< viali >>
rect 1026 347 1089 410
rect 1249 -162 1313 -98
rect 1112 -903 1176 -839
<< metal1 >>
rect 692 410 892 556
rect 1014 410 1101 416
rect 1192 410 1635 463
rect 692 356 1026 410
rect 0 0 200 200
rect 720 144 783 356
rect 841 347 1026 356
rect 1089 400 1635 410
rect 1089 347 1255 400
rect 1572 367 1635 400
rect 1014 341 1101 347
rect 350 78 627 141
rect 0 -400 200 -200
rect 350 -490 413 78
rect 764 -65 827 89
rect 1690 86 1952 150
rect 1566 -52 1630 -48
rect 547 -76 969 -65
rect 547 -128 903 -76
rect 547 -314 610 -128
rect 966 -128 969 -76
rect 1237 -98 1325 -92
rect 903 -146 966 -140
rect 1237 -162 1249 -98
rect 1313 -162 1325 -98
rect 1566 -112 1644 -52
rect 1888 -56 1952 86
rect 1237 -168 1325 -162
rect 546 -454 610 -314
rect 1098 -440 1200 -376
rect 246 -494 446 -490
rect 246 -558 872 -494
rect 0 -800 200 -600
rect 246 -690 446 -558
rect 1136 -706 1200 -440
rect 724 -770 1200 -706
rect 410 -998 626 -954
rect 724 -958 788 -770
rect 1106 -839 1182 -827
rect 1252 -839 1316 -168
rect 1580 -270 1644 -112
rect 1882 -120 1888 -56
rect 1952 -120 1958 -56
rect 1384 -334 1954 -270
rect 1384 -744 1448 -334
rect 1890 -416 1954 -334
rect 1862 -616 2062 -416
rect 1384 -808 1574 -744
rect 1106 -903 1112 -839
rect 1176 -903 1316 -839
rect 1106 -915 1182 -903
rect 1628 -920 1854 -856
rect 0 -1200 200 -1000
rect 240 -1010 626 -998
rect 240 -1074 1192 -1010
rect 240 -1198 440 -1074
rect 1128 -1136 1192 -1074
rect 1364 -1088 1370 -1024
rect 1434 -1026 1440 -1024
rect 1434 -1088 1634 -1026
rect 1366 -1092 1634 -1088
rect 1790 -1136 1854 -920
rect 1128 -1200 1854 -1136
<< via1 >>
rect 903 -140 966 -76
rect 1888 -120 1952 -56
rect 1370 -1088 1434 -1024
<< metal2 >>
rect 1888 -56 1952 -50
rect 897 -140 903 -76
rect 966 -140 1434 -76
rect 1370 -236 1434 -140
rect 1888 -236 1952 -120
rect 1370 -300 1952 -236
rect 1370 -1024 1434 -300
rect 1370 -1094 1434 -1088
use sky130_fd_pr__pfet_01v8_XGS3BL  XM0
timestamp 1704310947
transform 0 1 765 -1 0 -987
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_L6G859  XM1
timestamp 1704310896
transform 1 0 872 0 1 -412
box -426 -252 426 252
use sky130_fd_pr__pfet_01v8_XW9KDL  XM2
timestamp 1704311015
transform 0 -1 897 1 0 115
box -211 -449 211 449
use sky130_fd_pr__pfet_01v8_VZ9GC6  XM3
timestamp 1704310896
transform 0 1 1601 -1 0 160
box -396 -261 396 261
use sky130_fd_pr__nfet_01v8_ATLS57  XM4
timestamp 1704311096
transform -1 0 1599 0 -1 -784
box -211 -410 211 410
<< labels >>
flabel metal1 240 -1198 440 -998 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 692 356 892 556 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 246 -690 446 -490 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 1862 -616 2062 -416 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
<< end >>
