* NGSPICE file created from analog_therm.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X a_208_47# a_75_199#
+ a_544_297# a_315_47# a_201_297#
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_208_47# X 1.91e-19
C1 a_544_297# X 2.35e-19
C2 VPB C1 0.0394f
C3 a_201_297# X 0.0131f
C4 A2 A1 0.0689f
C5 a_75_199# X 0.0959f
C6 VGND C1 0.0181f
C7 A2 VPWR 0.0174f
C8 a_315_47# A2 0.00335f
C9 A1 C1 3.21e-19
C10 C1 VPWR 0.0146f
C11 a_208_47# A2 0.00102f
C12 a_201_297# A2 0.0112f
C13 VPB A3 0.0268f
C14 a_75_199# A2 0.0621f
C15 VGND A3 0.0161f
C16 a_201_297# C1 0.00243f
C17 VPB B1 0.0292f
C18 a_75_199# C1 0.0628f
C19 VGND B1 0.0171f
C20 A3 VPWR 0.0181f
C21 A2 X 3.01e-19
C22 A1 B1 0.0716f
C23 C1 X 5.14e-20
C24 B1 VPWR 0.0125f
C25 a_208_47# A3 3.65e-19
C26 a_201_297# A3 0.00642f
C27 a_75_199# A3 0.163f
C28 VGND VPB 0.00772f
C29 a_544_297# B1 1.13e-19
C30 a_201_297# B1 0.00594f
C31 VPB A1 0.0306f
C32 a_75_199# B1 0.102f
C33 VGND A1 0.0113f
C34 A3 X 0.00317f
C35 VPB VPWR 0.0749f
C36 VGND VPWR 0.0735f
C37 VGND a_315_47# 0.00427f
C38 A1 VPWR 0.0151f
C39 B1 X 7.79e-20
C40 a_315_47# A1 0.00313f
C41 a_201_297# VPB 0.00186f
C42 VGND a_208_47# 0.00302f
C43 a_75_199# VPB 0.0486f
C44 VGND a_544_297# 0.00256f
C45 a_315_47# VPWR 0.00154f
C46 VGND a_201_297# 0.00403f
C47 A3 A2 0.0747f
C48 VGND a_75_199# 0.362f
C49 a_201_297# A1 0.011f
C50 a_208_47# VPWR 8.35e-19
C51 a_75_199# A1 0.0696f
C52 a_544_297# VPWR 0.0105f
C53 a_201_297# VPWR 0.211f
C54 VPB X 0.0107f
C55 a_75_199# VPWR 0.109f
C56 VGND X 0.0609f
C57 a_75_199# a_315_47# 0.0202f
C58 A1 X 1.2e-19
C59 B1 C1 0.066f
C60 a_201_297# a_544_297# 0.00702f
C61 a_75_199# a_208_47# 0.0159f
C62 a_75_199# a_544_297# 0.0176f
C63 X VPWR 0.0676f
C64 a_75_199# a_201_297# 0.16f
C65 VPB A2 0.0376f
C66 VGND A2 0.0119f
C67 VGND VNB 0.437f
C68 VPWR VNB 0.365f
C69 X VNB 0.0906f
C70 C1 VNB 0.148f
C71 B1 VNB 0.0947f
C72 A1 VNB 0.101f
C73 A2 VNB 0.11f
C74 A3 VNB 0.0908f
C75 VPB VNB 0.782f
C76 a_201_297# VNB 0.00345f
C77 a_75_199# VNB 0.205f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_181_47# a_109_47# a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_27_47# a_109_47# 0.00517f
C1 VGND a_27_47# 0.134f
C2 a_27_47# B 0.0625f
C3 X a_27_47# 0.087f
C4 C a_27_47# 0.186f
C5 VPWR a_181_47# 3.97e-19
C6 a_27_47# VPB 0.0501f
C7 VPWR A 0.0185f
C8 VGND a_181_47# 0.00261f
C9 A a_109_47# 6.45e-19
C10 C a_181_47# 0.00151f
C11 VGND A 0.0154f
C12 A B 0.0869f
C13 VPWR a_109_47# 3.29e-19
C14 VPWR VGND 0.0475f
C15 VPWR B 0.128f
C16 VPWR X 0.0766f
C17 VPWR C 0.00464f
C18 VGND a_109_47# 0.00123f
C19 VGND B 0.00714f
C20 A VPB 0.0426f
C21 X VGND 0.0708f
C22 X B 0.00111f
C23 C VGND 0.0703f
C24 C B 0.0746f
C25 C X 0.0149f
C26 a_27_47# a_181_47# 0.00401f
C27 VPWR VPB 0.0795f
C28 A a_27_47# 0.157f
C29 VGND VPB 0.00604f
C30 VPB B 0.0836f
C31 X VPB 0.0121f
C32 C VPB 0.0347f
C33 VPWR a_27_47# 0.145f
C34 VGND VNB 0.3f
C35 X VNB 0.0923f
C36 C VNB 0.12f
C37 A VNB 0.174f
C38 VPWR VNB 0.274f
C39 B VNB 0.102f
C40 VPB VNB 0.516f
C41 a_27_47# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
C0 VGND VPWR 0.353f
C1 VPWR VPB 0.0625f
C2 VGND VPB 0.0797f
C3 VPWR VNB 0.47f
C4 VGND VNB 0.427f
C5 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VGND VPWR 0.546f
C1 VPWR VPB 0.0787f
C2 VGND VPB 0.116f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_384_47# a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
C0 X VPWR 0.0847f
C1 B1 X 3.04e-20
C2 VPB X 0.0108f
C3 VPWR A2 0.0201f
C4 A1 A2 0.0921f
C5 A2 a_299_297# 0.0468f
C6 VPB A2 0.0373f
C7 X a_81_21# 0.112f
C8 A2 a_81_21# 7.47e-19
C9 a_384_47# VGND 0.00366f
C10 VPWR VGND 0.0579f
C11 A1 VGND 0.0786f
C12 VGND a_299_297# 0.00772f
C13 B1 VGND 0.0181f
C14 VPB VGND 0.00713f
C15 a_384_47# VPWR 4.08e-19
C16 a_384_47# A1 0.00884f
C17 a_384_47# a_299_297# 1.48e-19
C18 A1 VPWR 0.0209f
C19 VPWR a_299_297# 0.202f
C20 B1 VPWR 0.0196f
C21 VPB VPWR 0.068f
C22 A1 a_299_297# 0.0585f
C23 B1 A1 0.0817f
C24 B1 a_299_297# 0.00863f
C25 VPB A1 0.0264f
C26 VPB a_299_297# 0.0111f
C27 VPB B1 0.0387f
C28 VGND a_81_21# 0.173f
C29 a_384_47# a_81_21# 0.00138f
C30 VPWR a_81_21# 0.146f
C31 A1 a_81_21# 0.0568f
C32 X VGND 0.0512f
C33 a_81_21# a_299_297# 0.0821f
C34 B1 a_81_21# 0.148f
C35 VPB a_81_21# 0.0593f
C36 VGND A2 0.0495f
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 Y VGND 0.155f
C1 A Y 0.0894f
C2 VPB Y 0.0061f
C3 VGND VPWR 0.0423f
C4 A VPWR 0.0631f
C5 VPB VPWR 0.0521f
C6 Y VPWR 0.209f
C7 A VGND 0.0638f
C8 VPB VGND 0.00649f
C9 VPB A 0.0742f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X a_29_53# a_183_297# a_111_297#
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 VPB VPWR 0.0649f
C1 VPB X 0.0109f
C2 a_29_53# VPB 0.0491f
C3 VGND B 0.0152f
C4 VPB A 0.0377f
C5 C VGND 0.0161f
C6 VGND VPWR 0.0459f
C7 a_183_297# VGND 5.75e-19
C8 C B 0.0802f
C9 VGND X 0.036f
C10 a_111_297# VGND 3.96e-19
C11 a_29_53# VGND 0.217f
C12 VPWR B 0.147f
C13 B X 6.52e-19
C14 a_29_53# B 0.121f
C15 C VPWR 0.00457f
C16 C a_29_53# 0.0857f
C17 a_183_297# VPWR 8.13e-19
C18 VPWR X 0.0885f
C19 a_111_297# VPWR 5.94e-19
C20 a_29_53# VPWR 0.0833f
C21 VGND A 0.0187f
C22 a_29_53# a_183_297# 0.00868f
C23 a_29_53# X 0.0991f
C24 a_29_53# a_111_297# 0.005f
C25 B A 0.0787f
C26 C A 0.0343f
C27 VGND VPB 0.00724f
C28 VPWR A 0.00936f
C29 a_183_297# A 0.00239f
C30 VPB B 0.0962f
C31 A X 0.00127f
C32 a_111_297# A 0.00223f
C33 a_29_53# A 0.242f
C34 C VPB 0.0396f
C35 VGND VNB 0.306f
C36 X VNB 0.0882f
C37 A VNB 0.117f
C38 C VNB 0.16f
C39 B VNB 0.117f
C40 VPWR VNB 0.253f
C41 VPB VNB 0.516f
C42 a_29_53# VNB 0.18f
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
C0 VPWR VGND 0.903f
C1 VPB VGND 0.161f
C2 VPWR VPB 0.0858f
C3 VPWR VNB 0.867f
C4 VGND VNB 0.761f
C5 VPB VNB 0.605f
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 B VGND 0.0451f
C1 a_109_297# Y 0.0113f
C2 VGND Y 0.154f
C3 VPWR VPB 0.0449f
C4 B VPWR 0.0148f
C5 VGND A 0.0486f
C6 B VPB 0.0367f
C7 VPWR Y 0.0995f
C8 VPB Y 0.0139f
C9 a_109_297# VGND 0.00128f
C10 B Y 0.0877f
C11 VPWR A 0.0528f
C12 VPB A 0.0415f
C13 B A 0.0584f
C14 VPWR a_109_297# 0.00638f
C15 VPWR VGND 0.0314f
C16 A Y 0.0471f
C17 VPB VGND 0.00456f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X a_193_297# a_465_47#
+ a_205_47# a_109_297# a_27_47#
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
C0 X VGND 0.061f
C1 C1 a_27_47# 0.0792f
C2 A2 VPB 0.027f
C3 B1 VPB 0.0321f
C4 VGND a_109_297# 0.00284f
C5 a_193_297# VPB 0.00774f
C6 B2 C1 0.0726f
C7 VGND B1 0.0133f
C8 X VPWR 0.0897f
C9 VGND A2 0.0168f
C10 a_27_47# VPB 0.0512f
C11 a_193_297# VGND 0.00438f
C12 VPWR a_109_297# 0.15f
C13 B2 VPB 0.0256f
C14 VGND a_27_47# 0.395f
C15 A1 C1 1.77e-20
C16 VGND a_465_47# 0.00257f
C17 A2 VPWR 0.0209f
C18 VPWR B1 0.00982f
C19 a_193_297# VPWR 0.169f
C20 VGND B2 0.0174f
C21 VPWR a_27_47# 0.099f
C22 A1 VPB 0.0343f
C23 X a_109_297# 3.99e-19
C24 VPWR a_465_47# 5.05e-19
C25 VPWR B2 0.00842f
C26 VGND A1 0.0126f
C27 X A2 0.00157f
C28 X B1 9.58e-20
C29 a_193_297# X 0.00367f
C30 B1 a_109_297# 0.00736f
C31 X a_27_47# 0.0921f
C32 a_193_297# a_109_297# 0.0927f
C33 X a_465_47# 1.56e-19
C34 VGND a_205_47# 0.00156f
C35 A1 VPWR 0.0161f
C36 a_27_47# a_109_297# 0.0961f
C37 a_193_297# A2 0.00683f
C38 a_193_297# B1 0.00869f
C39 X B2 6.77e-20
C40 B2 a_109_297# 0.0133f
C41 A2 a_27_47# 0.153f
C42 B1 a_27_47# 0.112f
C43 a_193_297# a_27_47# 0.144f
C44 C1 VPB 0.0367f
C45 VPWR a_205_47# 1.62e-19
C46 B2 B1 0.0784f
C47 X A1 2.77e-19
C48 a_193_297# B2 0.00126f
C49 VGND C1 0.0196f
C50 a_27_47# a_465_47# 0.013f
C51 A1 a_109_297# 1.05e-19
C52 B2 a_27_47# 0.0959f
C53 VGND VPB 0.00844f
C54 A1 B1 0.0609f
C55 A1 A2 0.0692f
C56 a_193_297# A1 0.0109f
C57 VPWR C1 0.0139f
C58 A1 a_27_47# 0.0984f
C59 VPWR VPB 0.0799f
C60 A1 a_465_47# 7.06e-19
C61 X C1 5.03e-20
C62 VGND VPWR 0.0722f
C63 a_27_47# a_205_47# 0.00762f
C64 C1 a_109_297# 0.00739f
C65 X VPB 0.0113f
C66 A2 C1 9.03e-21
C67 B1 C1 6.46e-19
C68 a_109_297# VPB 0.00421f
C69 VGND VNB 0.437f
C70 X VNB 0.0919f
C71 VPWR VNB 0.364f
C72 A2 VNB 0.0896f
C73 A1 VNB 0.106f
C74 B1 VNB 0.108f
C75 B2 VNB 0.0887f
C76 C1 VNB 0.139f
C77 VPB VNB 0.782f
C78 a_193_297# VNB 0.0011f
C79 a_109_297# VNB 7.11e-19
C80 a_27_47# VNB 0.216f
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X a_256_47# a_584_47#
+ a_93_21# a_250_297# a_346_47#
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
C0 A3 VPB 0.0291f
C1 A3 A2 0.0788f
C2 a_250_297# B2 0.0344f
C3 a_93_21# VGND 0.251f
C4 a_256_47# VGND 0.00394f
C5 B1 VGND 0.0344f
C6 A3 X 2.45e-19
C7 a_346_47# VPWR 0.00109f
C8 VGND VPB 0.00788f
C9 A2 VGND 0.0114f
C10 VGND X 0.06f
C11 a_346_47# A1 0.00465f
C12 a_250_297# A3 0.00602f
C13 a_584_47# VPWR 9.47e-19
C14 a_346_47# a_93_21# 0.0119f
C15 B1 a_346_47# 5.39e-20
C16 VPWR A1 0.016f
C17 a_346_47# A2 0.00252f
C18 a_250_297# VGND 0.0072f
C19 A3 B2 9.12e-20
C20 a_93_21# VPWR 0.0907f
C21 a_256_47# VPWR 9.47e-19
C22 B1 VPWR 0.01f
C23 a_584_47# a_93_21# 0.00278f
C24 VPWR VPB 0.0756f
C25 B1 a_584_47# 0.00143f
C26 VPWR A2 0.0133f
C27 VGND B2 0.0469f
C28 a_93_21# A1 0.0641f
C29 B1 A1 0.0965f
C30 VPWR X 0.0849f
C31 A1 VPB 0.0296f
C32 a_256_47# a_93_21# 0.0114f
C33 A2 A1 0.0971f
C34 B1 a_93_21# 0.0774f
C35 B1 a_256_47# 2.07e-20
C36 a_93_21# VPB 0.0485f
C37 B1 VPB 0.0276f
C38 A1 X 6.03e-20
C39 a_93_21# A2 0.0747f
C40 a_256_47# A2 0.00256f
C41 B1 A2 1.44e-20
C42 A3 VGND 0.00974f
C43 a_250_297# VPWR 0.313f
C44 A2 VPB 0.0287f
C45 a_93_21# X 0.0841f
C46 B1 X 3.83e-20
C47 a_584_47# a_250_297# 2.43e-19
C48 X VPB 0.0108f
C49 A2 X 1.19e-19
C50 a_250_297# A1 0.0129f
C51 VPWR B2 0.0108f
C52 a_250_297# a_93_21# 0.188f
C53 B1 a_250_297# 0.0125f
C54 a_250_297# VPB 0.00616f
C55 A1 B2 3.14e-19
C56 a_250_297# A2 0.0129f
C57 a_93_21# B2 0.0147f
C58 a_250_297# X 5.42e-19
C59 a_346_47# VGND 0.00514f
C60 B1 B2 0.0823f
C61 VPWR A3 0.0158f
C62 B2 VPB 0.0355f
C63 A2 B2 1.46e-19
C64 VPWR VGND 0.076f
C65 a_584_47# VGND 0.00683f
C66 a_93_21# A3 0.124f
C67 a_256_47# A3 4.42e-19
C68 B1 A3 7.88e-22
C69 A1 VGND 0.0133f
C70 VGND VNB 0.465f
C71 VPWR VNB 0.365f
C72 X VNB 0.0937f
C73 B2 VNB 0.14f
C74 B1 VNB 0.101f
C75 A1 VNB 0.0951f
C76 A2 VNB 0.0921f
C77 A3 VNB 0.0929f
C78 VPB VNB 0.782f
C79 a_250_297# VNB 0.0278f
C80 a_93_21# VNB 0.151f
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X a_277_297# a_205_297# a_27_297#
+ a_109_297#
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 B VGND 0.0159f
C1 B a_27_297# 0.159f
C2 C VPWR 0.00723f
C3 a_205_297# VPWR 5.16e-19
C4 A VPB 0.033f
C5 VPWR VGND 0.0546f
C6 X A 0.00133f
C7 a_27_297# VPWR 0.084f
C8 D B 0.00287f
C9 X VPB 0.0109f
C10 C A 0.028f
C11 A VGND 0.016f
C12 A a_27_297# 0.163f
C13 D VPWR 0.00503f
C14 B a_277_297# 2.29e-19
C15 C VPB 0.0338f
C16 VPB VGND 0.00796f
C17 X VGND 0.0354f
C18 VPB a_27_297# 0.0517f
C19 VPWR a_277_297# 7.48e-19
C20 C a_109_297# 0.00356f
C21 X a_27_297# 0.0991f
C22 a_109_297# VGND 7.58e-19
C23 D A 2.13e-19
C24 a_27_297# a_109_297# 0.00695f
C25 a_205_297# C 0.00261f
C26 C VGND 0.0191f
C27 a_205_297# VGND 3.36e-19
C28 C a_27_297# 0.158f
C29 a_205_297# a_27_297# 0.00412f
C30 B VPWR 0.193f
C31 D VPB 0.0405f
C32 a_27_297# VGND 0.235f
C33 A a_277_297# 2.28e-19
C34 X a_277_297# 6.43e-20
C35 D C 0.0954f
C36 A B 0.0639f
C37 D VGND 0.0517f
C38 D a_27_297# 0.054f
C39 C a_277_297# 5.54e-19
C40 A VPWR 0.00769f
C41 VPB B 0.106f
C42 a_277_297# VGND 4.65e-19
C43 X B 6.42e-19
C44 a_27_297# a_277_297# 0.00876f
C45 VPB VPWR 0.075f
C46 X VPWR 0.0878f
C47 C B 0.0917f
C48 a_109_297# VPWR 9.23e-19
C49 VGND VNB 0.367f
C50 X VNB 0.0883f
C51 A VNB 0.109f
C52 C VNB 0.105f
C53 D VNB 0.175f
C54 B VNB 0.115f
C55 VPWR VNB 0.29f
C56 VPB VNB 0.605f
C57 a_27_297# VNB 0.163f
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
C0 VGND VPB 0.35f
C1 VGND VPWR 1.57f
C2 VPWR VPB 0.137f
C3 VPWR VNB 1.67f
C4 VGND VNB 1.47f
C5 VPB VNB 1.14f
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X a_369_47# a_469_47#
+ a_297_47# a_193_413# a_27_47#
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_193_413# VPB 0.0644f
C1 a_193_413# B 0.144f
C2 a_297_47# VPWR 2.82e-19
C3 a_193_413# X 0.108f
C4 VGND A_N 0.0205f
C5 a_27_47# VPB 0.092f
C6 B a_27_47# 0.0794f
C7 a_469_47# C 0.00202f
C8 VGND C 0.0395f
C9 a_297_47# a_193_413# 0.00137f
C10 VGND a_369_47# 0.00505f
C11 D a_469_47# 0.00183f
C12 D VGND 0.0372f
C13 VGND VPB 0.0123f
C14 VGND B 0.037f
C15 a_193_413# VPWR 0.281f
C16 a_469_47# X 0.001f
C17 VGND X 0.0588f
C18 A_N VPB 0.0832f
C19 a_27_47# VPWR 0.106f
C20 a_369_47# C 0.00448f
C21 D C 0.183f
C22 C VPB 0.0742f
C23 VGND a_297_47# 0.00183f
C24 B C 0.164f
C25 D VPB 0.0763f
C26 C X 0.00479f
C27 a_369_47# B 0.00129f
C28 a_193_413# a_27_47# 0.125f
C29 B VPB 0.089f
C30 a_469_47# VPWR 7.77e-19
C31 VGND VPWR 0.0727f
C32 D X 0.0168f
C33 X VPB 0.0108f
C34 A_N VPWR 0.02f
C35 a_469_47# a_193_413# 0.00109f
C36 VGND a_193_413# 0.0915f
C37 C VPWR 0.0182f
C38 a_297_47# B 0.00353f
C39 a_369_47# VPWR 6.65e-19
C40 VGND a_27_47# 0.103f
C41 D VPWR 0.0186f
C42 A_N a_193_413# 0.00151f
C43 VPWR VPB 0.0818f
C44 B VPWR 0.0186f
C45 a_193_413# C 0.0389f
C46 A_N a_27_47# 0.237f
C47 VPWR X 0.0586f
C48 a_369_47# a_193_413# 0.00181f
C49 VGND a_469_47# 0.00551f
C50 D a_193_413# 0.155f
C51 VGND VNB 0.456f
C52 X VNB 0.0934f
C53 VPWR VNB 0.368f
C54 D VNB 0.123f
C55 C VNB 0.108f
C56 B VNB 0.12f
C57 A_N VNB 0.198f
C58 VPB VNB 0.782f
C59 a_193_413# VNB 0.136f
C60 a_27_47# VNB 0.224f
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X a_109_93# a_368_53# a_209_311#
+ a_296_53#
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
C0 C VPWR 0.005f
C1 C a_209_311# 0.19f
C2 VGND B 0.00796f
C3 C VPB 0.0339f
C4 B VPWR 0.131f
C5 A_N a_109_93# 0.117f
C6 a_209_311# B 0.0609f
C7 B VPB 0.0914f
C8 X C 0.0176f
C9 A_N VGND 0.045f
C10 A_N VPWR 0.0513f
C11 a_109_93# a_296_53# 1.84e-19
C12 X B 0.00119f
C13 A_N a_209_311# 0.00515f
C14 VGND a_109_93# 0.0784f
C15 A_N VPB 0.111f
C16 a_109_93# VPWR 0.0984f
C17 a_109_93# a_209_311# 0.168f
C18 VGND a_296_53# 6.07e-19
C19 a_109_93# VPB 0.0652f
C20 a_296_53# VPWR 1.15e-19
C21 A_N X 1.44e-19
C22 a_209_311# a_296_53# 0.0049f
C23 a_368_53# VGND 0.0031f
C24 VGND VPWR 0.0657f
C25 a_368_53# VPWR 4.26e-19
C26 VGND a_209_311# 0.131f
C27 a_368_53# a_209_311# 0.0026f
C28 C B 0.0671f
C29 a_209_311# VPWR 0.155f
C30 VGND VPB 0.00909f
C31 VPB VPWR 0.104f
C32 a_209_311# VPB 0.0515f
C33 X VGND 0.0647f
C34 A_N C 7.6e-19
C35 X VPWR 0.0732f
C36 X a_209_311# 0.0877f
C37 X VPB 0.0119f
C38 A_N B 2.03e-19
C39 a_109_93# C 3.91e-20
C40 a_109_93# B 0.0802f
C41 VGND C 0.0678f
C42 a_368_53# C 0.00415f
C43 VGND VNB 0.44f
C44 X VNB 0.0925f
C45 C VNB 0.114f
C46 B VNB 0.101f
C47 VPWR VNB 0.342f
C48 A_N VNB 0.197f
C49 VPB VNB 0.693f
C50 a_209_311# VNB 0.143f
C51 a_109_93# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
C0 VPB a_27_47# 0.139f
C1 VGND X 0.216f
C2 A VPB 0.0321f
C3 VPWR X 0.317f
C4 X a_27_47# 0.328f
C5 VGND VPWR 0.057f
C6 VGND a_27_47# 0.148f
C7 A X 0.014f
C8 VPWR a_27_47# 0.219f
C9 VGND A 0.0431f
C10 A VPWR 0.022f
C11 X VPB 0.0122f
C12 A a_27_47# 0.195f
C13 VGND VPB 0.00583f
C14 VPWR VPB 0.0632f
C15 VGND VNB 0.358f
C16 X VNB 0.067f
C17 VPWR VNB 0.308f
C18 A VNB 0.148f
C19 VPB VNB 0.605f
C20 a_27_47# VNB 0.543f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
C0 VPWR a_145_75# 6.31e-19
C1 A VGND 0.0147f
C2 a_145_75# a_59_75# 0.00658f
C3 X VGND 0.0993f
C4 B A 0.0971f
C5 B X 0.00276f
C6 B VGND 0.0115f
C7 VPWR A 0.0362f
C8 X VPWR 0.111f
C9 A a_59_75# 0.0809f
C10 X a_59_75# 0.109f
C11 VPWR VGND 0.0461f
C12 B VPWR 0.0117f
C13 VGND a_59_75# 0.116f
C14 B a_59_75# 0.143f
C15 VPB A 0.0806f
C16 X VPB 0.0127f
C17 VPWR a_59_75# 0.15f
C18 VPB VGND 0.008f
C19 B VPB 0.0629f
C20 VPB VPWR 0.0729f
C21 VPB a_59_75# 0.0563f
C22 X a_145_75# 5.76e-19
C23 VGND a_145_75# 0.00468f
C24 X A 1.68e-19
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y a_297_297# a_191_297#
+ a_109_297#
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPWR A 0.0483f
C1 VPWR a_297_297# 0.00317f
C2 VGND D 0.0456f
C3 VPB Y 0.0127f
C4 VPWR C 0.0509f
C5 Y A 0.0175f
C6 a_297_297# Y 1.24e-19
C7 Y C 0.125f
C8 VGND VPWR 0.0492f
C9 B a_191_297# 0.00223f
C10 VGND Y 0.151f
C11 VPWR D 0.0128f
C12 a_109_297# C 0.0062f
C13 VPB B 0.0304f
C14 B A 0.11f
C15 Y D 0.108f
C16 B a_297_297# 0.0132f
C17 a_191_297# C 0.0195f
C18 B C 0.173f
C19 a_109_297# VGND 0.00181f
C20 VPB A 0.041f
C21 VPWR Y 0.0561f
C22 VGND a_191_297# 9.29e-19
C23 a_297_297# A 3.16e-19
C24 VPB C 0.0299f
C25 B VGND 0.0191f
C26 C A 0.00268f
C27 VPB VGND 0.0048f
C28 a_109_297# VPWR 0.00576f
C29 VGND A 0.0526f
C30 VGND a_297_297# 8.1e-19
C31 VGND C 0.0184f
C32 a_109_297# Y 0.0122f
C33 VPB D 0.0376f
C34 a_191_297# VPWR 0.0049f
C35 B VPWR 0.0887f
C36 a_191_297# Y 0.00142f
C37 D C 0.0523f
C38 B Y 0.0403f
C39 VPB VPWR 0.0524f
C40 VGND VNB 0.322f
C41 VPWR VNB 0.276f
C42 Y VNB 0.0645f
C43 A VNB 0.174f
C44 B VNB 0.0968f
C45 C VNB 0.0911f
C46 D VNB 0.159f
C47 VPB VNB 0.516f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X a_75_212#
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 VPWR VPB 0.0355f
C1 a_75_212# VGND 0.105f
C2 X A 8.48e-19
C3 VPWR VGND 0.0289f
C4 X VPB 0.0128f
C5 a_75_212# VPWR 0.134f
C6 X VGND 0.0545f
C7 A VPB 0.0525f
C8 a_75_212# X 0.107f
C9 X VPWR 0.0896f
C10 VGND A 0.0184f
C11 VGND VPB 0.00507f
C12 a_75_212# A 0.178f
C13 a_75_212# VPB 0.0571f
C14 VPWR A 0.0217f
C15 VGND VNB 0.207f
C16 VPWR VNB 0.176f
C17 X VNB 0.0942f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_75_212# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 X VPB 0.0128f
C1 a_27_47# VGND 0.105f
C2 VPWR A 0.0215f
C3 X VGND 0.0546f
C4 VPWR VPB 0.0355f
C5 a_27_47# X 0.107f
C6 VPWR VGND 0.029f
C7 A VPB 0.0524f
C8 a_27_47# VPWR 0.135f
C9 VPWR X 0.0897f
C10 VGND A 0.0184f
C11 VGND VPB 0.00505f
C12 a_27_47# A 0.181f
C13 a_27_47# VPB 0.0592f
C14 X A 8.48e-19
C15 VGND VNB 0.207f
C16 X VNB 0.0941f
C17 VPWR VNB 0.175f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_27_47# VNB 0.208f
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X a_664_47# a_841_47#
+ a_381_47# a_62_47# a_558_47#
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_664_47# VGND 0.125f
C1 VPB VPWR 0.103f
C2 X VPWR 0.108f
C3 a_558_47# a_381_47# 0.16f
C4 a_62_47# VPB 0.0515f
C5 a_62_47# X 0.156f
C6 VGND a_558_47# 0.0816f
C7 a_841_47# a_664_47# 0.134f
C8 a_62_47# VPWR 0.149f
C9 VPB a_381_47# 0.0447f
C10 X a_381_47# 0.318f
C11 VPB VGND 0.008f
C12 a_841_47# a_558_47# 0.00368f
C13 X VGND 0.106f
C14 VPB A 0.105f
C15 X A 0.0142f
C16 VPWR a_381_47# 0.134f
C17 VPWR VGND 0.0902f
C18 a_62_47# VGND 0.144f
C19 VPWR A 0.0174f
C20 a_62_47# A 0.244f
C21 a_841_47# VPB 0.0108f
C22 a_664_47# a_558_47# 0.314f
C23 a_841_47# VPWR 0.0614f
C24 VGND a_381_47# 0.125f
C25 A a_381_47# 5.42e-19
C26 VGND A 0.0176f
C27 VPB a_664_47# 0.043f
C28 X a_664_47# 6.67e-19
C29 a_841_47# VGND 0.0585f
C30 VPB a_558_47# 0.115f
C31 X a_558_47# 0.0144f
C32 VPWR a_664_47# 0.131f
C33 VPWR a_558_47# 0.084f
C34 X VPB 0.126f
C35 VGND VNB 0.537f
C36 VPWR VNB 0.439f
C37 X VNB 0.163f
C38 A VNB 0.198f
C39 VPB VNB 0.959f
C40 a_841_47# VNB 0.0929f
C41 a_664_47# VNB 0.13f
C42 a_558_47# VNB 0.164f
C43 a_381_47# VNB 0.11f
C44 a_62_47# VNB 0.169f
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y a_129_47# a_47_47# a_285_47#
+ a_377_297#
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VPB VGND 0.00568f
C1 VGND Y 0.0381f
C2 VPWR A 0.0349f
C3 VPWR a_377_297# 0.00559f
C4 a_285_47# VGND 0.211f
C5 VGND a_47_47# 0.104f
C6 VPWR a_129_47# 9.47e-19
C7 VPB A 0.0822f
C8 A Y 0.00181f
C9 a_377_297# Y 0.00188f
C10 A a_285_47# 0.0353f
C11 A a_47_47# 0.0307f
C12 a_377_297# a_47_47# 0.00899f
C13 VPB VPWR 0.0718f
C14 VPWR Y 0.107f
C15 VGND B 0.0389f
C16 VPWR a_285_47# 0.00255f
C17 a_129_47# a_47_47# 0.00369f
C18 VPWR a_47_47# 0.273f
C19 VPB Y 0.00878f
C20 VPB a_285_47# 5.53e-19
C21 a_285_47# Y 0.0439f
C22 A B 0.236f
C23 a_377_297# B 0.00254f
C24 VPB a_47_47# 0.0444f
C25 a_47_47# Y 0.143f
C26 a_285_47# a_47_47# 0.0175f
C27 a_129_47# B 0.00236f
C28 VPWR B 0.0408f
C29 A VGND 0.0635f
C30 a_377_297# VGND 0.00125f
C31 VPB B 0.0643f
C32 B Y 0.00334f
C33 a_285_47# B 0.067f
C34 a_129_47# VGND 0.00547f
C35 B a_47_47# 0.356f
C36 VPWR VGND 0.0665f
C37 VGND VNB 0.4f
C38 Y VNB 0.0783f
C39 VPWR VNB 0.352f
C40 A VNB 0.217f
C41 B VNB 0.212f
C42 VPB VNB 0.693f
C43 a_285_47# VNB 0.0174f
C44 a_47_47# VNB 0.199f
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X a_472_297# a_80_21#
+ a_300_47# a_217_297#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
C0 VPB A1 0.0266f
C1 a_80_21# X 0.118f
C2 C1 X 7.15e-20
C3 a_217_297# a_80_21# 0.127f
C4 a_217_297# C1 0.00262f
C5 VPWR a_300_47# 8.53e-19
C6 a_80_21# VGND 0.293f
C7 C1 VGND 0.0176f
C8 a_217_297# X 0.00271f
C9 A2 a_80_21# 0.128f
C10 a_80_21# a_472_297# 0.0164f
C11 X VGND 0.0654f
C12 a_80_21# VPWR 0.119f
C13 a_217_297# VGND 0.00342f
C14 C1 VPWR 0.0137f
C15 A2 X 6.82e-19
C16 a_80_21# B1 0.0964f
C17 C1 B1 0.0846f
C18 a_217_297# A2 0.0135f
C19 X a_472_297# 2.6e-19
C20 a_217_297# a_472_297# 0.00517f
C21 X VPWR 0.0884f
C22 a_300_47# A1 5.95e-19
C23 A2 VGND 0.0191f
C24 a_217_297# VPWR 0.197f
C25 X B1 1.18e-19
C26 VGND a_472_297# 0.00188f
C27 a_217_297# B1 0.00651f
C28 VPB a_80_21# 0.0661f
C29 C1 VPB 0.0379f
C30 VPWR VGND 0.0665f
C31 VGND B1 0.0175f
C32 A2 VPWR 0.0161f
C33 VPB X 0.0118f
C34 VPWR a_472_297# 0.00703f
C35 a_80_21# A1 0.111f
C36 a_217_297# VPB 0.00494f
C37 B1 a_472_297# 1.87e-19
C38 VPWR B1 0.0129f
C39 VPB VGND 0.00775f
C40 X A1 3.62e-19
C41 a_217_297# A1 0.0124f
C42 VPB A2 0.0384f
C43 VGND A1 0.0147f
C44 VPB VPWR 0.0754f
C45 A2 A1 0.0881f
C46 VPB B1 0.0267f
C47 a_80_21# a_300_47# 0.00997f
C48 VPWR A1 0.0149f
C49 X a_300_47# 5.31e-19
C50 A1 B1 0.0834f
C51 C1 a_80_21# 0.079f
C52 VGND a_300_47# 0.00536f
C53 VGND VNB 0.385f
C54 VPWR VNB 0.325f
C55 X VNB 0.0899f
C56 C1 VNB 0.144f
C57 B1 VNB 0.0899f
C58 A1 VNB 0.0905f
C59 A2 VNB 0.108f
C60 VPB VNB 0.693f
C61 a_217_297# VNB 0.00117f
C62 a_80_21# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VGND VPWR 0.0662f
C1 VGND a_109_47# 0.00223f
C2 C a_303_47# 0.00527f
C3 X VPWR 0.0945f
C4 D C 0.18f
C5 C VPB 0.0609f
C6 D a_303_47# 0.00119f
C7 B C 0.161f
C8 a_197_47# B 0.00623f
C9 C VPWR 0.021f
C10 a_197_47# VPWR 5.24e-19
C11 D VPB 0.0782f
C12 VGND a_27_47# 0.132f
C13 C a_109_47# 1.72e-20
C14 a_303_47# VPWR 4.83e-19
C15 D VPWR 0.0207f
C16 X a_27_47# 0.0754f
C17 B VPB 0.0643f
C18 A VPB 0.0907f
C19 VPB VPWR 0.077f
C20 A B 0.0839f
C21 B VPWR 0.0231f
C22 A VPWR 0.044f
C23 VGND X 0.0903f
C24 B a_109_47# 0.00153f
C25 C a_27_47# 0.0516f
C26 a_197_47# a_27_47# 0.00167f
C27 a_109_47# VPWR 4.66e-19
C28 a_303_47# a_27_47# 0.00119f
C29 D a_27_47# 0.107f
C30 C VGND 0.0408f
C31 a_197_47# VGND 0.00387f
C32 VPB a_27_47# 0.082f
C33 B a_27_47# 0.13f
C34 A a_27_47# 0.153f
C35 a_303_47# VGND 0.00381f
C36 a_27_47# VPWR 0.326f
C37 D VGND 0.0898f
C38 VGND VPB 0.00852f
C39 a_27_47# a_109_47# 0.00578f
C40 D X 0.00746f
C41 B VGND 0.0453f
C42 a_197_47# C 0.00123f
C43 A VGND 0.0151f
C44 VPB X 0.0111f
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X a_489_413# a_226_47#
+ a_556_47# a_226_297# a_76_199#
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPB B1 0.0803f
C1 a_76_199# a_556_47# 0.0017f
C2 B2 a_556_47# 0.00291f
C3 a_226_47# A1_N 0.0209f
C4 VPWR A1_N 0.00672f
C5 a_489_413# a_226_47# 0.00579f
C6 a_489_413# VPWR 0.143f
C7 a_226_47# VGND 0.149f
C8 VPWR VGND 0.0743f
C9 a_76_199# a_226_47# 0.188f
C10 VPWR a_76_199# 0.2f
C11 B2 a_226_47# 0.0975f
C12 B2 VPWR 0.0161f
C13 a_226_47# a_226_297# 0.00128f
C14 VPWR a_226_297# 8.54e-19
C15 A1_N VGND 0.0261f
C16 a_226_47# A2_N 0.141f
C17 VPWR A2_N 0.00449f
C18 a_489_413# VGND 0.0058f
C19 a_76_199# A1_N 0.119f
C20 a_226_47# X 0.0108f
C21 VPWR X 0.0589f
C22 a_489_413# a_76_199# 0.0473f
C23 A1_N a_226_297# 0.00184f
C24 B2 a_489_413# 0.0541f
C25 A1_N A2_N 0.11f
C26 a_76_199# VGND 0.108f
C27 B2 VGND 0.0335f
C28 A1_N X 0.00211f
C29 VGND a_226_297# 5.63e-19
C30 VPB a_226_47# 0.111f
C31 VPWR VPB 0.0951f
C32 A2_N VGND 0.0174f
C33 B2 a_76_199# 0.0626f
C34 a_76_199# a_226_297# 0.00354f
C35 VGND X 0.0627f
C36 a_76_199# A2_N 0.0125f
C37 VPB A1_N 0.0339f
C38 a_76_199# X 0.0995f
C39 VPWR B1 0.0188f
C40 a_489_413# VPB 0.015f
C41 A2_N X 2.55e-19
C42 VPB VGND 0.0128f
C43 a_489_413# B1 0.0382f
C44 VPB a_76_199# 0.0817f
C45 B2 VPB 0.0645f
C46 VGND B1 0.0471f
C47 VPB A2_N 0.0327f
C48 a_76_199# B1 0.00185f
C49 VPB X 0.0113f
C50 VPWR a_556_47# 7.24e-19
C51 B2 B1 0.182f
C52 VPWR a_226_47# 0.0187f
C53 VGND a_556_47# 0.00639f
C54 VGND VNB 0.462f
C55 A2_N VNB 0.103f
C56 A1_N VNB 0.111f
C57 VPWR VNB 0.369f
C58 X VNB 0.0975f
C59 B1 VNB 0.206f
C60 B2 VNB 0.106f
C61 VPB VNB 0.782f
C62 a_489_413# VNB 0.0254f
C63 a_226_47# VNB 0.162f
C64 a_76_199# VNB 0.141f
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X a_515_93# a_223_47#
+ a_615_93# a_343_93# a_429_93# a_27_47#
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
C0 X D 0.0193f
C1 VGND a_343_93# 0.0548f
C2 VPB a_223_47# 0.0799f
C3 A_N VPWR 0.0318f
C4 a_27_47# VPWR 0.0897f
C5 X a_343_93# 0.126f
C6 VPWR D 0.0143f
C7 C B_N 9.56e-20
C8 a_615_93# VPWR 8.49e-19
C9 VPB VGND 0.0167f
C10 VPWR a_343_93# 0.255f
C11 VPB X 0.0103f
C12 C a_515_93# 0.00389f
C13 A_N B_N 0.117f
C14 a_27_47# B_N 0.138f
C15 VGND a_223_47# 0.199f
C16 B_N D 6.67e-20
C17 VPB VPWR 0.106f
C18 B_N a_343_93# 0.00112f
C19 a_429_93# a_343_93# 0.00484f
C20 C D 0.163f
C21 VPWR a_223_47# 0.114f
C22 X VGND 0.0609f
C23 C a_615_93# 0.00407f
C24 a_515_93# a_343_93# 0.00115f
C25 C a_343_93# 0.0397f
C26 VPB B_N 0.0646f
C27 a_27_47# A_N 0.0906f
C28 VGND VPWR 0.0906f
C29 X VPWR 0.0582f
C30 a_615_93# D 0.00564f
C31 B_N a_223_47# 0.0431f
C32 a_429_93# a_223_47# 0.00492f
C33 a_27_47# a_343_93# 0.0406f
C34 C VPB 0.0686f
C35 a_343_93# D 0.114f
C36 a_615_93# a_343_93# 0.00103f
C37 B_N VGND 0.0427f
C38 a_429_93# VGND 0.00122f
C39 a_515_93# a_223_47# 0.00482f
C40 C a_223_47# 0.151f
C41 VPB A_N 0.0848f
C42 a_27_47# VPB 0.154f
C43 B_N X 4.64e-20
C44 VPB D 0.081f
C45 a_515_93# VGND 0.00408f
C46 C VGND 0.025f
C47 B_N VPWR 0.0168f
C48 VPB a_343_93# 0.0857f
C49 A_N a_223_47# 0.00833f
C50 a_429_93# VPWR 5.19e-19
C51 a_27_47# a_223_47# 0.267f
C52 a_223_47# D 4.03e-19
C53 A_N VGND 0.0146f
C54 a_515_93# VPWR 7.86e-19
C55 a_27_47# VGND 0.0715f
C56 a_223_47# a_343_93# 0.269f
C57 VGND D 0.0414f
C58 C VPWR 0.012f
C59 VGND a_615_93# 0.0044f
C60 VGND VNB 0.553f
C61 X VNB 0.0908f
C62 VPWR VNB 0.453f
C63 D VNB 0.124f
C64 C VNB 0.107f
C65 B_N VNB 0.134f
C66 A_N VNB 0.144f
C67 VPB VNB 0.959f
C68 a_343_93# VNB 0.172f
C69 a_223_47# VNB 0.141f
C70 a_27_47# VNB 0.259f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 B VGND 0.0304f
C1 A X 0.00166f
C2 VPB VGND 0.00696f
C3 A B 0.221f
C4 A VPB 0.051f
C5 a_35_297# a_117_297# 0.00641f
C6 VPWR a_117_297# 0.00852f
C7 B X 0.0149f
C8 VPB X 0.0154f
C9 a_117_297# VGND 0.00177f
C10 a_285_297# a_35_297# 0.025f
C11 VPWR a_285_297# 0.246f
C12 VPB B 0.0697f
C13 a_285_297# VGND 0.00394f
C14 VPWR a_35_297# 0.096f
C15 a_35_297# a_285_47# 0.00723f
C16 VPWR a_285_47# 8.6e-19
C17 a_35_297# VGND 0.177f
C18 a_117_297# X 2.25e-19
C19 VPWR VGND 0.0643f
C20 a_285_297# A 0.00749f
C21 VGND a_285_47# 0.00552f
C22 a_117_297# B 0.00777f
C23 a_285_297# X 0.0712f
C24 A a_35_297# 0.0633f
C25 VPWR A 0.0348f
C26 a_285_297# B 0.0553f
C27 A VGND 0.0325f
C28 a_35_297# X 0.166f
C29 VPWR X 0.0537f
C30 X a_285_47# 0.00206f
C31 a_285_297# VPB 0.0133f
C32 a_35_297# B 0.203f
C33 VPWR B 0.0703f
C34 X VGND 0.173f
C35 B a_285_47# 3.98e-19
C36 a_35_297# VPB 0.0699f
C37 VPWR VPB 0.0689f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X a_465_297# a_297_297#
+ a_215_297# a_392_297# a_109_53#
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 VGND A 0.0158f
C1 VPWR a_109_53# 0.0418f
C2 B X 6.65e-19
C3 a_215_297# X 0.0991f
C4 VGND a_297_297# 6.5e-19
C5 X A 0.00127f
C6 C a_392_297# 0.00267f
C7 D_N VPB 0.0461f
C8 VPWR VGND 0.075f
C9 C a_465_297# 6.89e-19
C10 a_215_297# D_N 3.19e-19
C11 a_215_297# a_392_297# 0.00419f
C12 VPWR X 0.0885f
C13 C VPB 0.0337f
C14 VGND a_109_53# 0.118f
C15 a_215_297# a_465_297# 0.00827f
C16 C B 0.0893f
C17 a_465_297# A 5.42e-19
C18 a_215_297# C 0.161f
C19 C A 0.0281f
C20 B VPB 0.116f
C21 a_215_297# VPB 0.0508f
C22 VPB A 0.0325f
C23 C a_297_297# 0.00375f
C24 VPWR D_N 0.0412f
C25 a_392_297# VPWR 5.29e-19
C26 a_215_297# B 0.159f
C27 B A 0.0666f
C28 a_215_297# A 0.157f
C29 VGND X 0.0359f
C30 VPWR a_465_297# 7.08e-19
C31 D_N a_109_53# 0.0889f
C32 a_215_297# a_297_297# 0.00659f
C33 C VPWR 0.00753f
C34 VPWR VPB 0.122f
C35 C a_109_53# 0.0984f
C36 VPWR B 0.255f
C37 a_215_297# VPWR 0.0871f
C38 D_N VGND 0.0531f
C39 a_392_297# VGND 3.44e-19
C40 VPWR A 0.0073f
C41 VPB a_109_53# 0.0547f
C42 B a_109_53# 0.0246f
C43 VPWR a_297_297# 8.59e-19
C44 a_215_297# a_109_53# 0.0807f
C45 a_465_297# VGND 5.02e-19
C46 a_109_53# A 1.19e-19
C47 C VGND 0.0202f
C48 VGND VPB 0.0115f
C49 a_109_53# a_297_297# 7.06e-21
C50 B VGND 0.0161f
C51 a_215_297# VGND 0.237f
C52 VPB X 0.011f
C53 VGND VNB 0.469f
C54 X VNB 0.0884f
C55 A VNB 0.108f
C56 C VNB 0.101f
C57 D_N VNB 0.185f
C58 B VNB 0.101f
C59 VPWR VNB 0.399f
C60 VPB VNB 0.782f
C61 a_109_53# VNB 0.159f
C62 a_215_297# VNB 0.142f
.ends

.subckt therm_raw b[0] b[2] b[3] p[11] p[12] p[13] p[14] p[1] p[2] p[4] p[5] p[8]
+ p[9] input3/a_27_47# net7 input13/a_27_47# net3 net15 net14 input7/a_27_47# _04_
+ input9/a_75_212# b[1] _27_/a_27_297# input1/a_75_212# input5/a_62_47# net2 p[0]
+ input5/a_381_47# _19_ net8 input8/a_27_47# p[7] output17/a_27_47# _01_ _02_ input15/a_27_47#
+ input5/a_558_47# _15_ p[3] input5/a_664_47# _08_ input6/a_27_47# net17 net5 VPWR
+ p[10] VGND p[6]
X_49_ net7 _02_ _19_ _20_ _21_ VGND VGND VPWR VPWR net17 _49_/a_208_47# _49_/a_75_199#
+ _49_/a_544_297# _49_/a_315_47# _49_/a_201_297# sky130_fd_sc_hd__a311o_1
X_48_ net11 _02_ _07_ VGND VGND VPWR VPWR _21_ _48_/a_181_47# _48_/a_109_47# _48_/a_27_47#
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ net5 _12_ _17_ VGND VGND VPWR VPWR _20_ _47_/a_384_47# _47_/a_81_21# _47_/a_299_297#
+ sky130_fd_sc_hd__a21o_1
X_46_ _04_ VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__inv_2
X_29_ net11 net13 net12 VGND VGND VPWR VPWR _03_ _29_/a_29_53# _29_/a_183_297# _29_/a_111_297#
+ sky130_fd_sc_hd__or3_1
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28_ _00_ _01_ VGND VGND VPWR VPWR _02_ _28_/a_109_297# sky130_fd_sc_hd__nor2_1
X_45_ _02_ _09_ _12_ _13_ _18_ VGND VGND VPWR VPWR net16 _45_/a_193_297# _45_/a_465_47#
+ _45_/a_205_47# _45_/a_109_297# _45_/a_27_47# sky130_fd_sc_hd__a221o_1
X_44_ net14 _14_ _15_ _17_ net2 VGND VGND VPWR VPWR _18_ _44_/a_256_47# _44_/a_584_47#
+ _44_/a_93_21# _44_/a_250_297# _44_/a_346_47# sky130_fd_sc_hd__a32o_1
X_27_ net14 net15 net3 net2 VGND VGND VPWR VPWR _01_ _27_/a_277_297# _27_/a_205_297#
+ _27_/a_27_297# _27_/a_109_297# sky130_fd_sc_hd__or4_1
XFILLER_0_7_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_26_ net5 net4 net6 VGND VGND VPWR VPWR _00_ _26_/a_29_53# _26_/a_183_297# _26_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_43_ _00_ _06_ _10_ _16_ VGND VGND VPWR VPWR _17_ _43_/a_369_47# _43_/a_469_47# _43_/a_297_47#
+ _43_/a_193_413# _43_/a_27_47# sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_42_ net3 net15 net14 VGND VGND VPWR VPWR _16_ _42_/a_109_93# _42_/a_368_53# _42_/a_209_311#
+ _42_/a_296_53# sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_3_Left_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND VPWR VPWR b[0] output16/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_41_ _06_ _10_ VGND VGND VPWR VPWR _15_ _41_/a_145_75# _41_/a_59_75# sky130_fd_sc_hd__and2_1
Xoutput17 net17 VGND VGND VPWR VPWR b[1] output17/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_40_ net15 net3 net2 _00_ VGND VGND VPWR VPWR _14_ _40_/a_297_297# _40_/a_191_297#
+ _40_/a_109_297# sky130_fd_sc_hd__nor4_1
Xoutput18 net18 VGND VGND VPWR VPWR b[2] output18/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR b[3] output19/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_7_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 p[0] VGND VGND VPWR VPWR net1 input1/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput2 p[10] VGND VGND VPWR VPWR net2 input2/a_27_47# sky130_fd_sc_hd__buf_1
Xinput3 p[11] VGND VGND VPWR VPWR net3 input3/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 p[12] VGND VGND VPWR VPWR net4 input4/a_75_212# sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 p[13] VGND VGND VPWR VPWR net5 input5/a_664_47# input5/a_841_47# input5/a_381_47#
+ input5/a_62_47# input5/a_558_47# sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_1_Left_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 p[14] VGND VGND VPWR VPWR net6 input6/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 p[1] VGND VGND VPWR VPWR net7 input7/a_27_47# sky130_fd_sc_hd__buf_1
Xinput10 p[4] VGND VGND VPWR VPWR net10 input10/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 p[2] VGND VGND VPWR VPWR net8 input8/a_27_47# sky130_fd_sc_hd__buf_1
Xinput11 p[5] VGND VGND VPWR VPWR net11 input11/a_27_47# sky130_fd_sc_hd__buf_1
X_39_ net5 net6 VGND VGND VPWR VPWR _13_ _39_/a_129_47# _39_/a_47_47# _39_/a_285_47#
+ _39_/a_377_297# sky130_fd_sc_hd__xnor2_1
Xinput9 p[3] VGND VGND VPWR VPWR net9 input9/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput12 p[6] VGND VGND VPWR VPWR net12 input12/a_27_47# sky130_fd_sc_hd__buf_1
X_55_ _14_ _15_ _20_ _22_ VGND VGND VPWR VPWR net19 _55_/a_472_297# _55_/a_80_21#
+ _55_/a_300_47# _55_/a_217_297# sky130_fd_sc_hd__a211o_1
X_38_ net4 _06_ _10_ _11_ VGND VGND VPWR VPWR _12_ _38_/a_109_47# _38_/a_197_47# _38_/a_303_47#
+ _38_/a_27_47# sky130_fd_sc_hd__and4_1
X_54_ _25_ VGND VGND VPWR VPWR net18 _54_/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput13 p[7] VGND VGND VPWR VPWR net13 input13/a_27_47# sky130_fd_sc_hd__buf_1
X_37_ net14 net15 net3 net2 VGND VGND VPWR VPWR _11_ _37_/a_109_47# _37_/a_197_47#
+ _37_/a_303_47# _37_/a_27_47# sky130_fd_sc_hd__and4_1
X_53_ _21_ _22_ _24_ VGND VGND VPWR VPWR _25_ _53_/a_29_53# _53_/a_183_297# _53_/a_111_297#
+ sky130_fd_sc_hd__or3_1
Xinput14 p[8] VGND VGND VPWR VPWR net14 input14/a_27_47# sky130_fd_sc_hd__buf_1
X_36_ net11 net10 net13 net12 VGND VGND VPWR VPWR _10_ _36_/a_109_47# _36_/a_197_47#
+ _36_/a_303_47# _36_/a_27_47# sky130_fd_sc_hd__and4_1
X_52_ _02_ _06_ _23_ _12_ net5 VGND VGND VPWR VPWR _24_ _52_/a_256_47# _52_/a_584_47#
+ _52_/a_93_21# _52_/a_250_297# _52_/a_346_47# sky130_fd_sc_hd__a32o_1
X_35_ _04_ _05_ _07_ _08_ VGND VGND VPWR VPWR _09_ _35_/a_489_413# _35_/a_226_47#
+ _35_/a_556_47# _35_/a_226_297# _35_/a_76_199# sky130_fd_sc_hd__a2bb2o_1
Xinput15 p[9] VGND VGND VPWR VPWR net15 input15/a_27_47# sky130_fd_sc_hd__buf_1
X_51_ _03_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__inv_2
X_34_ net11 net12 VGND VGND VPWR VPWR _08_ _34_/a_129_47# _34_/a_47_47# _34_/a_285_47#
+ _34_/a_377_297# sky130_fd_sc_hd__xnor2_1
X_33_ net13 _06_ net10 VGND VGND VPWR VPWR _07_ _33_/a_109_93# _33_/a_368_53# _33_/a_209_311#
+ _33_/a_296_53# sky130_fd_sc_hd__and3b_1
X_50_ net5 net6 _15_ _11_ VGND VGND VPWR VPWR _22_ _50_/a_515_93# _50_/a_223_47# _50_/a_615_93#
+ _50_/a_343_93# _50_/a_429_93# _50_/a_27_47# sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ net7 net1 net9 net8 VGND VGND VPWR VPWR _06_ _32_/a_109_47# _32_/a_197_47# _32_/a_303_47#
+ _32_/a_27_47# sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_5_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31_ net7 net8 VGND VGND VPWR VPWR _05_ _31_/a_117_297# _31_/a_285_297# _31_/a_285_47#
+ _31_/a_35_297# sky130_fd_sc_hd__xor2_1
X_30_ net9 net10 _03_ net1 VGND VGND VPWR VPWR _04_ _30_/a_465_297# _30_/a_297_297#
+ _30_/a_215_297# _30_/a_392_297# _30_/a_109_53# sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
C0 VPWR _31_/a_285_47# -2.91e-19
C1 net9 _09_ 2.62e-19
C2 _06_ net18 0.0211f
C3 _55_/a_80_21# net3 2.35e-19
C4 _16_ _06_ 0.00162f
C5 _26_/a_29_53# _12_ 0.00243f
C6 b[1] output17/a_27_47# 0.00945f
C7 _50_/a_615_93# net14 1.69e-20
C8 net11 _53_/a_29_53# 8.31e-19
C9 _06_ _43_/a_193_413# 0.0138f
C10 VPWR _44_/a_93_21# 0.005f
C11 _37_/a_27_47# net6 4.3e-20
C12 _11_ input15/a_27_47# 4.4e-19
C13 _10_ _17_ 0.0233f
C14 b[0] output16/a_27_47# 0.014f
C15 _22_ _09_ 0.0279f
C16 p[5] input10/a_27_47# 0.0172f
C17 p[10] _01_ 7.94e-20
C18 net9 net13 0.035f
C19 _55_/a_80_21# _42_/a_209_311# 0.0175f
C20 b[1] input3/a_27_47# 1.31e-20
C21 _42_/a_109_93# net15 4.62e-19
C22 VPWR p[13] 0.183f
C23 _00_ _45_/a_27_47# 4.84e-20
C24 _17_ p[9] 1.03e-20
C25 _22_ net6 0.163f
C26 _36_/a_27_47# _05_ 3.67e-21
C27 _50_/a_223_47# _36_/a_27_47# 1.27e-20
C28 _39_/a_285_47# _12_ 0.0221f
C29 _35_/a_226_47# _45_/a_193_297# 8.15e-21
C30 b[3] _55_/a_80_21# 3.55e-19
C31 _08_ _09_ 0.103f
C32 _36_/a_197_47# _25_ 2.37e-21
C33 net19 _44_/a_250_297# 0.00592f
C34 output17/a_27_47# net8 0.0043f
C35 _34_/a_47_47# net12 0.0385f
C36 _16_ _18_ 0.144f
C37 _21_ net18 0.00215f
C38 output17/a_27_47# _19_ 7.69e-19
C39 net4 _02_ 0.00376f
C40 _44_/a_93_21# net15 0.00573f
C41 _41_/a_59_75# _12_ 0.00101f
C42 p[2] _05_ 3.69e-19
C43 _01_ _35_/a_76_199# 3.08e-21
C44 _04_ _49_/a_201_297# 0.0253f
C45 VPWR _52_/a_346_47# -0.00109f
C46 _43_/a_193_413# _18_ 0.0413f
C47 net18 _24_ 5.57e-21
C48 p[10] p[11] 0.00241f
C49 _27_/a_277_297# VPWR -3.63e-19
C50 _32_/a_27_47# _30_/a_109_53# 1.51e-19
C51 _22_ net13 4.63e-20
C52 input14/a_27_47# p[13] 1.37e-19
C53 _32_/a_197_47# net1 0.00142f
C54 p[13] net15 1.48e-19
C55 net7 p[1] 0.00514f
C56 net5 _55_/a_80_21# 2.78e-19
C57 VPWR _35_/a_556_47# -7.24e-19
C58 p[8] _11_ 7.7e-20
C59 _08_ net13 1.82e-19
C60 _40_/a_297_297# _06_ 1.64e-19
C61 input9/a_75_212# _30_/a_215_297# 6.24e-21
C62 net3 input15/a_27_47# 8.74e-20
C63 _07_ _02_ 0.0083f
C64 b[0] _39_/a_285_47# 1.88e-19
C65 _04_ _06_ 0.0136f
C66 _03_ _07_ 0.0113f
C67 _29_/a_111_297# _09_ 5.79e-20
C68 _15_ _44_/a_250_297# 0.00517f
C69 _32_/a_27_47# net8 0.0275f
C70 input5/a_381_47# net14 0.00479f
C71 VPWR _12_ 0.28f
C72 _27_/a_277_297# net15 1.93e-19
C73 p[14] input6/a_27_47# 0.0155f
C74 net6 _09_ 5.43e-20
C75 _22_ _13_ 0.00309f
C76 VPWR _30_/a_297_297# -4.57e-19
C77 _43_/a_297_47# _06_ 4.81e-20
C78 _03_ _33_/a_209_311# 8.38e-19
C79 net14 _01_ 8.29e-19
C80 _29_/a_29_53# _36_/a_27_47# 6.92e-20
C81 _48_/a_27_47# _07_ 0.0524f
C82 VPWR p[1] 0.08f
C83 _09_ net13 0.0379f
C84 b[3] input15/a_27_47# 1.77e-19
C85 input10/a_27_47# p[6] 0.00214f
C86 net9 _35_/a_226_47# 1.22e-20
C87 _12_ net15 8.14e-21
C88 input3/a_27_47# output17/a_27_47# 3.15e-19
C89 net11 _52_/a_93_21# 2.8e-19
C90 net6 net13 0.00188f
C91 _04_ _18_ 1.94e-21
C92 VPWR _52_/a_250_297# 0.019f
C93 _17_ net4 7.52e-21
C94 _21_ _04_ 0.39f
C95 p[8] net3 2.53e-19
C96 p[2] _31_/a_35_297# 0.00264f
C97 net11 net8 1.5e-19
C98 net11 _19_ 6.27e-21
C99 VPWR b[0] 0.142f
C100 p[11] net14 0.00182f
C101 net10 _33_/a_368_53# 0.00171f
C102 _40_/a_109_297# _14_ -1.78e-33
C103 _10_ output19/a_27_47# 3.23e-20
C104 p[10] _02_ 2.17e-19
C105 _22_ _35_/a_226_47# 1.39e-20
C106 _30_/a_465_297# net12 8.01e-20
C107 _26_/a_111_297# VPWR -5.92e-20
C108 net16 _06_ 0.0511f
C109 net10 _06_ 0.184f
C110 net15 p[1] 6.22e-20
C111 p[10] _03_ 8.74e-20
C112 output19/a_27_47# p[9] 0.0852f
C113 input5/a_381_47# net9 3.4e-19
C114 _10_ _45_/a_465_47# 3.32e-19
C115 _09_ _13_ 0.0927f
C116 _08_ _35_/a_226_47# 0.00117f
C117 _00_ _47_/a_299_297# 7.59e-21
C118 _10_ _47_/a_81_21# 0.0061f
C119 _26_/a_29_53# _11_ 1.09e-19
C120 _35_/a_76_199# _02_ 5.73e-19
C121 _12_ _53_/a_29_53# 3.46e-20
C122 net6 _13_ 0.0106f
C123 p[8] b[3] 0.226f
C124 _03_ _35_/a_76_199# 0.0733f
C125 input6/a_27_47# _17_ 7.13e-22
C126 _10_ _47_/a_384_47# 3.53e-19
C127 _33_/a_296_53# net13 3.71e-20
C128 _50_/a_615_93# net6 1.43e-19
C129 net1 _49_/a_201_297# 0.00304f
C130 _45_/a_109_297# _06_ 0.0023f
C131 net9 _01_ 0.157f
C132 _13_ net13 4e-21
C133 net10 _18_ 1.47e-21
C134 _04_ _50_/a_27_47# 2.07e-21
C135 net16 _18_ 8.17e-21
C136 b[1] p[13] 0.00115f
C137 _21_ net10 0.0254f
C138 _32_/a_303_47# _20_ 1.54e-19
C139 net16 _21_ 1.89e-19
C140 VPWR _54_/a_75_212# 0.0475f
C141 _31_/a_35_297# _55_/a_80_21# 5.9e-21
C142 net5 _30_/a_215_297# 8.27e-21
C143 _37_/a_109_47# net14 1.71e-19
C144 _31_/a_285_47# net8 0.00129f
C145 _42_/a_109_93# _19_ 1.14e-21
C146 net16 _24_ 6.93e-19
C147 _10_ _25_ 0.0109f
C148 _00_ _16_ 0.00613f
C149 net1 _06_ 0.0115f
C150 _22_ _01_ 0.15f
C151 _41_/a_59_75# _11_ 8.7e-19
C152 _33_/a_109_93# input13/a_27_47# 0.00348f
C153 _04_ net12 0.267f
C154 _09_ _35_/a_226_47# 0.058f
C155 _10_ _43_/a_27_47# 0.0279f
C156 _00_ _43_/a_193_413# 0.00721f
C157 _37_/a_27_47# p[11] 4.41e-19
C158 _02_ _45_/a_193_297# 0.00988f
C159 _35_/a_226_297# _12_ 3.35e-20
C160 _03_ _45_/a_193_297# 2.57e-20
C161 net2 input15/a_27_47# 0.00296f
C162 _26_/a_29_53# net3 2.83e-21
C163 net14 _02_ 0.00952f
C164 _38_/a_27_47# output16/a_27_47# 9.02e-19
C165 p[13] net8 0.00345f
C166 _03_ net14 1.5e-19
C167 VPWR _32_/a_109_47# 0.00124f
C168 p[14] net14 6.11e-20
C169 _22_ p[11] 3.13e-20
C170 _04_ net17 0.0218f
C171 VPWR p[5] 0.092f
C172 _35_/a_226_47# net13 0.00709f
C173 VPWR _44_/a_256_47# -7.56e-19
C174 _52_/a_346_47# _52_/a_93_21# -5.12e-20
C175 _28_/a_109_297# _11_ 6.29e-19
C176 _30_/a_215_297# _05_ 0.0453f
C177 _16_ _14_ 0.0584f
C178 _10_ _20_ 0.179f
C179 b[2] _25_ 0.0015f
C180 VPWR _11_ 0.352f
C181 VPWR input9/a_75_212# 0.0641f
C182 _27_/a_277_297# net8 7.99e-20
C183 _21_ net1 0.0252f
C184 net10 _50_/a_27_47# 3.78e-21
C185 output17/a_27_47# _42_/a_109_93# 8.6e-21
C186 net16 _50_/a_27_47# 2.35e-20
C187 net7 net3 7.45e-20
C188 _49_/a_315_47# _49_/a_75_199# 1.78e-33
C189 _06_ _34_/a_377_297# 0.00427f
C190 _14_ _43_/a_193_413# 0.0297f
C191 net5 output16/a_27_47# 4.08e-20
C192 input2/a_27_47# _30_/a_215_297# 3.51e-20
C193 net19 _55_/a_80_21# 0.00423f
C194 net6 _45_/a_205_47# 2.59e-20
C195 p[8] net2 0.00102f
C196 _01_ _09_ 4.69e-21
C197 _39_/a_47_47# _12_ 0.0317f
C198 net10 net12 0.539f
C199 input3/a_27_47# _42_/a_109_93# 0.00249f
C200 _35_/a_226_47# _13_ 5.62e-21
C201 _52_/a_93_21# _12_ 0.0157f
C202 input14/a_27_47# _11_ 1.42e-19
C203 net15 _11_ 0.145f
C204 p[13] output17/a_27_47# 0.00118f
C205 input5/a_841_47# _06_ 1.66e-19
C206 _26_/a_29_53# net5 0.0237f
C207 _00_ _04_ 1.98e-20
C208 input6/a_27_47# output19/a_27_47# 0.107f
C209 _30_/a_297_297# net8 2.42e-21
C210 _00_ _43_/a_297_47# 1.26e-19
C211 net9 _02_ 0.00611f
C212 input8/a_27_47# net9 3.71e-20
C213 net10 net17 8.67e-21
C214 _03_ net9 0.15f
C215 _01_ net13 0.00228f
C216 _21_ _34_/a_377_297# 2.37e-19
C217 _17_ net14 0.104f
C218 p[13] input3/a_27_47# 0.00499f
C219 _26_/a_29_53# _52_/a_584_47# 7.45e-20
C220 VPWR net3 0.351f
C221 VPWR _55_/a_300_47# -4.61e-19
C222 _40_/a_297_297# _14_ 1.58e-19
C223 _37_/a_27_47# p[14] 1.37e-19
C224 _15_ _55_/a_80_21# 0.107f
C225 _39_/a_47_47# b[0] 2.04e-19
C226 _52_/a_93_21# _52_/a_250_297# -6.97e-22
C227 _19_ p[1] 2.82e-20
C228 p[2] _49_/a_201_297# 4.58e-20
C229 net5 net7 0.195f
C230 net5 _39_/a_285_47# 0.0405f
C231 _29_/a_29_53# _30_/a_215_297# 1.72e-19
C232 _22_ _02_ 0.552f
C233 _32_/a_27_47# p[13] 6.49e-20
C234 _31_/a_35_297# _30_/a_215_297# 6.37e-19
C235 _04_ _14_ 2.04e-21
C236 _03_ _22_ 2.55e-20
C237 _11_ _53_/a_29_53# 2.33e-20
C238 _21_ input5/a_841_47# 1.59e-21
C239 net5 _36_/a_109_47# 0.00144f
C240 net5 _41_/a_59_75# 2.41e-19
C241 VPWR p[6] 0.0738f
C242 _45_/a_205_47# _13_ 7.51e-20
C243 _08_ _02_ 2.26e-20
C244 VPWR _42_/a_209_311# -0.00753f
C245 net1 net12 1.17e-19
C246 _26_/a_29_53# _50_/a_223_47# 0.00124f
C247 _06_ _36_/a_27_47# 0.0501f
C248 VPWR _38_/a_27_47# -0.0142f
C249 _29_/a_183_297# net9 3.51e-19
C250 _03_ _08_ 0.0144f
C251 _43_/a_297_47# _14_ 9.11e-19
C252 _28_/a_109_297# b[3] 7.49e-20
C253 input14/a_27_47# net3 9.36e-19
C254 _55_/a_300_47# net15 1.09e-19
C255 net19 input15/a_27_47# 0.00236f
C256 _55_/a_217_297# net3 5.78e-20
C257 net15 net3 0.394f
C258 input5/a_558_47# p[10] 1.09e-19
C259 VPWR b[3] 0.367f
C260 b[2] output18/a_27_47# 0.0141f
C261 _06_ p[7] 0.00864f
C262 net4 _20_ 3.01e-20
C263 _04_ _49_/a_75_199# 0.0782f
C264 net1 net17 2.89e-19
C265 _48_/a_27_47# _08_ 2.58e-19
C266 _05_ net7 0.0129f
C267 VPWR net5 0.612f
C268 net17 input7/a_27_47# 4.99e-20
C269 _42_/a_209_311# net15 0.0157f
C270 _00_ _45_/a_109_297# 4.86e-20
C271 _10_ _45_/a_27_47# 0.0143f
C272 _27_/a_27_297# p[10] 6.35e-19
C273 _18_ _36_/a_27_47# 5.46e-20
C274 input14/a_27_47# b[3] 0.0211f
C275 net9 _17_ 2.89e-23
C276 _36_/a_303_47# _25_ 2.03e-21
C277 b[3] net15 0.00408f
C278 net7 _49_/a_544_297# 2.72e-19
C279 b[3] _55_/a_217_297# 3.41e-19
C280 _00_ _44_/a_250_297# 6.39e-20
C281 _21_ _36_/a_27_47# 0.0276f
C282 _06_ _53_/a_111_297# 3.82e-19
C283 _09_ _02_ 0.297f
C284 _29_/a_111_297# _03_ 7.48e-19
C285 _34_/a_377_297# net12 0.00251f
C286 _03_ _09_ 0.326f
C287 _37_/a_27_47# _17_ 0.00277f
C288 input2/a_27_47# net7 0.00213f
C289 _07_ _20_ 1.28e-21
C290 VPWR _52_/a_584_47# -9.47e-19
C291 _10_ _23_ 0.00192f
C292 _15_ input15/a_27_47# 2.15e-20
C293 net6 _02_ 0.00427f
C294 net2 net7 0.00234f
C295 _03_ net6 2.9e-20
C296 p[8] net19 0.0268f
C297 p[14] net6 0.00237f
C298 net16 _38_/a_109_47# 4.17e-19
C299 net5 net15 0.0226f
C300 _22_ _17_ 0.00334f
C301 net5 _55_/a_217_297# 8.84e-20
C302 _00_ net1 9.43e-19
C303 p[3] input13/a_27_47# 0.00101f
C304 _02_ net13 0.00154f
C305 _29_/a_29_53# _26_/a_29_53# 0.00121f
C306 _06_ _55_/a_80_21# 5.15e-19
C307 _38_/a_27_47# _53_/a_29_53# 1.29e-19
C308 _48_/a_27_47# _09_ 0.00541f
C309 _42_/a_109_93# _44_/a_93_21# 1.25e-19
C310 _03_ net13 0.271f
C311 VPWR _05_ 0.127f
C312 VPWR _50_/a_223_47# -0.00601f
C313 output19/a_27_47# net14 0.00142f
C314 _32_/a_109_47# net8 0.0011f
C315 _29_/a_183_297# _09_ 4.51e-20
C316 input5/a_558_47# net14 0.0325f
C317 _14_ _44_/a_250_297# 4.82e-19
C318 net11 _12_ 0.00799f
C319 _21_ _53_/a_111_297# 4.38e-19
C320 _27_/a_205_297# net3 4.37e-19
C321 _39_/a_47_47# _11_ 3.9e-19
C322 _24_ _53_/a_111_297# 9.08e-21
C323 VPWR _49_/a_544_297# 0.00569f
C324 _43_/a_369_47# _06_ -2.02e-19
C325 b[2] _23_ 2.87e-20
C326 net12 p[4] 5.33e-19
C327 VPWR input2/a_27_47# 0.00872f
C328 _04_ _33_/a_109_93# 0.0299f
C329 _50_/a_27_47# _36_/a_27_47# 6.08e-19
C330 _45_/a_27_47# input4/a_75_212# 2.18e-20
C331 net8 _11_ 1.81e-20
C332 _29_/a_29_53# net7 6.01e-19
C333 _31_/a_35_297# net7 0.0384f
C334 VPWR net2 0.918f
C335 _55_/a_80_21# _18_ 1.44e-20
C336 _02_ _13_ 0.0676f
C337 _27_/a_27_297# net14 0.0118f
C338 _03_ _13_ 1.74e-20
C339 net11 _52_/a_250_297# 1.2e-19
C340 VPWR _52_/a_256_47# -9.47e-19
C341 _36_/a_27_47# net12 0.0185f
C342 _17_ net6 3.12e-19
C343 _35_/a_76_199# _20_ 3.21e-20
C344 input2/a_27_47# net15 1.61e-19
C345 _43_/a_369_47# _18_ 1.49e-19
C346 input14/a_27_47# net2 0.0176f
C347 net2 net15 0.324f
C348 net12 p[7] 0.0343f
C349 net1 _49_/a_75_199# 0.00799f
C350 _45_/a_27_47# net4 0.024f
C351 _26_/a_183_297# VPWR -3.03e-19
C352 _39_/a_47_47# net3 1.66e-20
C353 _06_ input15/a_27_47# 4.73e-19
C354 _29_/a_29_53# VPWR 0.0299f
C355 VPWR _31_/a_35_297# 0.0333f
C356 _43_/a_27_47# net14 4.87e-20
C357 input5/a_558_47# net9 4.42e-19
C358 net10 _33_/a_109_93# 0.0336f
C359 _35_/a_226_47# _02_ 2.21e-19
C360 _10_ _47_/a_299_297# 0.0134f
C361 net8 net3 9.23e-19
C362 b[1] b[3] 6.12e-20
C363 _06_ _35_/a_489_413# 9.22e-19
C364 _03_ _35_/a_226_47# 0.028f
C365 net3 _19_ 0.0129f
C366 _45_/a_27_47# _07_ 1.02e-20
C367 _47_/a_81_21# net9 3.49e-19
C368 _00_ _39_/a_129_47# 1.63e-20
C369 _18_ input15/a_27_47# 8.27e-21
C370 _37_/a_197_47# net14 7e-19
C371 net11 _54_/a_75_212# 0.00956f
C372 net14 _20_ 8.01e-20
C373 net19 _41_/a_59_75# 3.1e-20
C374 net5 _30_/a_109_53# 5.84e-22
C375 _07_ _23_ 1.27e-19
C376 _42_/a_209_311# net8 7.7e-21
C377 _26_/a_29_53# _15_ 0.00192f
C378 _48_/a_109_47# _06_ 9.47e-19
C379 _06_ _30_/a_215_297# 2.03e-20
C380 _32_/a_27_47# _11_ 1.65e-20
C381 _10_ _16_ 0.00486f
C382 _52_/a_346_47# _12_ 3.8e-19
C383 _47_/a_81_21# _22_ 7.25e-19
C384 _34_/a_285_47# p[6] 8.31e-20
C385 net5 _39_/a_47_47# 0.0352f
C386 _33_/a_209_311# input13/a_27_47# 5.85e-20
C387 _21_ _35_/a_489_413# 0.0448f
C388 _10_ _43_/a_193_413# 0.0174f
C389 _37_/a_109_47# p[11] 2.84e-20
C390 net5 _52_/a_93_21# 0.0124f
C391 output17/a_27_47# net3 0.00248f
C392 _15_ net7 8.4e-20
C393 _01_ _02_ 0.106f
C394 net5 net8 0.48f
C395 net5 _19_ 6.41e-21
C396 input8/a_27_47# _01_ 1.43e-19
C397 _03_ _01_ 2.85e-19
C398 _43_/a_193_413# p[9] 1.09e-19
C399 VPWR _32_/a_197_47# 0.00146f
C400 VPWR net19 0.181f
C401 net11 p[5] 0.0598f
C402 VPWR _44_/a_346_47# -8.74e-19
C403 _15_ _41_/a_59_75# 0.0139f
C404 b[1] _05_ 5.29e-20
C405 _22_ _25_ 5.39e-19
C406 b[2] net18 0.0131f
C407 _21_ _30_/a_215_297# 1.48e-19
C408 _30_/a_109_53# _05_ 0.033f
C409 input3/a_27_47# net3 0.03f
C410 output19/a_27_47# net6 0.00112f
C411 p[14] p[11] 3.13e-20
C412 input9/a_75_212# net11 1.1e-20
C413 _22_ _43_/a_27_47# 0.091f
C414 _45_/a_27_47# _35_/a_76_199# 2.04e-21
C415 _07_ _34_/a_47_47# 0.011f
C416 _06_ _34_/a_129_47# 5.3e-19
C417 b[3] output17/a_27_47# 4.01e-20
C418 _09_ _45_/a_465_47# 2.77e-19
C419 b[1] input2/a_27_47# 8.55e-19
C420 net9 _20_ 0.328f
C421 net19 net15 0.0501f
C422 input14/a_27_47# net19 1.44e-19
C423 input2/a_27_47# _30_/a_109_53# 1.54e-20
C424 b[1] net2 0.0191f
C425 net10 _31_/a_285_297# 1.68e-19
C426 net6 _45_/a_465_47# 6.06e-20
C427 p[0] p[10] 8.21e-20
C428 _05_ _52_/a_93_21# 1.12e-20
C429 _39_/a_377_297# _12_ 6.77e-19
C430 _28_/a_109_297# _15_ 0.00346f
C431 _00_ _55_/a_80_21# 5.5e-19
C432 _47_/a_299_297# net4 3.28e-19
C433 _47_/a_81_21# net6 2.14e-19
C434 _34_/a_47_47# _33_/a_209_311# 0.017f
C435 input3/a_27_47# _42_/a_209_311# 1.56e-19
C436 _05_ net8 0.0146f
C437 _52_/a_250_297# _12_ 0.0139f
C438 VPWR _15_ 0.912f
C439 _10_ _04_ 9.24e-20
C440 input5/a_62_47# net14 5.28e-20
C441 input3/a_27_47# b[3] 0.012f
C442 b[0] _12_ 2.61e-20
C443 p[2] _49_/a_75_199# 1.06e-19
C444 net5 output17/a_27_47# 5.01e-20
C445 _22_ _20_ 0.183f
C446 _49_/a_201_297# net7 0.00419f
C447 _26_/a_29_53# _06_ 0.0135f
C448 net12 input10/a_27_47# 0.00115f
C449 _35_/a_489_413# net12 3.97e-20
C450 _10_ _43_/a_297_47# 0.00118f
C451 _04_ p[3] 8.93e-22
C452 input2/a_27_47# _19_ 5.26e-20
C453 input2/a_27_47# net8 0.0207f
C454 _34_/a_285_47# _05_ 7.85e-21
C455 _17_ _01_ 1.46e-20
C456 _09_ _25_ 1.49e-19
C457 net2 net8 0.0525f
C458 net2 _19_ 0.101f
C459 _15_ net15 0.156f
C460 _14_ _55_/a_80_21# 0.0175f
C461 _16_ net4 2.73e-20
C462 _15_ _55_/a_217_297# 0.0474f
C463 _52_/a_93_21# _52_/a_256_47# -6.6e-20
C464 b[1] _31_/a_35_297# 3.21e-19
C465 _29_/a_29_53# _30_/a_109_53# 0.0103f
C466 _44_/a_256_47# _44_/a_93_21# -6.6e-20
C467 _43_/a_27_47# net6 9.07e-20
C468 _31_/a_35_297# _30_/a_109_53# 2.89e-20
C469 _06_ net7 0.00447f
C470 _06_ _39_/a_285_47# 1.23e-20
C471 _32_/a_27_47# net5 0.0961f
C472 p[11] _17_ 1.93e-19
C473 net11 p[6] 0.0099f
C474 net1 _31_/a_285_297# 5.85e-19
C475 _30_/a_215_297# net12 0.00676f
C476 _44_/a_93_21# _11_ 4.78e-20
C477 _45_/a_193_297# _23_ 4.13e-19
C478 _45_/a_465_47# _13_ 0.00134f
C479 _38_/a_27_47# net11 1.68e-20
C480 _26_/a_29_53# _50_/a_343_93# 2.61e-19
C481 _26_/a_29_53# _18_ 5.26e-20
C482 _25_ net13 0.00297f
C483 output17/a_27_47# _05_ 1.12e-19
C484 VPWR _42_/a_296_53# -6.37e-20
C485 _06_ _36_/a_109_47# 0.00168f
C486 _06_ _41_/a_59_75# 0.0429f
C487 input8/a_27_47# _02_ 5.08e-20
C488 _43_/a_369_47# _14_ 0.00135f
C489 _03_ _02_ 0.00474f
C490 VPWR _49_/a_201_297# 0.0185f
C491 _10_ net10 4.45e-19
C492 _10_ net16 0.0338f
C493 _26_/a_29_53# _24_ 2.11e-20
C494 net1 _32_/a_303_47# 1.45e-19
C495 _22_ output18/a_27_47# 7.51e-19
C496 _09_ _20_ 7.11e-19
C497 net17 _30_/a_215_297# 4.69e-20
C498 _31_/a_35_297# net8 0.0408f
C499 input5/a_62_47# net9 3.12e-19
C500 _31_/a_35_297# _19_ 1.47e-19
C501 input2/a_27_47# output17/a_27_47# 0.107f
C502 net6 _20_ 9.69e-20
C503 net10 p[3] 8.58e-19
C504 net2 output17/a_27_47# 0.0285f
C505 _18_ net7 2.58e-20
C506 VPWR _33_/a_368_53# -4.26e-19
C507 _21_ net7 3e-19
C508 _48_/a_27_47# _02_ 0.00435f
C509 _42_/a_109_93# net3 0.0435f
C510 net5 net11 0.0129f
C511 _33_/a_109_93# p[7] 1.15e-19
C512 _10_ _45_/a_109_297# 0.00202f
C513 _32_/a_27_47# _05_ 2.2e-20
C514 VPWR _06_ 1.4f
C515 _40_/a_191_297# net6 1.16e-20
C516 _41_/a_59_75# _50_/a_343_93# 6.13e-22
C517 _49_/a_201_297# net15 1.41e-19
C518 b[3] _55_/a_472_297# 1.51e-19
C519 _20_ net13 5.95e-19
C520 _06_ _53_/a_183_297# 0.00146f
C521 _29_/a_183_297# _03_ 7.36e-19
C522 net2 input3/a_27_47# 0.0222f
C523 _37_/a_109_47# _17_ 8.86e-21
C524 _43_/a_27_47# _13_ 1.66e-20
C525 _44_/a_93_21# net3 0.0102f
C526 _14_ input15/a_27_47# 9.48e-21
C527 _26_/a_29_53# _50_/a_27_47# 5.56e-19
C528 net16 _38_/a_197_47# 5.89e-19
C529 p[13] net3 3.65e-19
C530 _27_/a_205_297# _15_ 5.5e-20
C531 _12_ _11_ 0.195f
C532 _10_ net1 4.34e-19
C533 net9 input13/a_27_47# 2.42e-19
C534 net9 _23_ 1.21e-19
C535 b[3] _42_/a_109_93# 3.29e-19
C536 input12/a_27_47# _02_ 1.88e-19
C537 _06_ _55_/a_217_297# 3.46e-19
C538 _45_/a_27_47# _22_ 0.0131f
C539 _06_ net15 0.033f
C540 _42_/a_209_311# _44_/a_93_21# 2.21e-19
C541 VPWR _50_/a_343_93# -0.0126f
C542 _17_ _02_ 0.00482f
C543 VPWR _18_ 0.0721f
C544 _13_ _20_ 7.38e-21
C545 net11 _05_ 2.76e-19
C546 net1 p[3] 6.54e-19
C547 _04_ _07_ 9.74e-20
C548 _26_/a_29_53# net12 6.55e-19
C549 _21_ VPWR 0.871f
C550 p[14] _17_ 5.46e-21
C551 net19 net8 1.15e-19
C552 input5/a_558_47# _01_ 3.97e-20
C553 _32_/a_197_47# net8 3.39e-20
C554 b[3] _44_/a_93_21# 0.00491f
C555 input5/a_664_47# net14 0.0179f
C556 _50_/a_615_93# _20_ 8.8e-19
C557 VPWR _24_ 0.0129f
C558 _39_/a_377_297# _11_ 2.57e-20
C559 _27_/a_277_297# net3 2.71e-19
C560 _27_/a_27_297# input5/a_381_47# 1.47e-19
C561 net5 _42_/a_109_93# 0.00109f
C562 _22_ _23_ 0.0186f
C563 _04_ _33_/a_209_311# 0.00133f
C564 p[13] b[3] 0.165f
C565 _50_/a_27_47# _41_/a_59_75# 9.59e-22
C566 _31_/a_117_297# net7 0.00472f
C567 net5 _44_/a_93_21# 3.61e-20
C568 _08_ _23_ 1.81e-19
C569 _18_ net15 0.0382f
C570 _47_/a_81_21# _01_ 6.05e-21
C571 net12 net7 1.57e-19
C572 _06_ _53_/a_29_53# 0.0709f
C573 _27_/a_27_297# _01_ 8.04e-19
C574 _27_/a_109_297# net14 1.32e-19
C575 _32_/a_27_47# _31_/a_35_297# 9.17e-20
C576 net10 net4 8.28e-22
C577 net16 net4 0.155f
C578 p[13] net5 0.0069f
C579 _12_ net3 3.09e-20
C580 p[2] _31_/a_285_297# 0.00156f
C581 net9 _34_/a_47_47# 1.41e-20
C582 _35_/a_226_47# _20_ 5.19e-20
C583 net17 net7 0.2f
C584 _15_ net8 1.79e-19
C585 _15_ _19_ 1.46e-20
C586 _43_/a_469_47# _18_ 1.59e-19
C587 _45_/a_27_47# _09_ 0.00823f
C588 _45_/a_109_297# net4 6.43e-20
C589 VPWR _50_/a_27_47# -0.00335f
C590 _45_/a_27_47# net6 0.021f
C591 net10 _07_ 0.057f
C592 net5 _52_/a_346_47# 7.03e-19
C593 p[10] _04_ 0.00306f
C594 _05_ _31_/a_285_47# 5.61e-19
C595 _16_ net14 0.00266f
C596 _38_/a_27_47# _12_ 0.0527f
C597 _00_ _26_/a_29_53# 0.0466f
C598 _43_/a_27_47# _01_ 9.77e-20
C599 _29_/a_29_53# net11 0.00514f
C600 _34_/a_47_47# _22_ 3.9e-21
C601 _43_/a_193_413# net14 1.11e-19
C602 _09_ _23_ 0.207f
C603 _09_ input13/a_27_47# 1.27e-21
C604 VPWR _31_/a_117_297# 8.41e-19
C605 input5/a_664_47# net9 5.29e-19
C606 _21_ _53_/a_29_53# 0.00959f
C607 net10 _33_/a_209_311# 0.0419f
C608 net6 _23_ 2.13e-19
C609 _24_ _53_/a_29_53# 0.0835f
C610 _54_/a_75_212# _11_ 3.22e-20
C611 _04_ _35_/a_76_199# 0.0269f
C612 input3/a_27_47# net19 0.00105f
C613 VPWR net12 0.817f
C614 _06_ _35_/a_226_297# 1.28e-19
C615 _34_/a_47_47# _08_ 0.00123f
C616 net2 _42_/a_109_93# 0.00507f
C617 _00_ net7 8.12e-21
C618 net5 _12_ 0.983f
C619 _00_ _39_/a_285_47# 1.47e-21
C620 _10_ _39_/a_129_47# 2.51e-19
C621 _23_ net13 4.11e-19
C622 input13/a_27_47# net13 0.00139f
C623 VPWR net17 0.0371f
C624 net2 _44_/a_93_21# 0.0273f
C625 _10_ _36_/a_27_47# 0.00109f
C626 _01_ _20_ 0.161f
C627 _37_/a_303_47# net14 0.00112f
C628 _26_/a_29_53# _14_ 3.67e-19
C629 _00_ _41_/a_59_75# 2.43e-20
C630 _48_/a_181_47# _06_ 6.4e-19
C631 net8 _49_/a_201_297# 7.3e-19
C632 _06_ _30_/a_109_53# 1.96e-19
C633 p[13] net2 0.0247f
C634 _45_/a_27_47# _13_ 0.0703f
C635 p[14] output19/a_27_47# 0.0932f
C636 p[12] input15/a_27_47# 5.48e-19
C637 net1 _07_ 6.08e-22
C638 _40_/a_109_297# net6 2.53e-20
C639 net5 _39_/a_377_297# 0.00234f
C640 input3/a_27_47# _15_ 7.53e-19
C641 _30_/a_215_297# _33_/a_109_93# 0.00104f
C642 _37_/a_197_47# p[11] 1.59e-19
C643 net5 _52_/a_250_297# 0.018f
C644 _39_/a_47_47# _06_ 1.44e-19
C645 net17 net15 5.19e-19
C646 _47_/a_81_21# _02_ 1.59e-20
C647 p[2] p[3] 0.188f
C648 _14_ net7 0.00251f
C649 _13_ _23_ 2.08e-20
C650 net5 b[0] 2.76e-19
C651 p[3] p[7] 0.169f
C652 _27_/a_27_297# _02_ 0.00179f
C653 net10 _35_/a_76_199# 0.0146f
C654 _04_ net14 0.0863f
C655 _06_ _52_/a_93_21# 0.0574f
C656 _37_/a_27_47# _16_ 2.07e-19
C657 _30_/a_465_297# net9 0.00138f
C658 _27_/a_27_297# _03_ 2.68e-19
C659 _32_/a_27_47# _15_ 1.19e-19
C660 _50_/a_223_47# _12_ 0.00327f
C661 _06_ net8 0.00282f
C662 _05_ _12_ 2.52e-19
C663 _00_ VPWR 0.416f
C664 _37_/a_27_47# _43_/a_193_413# 0.0102f
C665 VPWR _44_/a_584_47# -2.28e-19
C666 _10_ _53_/a_111_297# 2.06e-19
C667 _43_/a_297_47# net14 1.09e-21
C668 _22_ net18 1.68e-19
C669 _21_ _30_/a_109_53# 3.31e-20
C670 _34_/a_47_47# net13 1.68e-19
C671 _16_ _22_ 3.8e-19
C672 _38_/a_27_47# _54_/a_75_212# 2.67e-19
C673 _22_ _43_/a_193_413# 0.00133f
C674 net7 _49_/a_75_199# 0.09f
C675 _45_/a_27_47# _35_/a_226_47# 5.71e-21
C676 _07_ _34_/a_377_297# 5.8e-19
C677 _06_ _34_/a_285_47# 0.00598f
C678 _39_/a_47_47# _18_ 1.23e-19
C679 _25_ _02_ 0.0156f
C680 _03_ _25_ 0.00422f
C681 net2 _12_ 1.02e-20
C682 _18_ _52_/a_93_21# 1.97e-19
C683 _05_ _52_/a_250_297# 8.86e-22
C684 _43_/a_27_47# _02_ 1.88e-21
C685 _28_/a_109_297# _14_ 5.66e-19
C686 _10_ _55_/a_80_21# 5.49e-19
C687 _00_ net15 0.00147f
C688 net1 p[10] 1.22e-19
C689 _18_ net8 1.15e-21
C690 _44_/a_256_47# net3 0.00101f
C691 _21_ _52_/a_93_21# 9.4e-19
C692 _47_/a_299_297# net6 3.63e-19
C693 _50_/a_343_93# net8 7.25e-19
C694 _35_/a_226_47# _23_ 4.21e-19
C695 output19/a_27_47# _17_ 0.00122f
C696 input5/a_558_47# _17_ 2.13e-21
C697 _35_/a_226_47# input13/a_27_47# 3.94e-20
C698 _21_ net8 0.00656f
C699 _52_/a_93_21# _24_ 0.0211f
C700 net3 _11_ 0.165f
C701 VPWR _14_ 0.186f
C702 input2/a_27_47# p[1] 0.0119f
C703 _49_/a_315_47# _09_ 1.11e-20
C704 net16 _45_/a_193_297# 0.00187f
C705 net2 p[1] 5.99e-20
C706 VPWR _38_/a_109_47# -4.66e-19
C707 _10_ _43_/a_369_47# 0.00199f
C708 net19 _42_/a_109_93# 0.0448f
C709 p[5] p[6] 0.198f
C710 _04_ net9 0.0213f
C711 _21_ _34_/a_285_47# 6.94e-20
C712 _47_/a_81_21# _17_ 0.0456f
C713 _02_ _20_ 0.1f
C714 net4 _36_/a_27_47# 0.0103f
C715 _09_ net18 1.97e-21
C716 _27_/a_27_297# _17_ 6.78e-22
C717 input5/a_62_47# p[11] 0.00153f
C718 _17_ _47_/a_384_47# 1.1e-20
C719 _03_ _20_ 0.0794f
C720 _38_/a_27_47# _11_ 0.071f
C721 VPWR _49_/a_75_199# 0.0177f
C722 _14_ _55_/a_217_297# 0.0116f
C723 _15_ _55_/a_472_297# 0.00626f
C724 net19 _44_/a_93_21# 0.0074f
C725 _14_ net15 0.0538f
C726 _16_ net6 1.62e-20
C727 b[3] _11_ 2.37e-20
C728 b[1] _31_/a_117_297# 2.34e-19
C729 _44_/a_346_47# _44_/a_93_21# -5.12e-20
C730 _43_/a_193_413# net6 2.41e-20
C731 _32_/a_109_47# net5 5.69e-21
C732 _04_ _22_ 1.76e-20
C733 _30_/a_109_53# net12 4.25e-20
C734 _44_/a_250_297# net14 4.24e-20
C735 _32_/a_27_47# _06_ 0.00663f
C736 _04_ _08_ 5.99e-19
C737 VPWR _42_/a_368_53# -3.03e-19
C738 _43_/a_469_47# _14_ 0.00259f
C739 _15_ _42_/a_109_93# 0.00367f
C740 net5 _11_ 0.207f
C741 net15 _49_/a_75_199# 5.13e-20
C742 net11 _49_/a_201_297# 1.42e-19
C743 _10_ input15/a_27_47# 4.5e-19
C744 b[1] net17 0.00766f
C745 _30_/a_465_297# net13 6.36e-20
C746 net1 net14 6.64e-20
C747 net17 _30_/a_109_53# 4.18e-20
C748 _43_/a_27_47# _17_ 0.00131f
C749 net4 _53_/a_111_297# 2.09e-19
C750 _31_/a_117_297# net8 5.91e-19
C751 _15_ _44_/a_93_21# 0.0168f
C752 net14 input7/a_27_47# 3.48e-19
C753 net10 net9 0.111f
C754 net12 net8 0.00458f
C755 output18/a_27_47# _02_ 3.6e-19
C756 p[9] input15/a_27_47# 0.0196f
C757 _10_ _35_/a_489_413# 3.41e-19
C758 _33_/a_209_311# p[7] 1.34e-19
C759 _42_/a_209_311# net3 0.029f
C760 _32_/a_27_47# _50_/a_343_93# 6.48e-20
C761 _32_/a_27_47# _18_ 1.18e-20
C762 _21_ _32_/a_27_47# 8.95e-19
C763 net11 _06_ 0.546f
C764 _40_/a_297_297# net6 7.47e-22
C765 b[3] net3 0.0026f
C766 _55_/a_80_21# net4 1.06e-19
C767 net17 net8 0.18f
C768 _29_/a_111_297# _04_ 9.25e-19
C769 _34_/a_285_47# net12 8.07e-20
C770 _37_/a_197_47# _17_ 9.19e-21
C771 _43_/a_193_413# _13_ 5.58e-21
C772 _17_ _20_ 0.102f
C773 net17 _19_ 0.0211f
C774 _04_ _09_ 0.0904f
C775 net16 _22_ 0.00606f
C776 _04_ net6 2.61e-20
C777 _50_/a_223_47# _11_ 0.0329f
C778 p[12] _41_/a_59_75# 0.0547f
C779 VPWR _33_/a_109_93# -0.00817f
C780 input9/a_75_212# _05_ 1.24e-21
C781 _00_ _30_/a_109_53# 3.67e-20
C782 net10 _08_ 0.189f
C783 _10_ _30_/a_215_297# 5.66e-20
C784 net16 _38_/a_303_47# 6.47e-19
C785 net5 net3 0.0365f
C786 b[3] _42_/a_209_311# 3.71e-19
C787 _43_/a_297_47# net6 8.23e-22
C788 _40_/a_191_297# _17_ 4.35e-19
C789 p[8] p[9] 0.0518f
C790 _45_/a_109_297# _22_ 0.0425f
C791 input4/a_75_212# input15/a_27_47# 1.1e-21
C792 p[3] _30_/a_215_297# 2.01e-19
C793 _04_ net13 0.569f
C794 VPWR _36_/a_197_47# -5.24e-19
C795 _00_ _39_/a_47_47# 1.85e-20
C796 VPWR _50_/a_429_93# -3.61e-19
C797 _36_/a_27_47# _35_/a_76_199# 3.22e-19
C798 _21_ net11 0.586f
C799 net1 net9 0.47f
C800 net2 _11_ 0.234f
C801 net5 _38_/a_27_47# 1.76e-19
C802 _27_/a_27_297# input5/a_558_47# 1.57e-19
C803 net5 _42_/a_209_311# 3.27e-21
C804 _45_/a_27_47# _02_ 0.00449f
C805 VPWR p[12] 0.0375f
C806 _15_ _12_ 0.00833f
C807 _00_ net8 3.23e-19
C808 _45_/a_27_47# _03_ 2.06e-20
C809 _06_ _42_/a_109_93# 5.53e-20
C810 output17/a_27_47# net17 0.0149f
C811 _31_/a_285_297# net7 0.00227f
C812 net1 _22_ 0.0129f
C813 net10 _09_ 0.037f
C814 net16 _09_ 0.00707f
C815 _02_ _23_ 0.0641f
C816 _03_ _23_ 0.0564f
C817 net10 net6 1.35e-20
C818 _04_ _13_ 1.17e-21
C819 net16 net6 8.27e-20
C820 _32_/a_27_47# net12 1.52e-19
C821 _49_/a_315_47# _01_ 1.82e-19
C822 p[12] net15 2.99e-19
C823 _41_/a_145_75# VPWR -2.46e-19
C824 _29_/a_29_53# input9/a_75_212# 9.7e-21
C825 _14_ net8 4.23e-19
C826 _14_ _19_ 2.71e-21
C827 net10 net13 0.375f
C828 net11 _50_/a_27_47# 6.05e-21
C829 net2 net3 0.519f
C830 _45_/a_109_297# net6 7.82e-19
C831 net5 _52_/a_584_47# 0.0022f
C832 _10_ _26_/a_29_53# 0.0265f
C833 _16_ _01_ 3.24e-19
C834 _06_ _52_/a_346_47# 0.0031f
C835 input6/a_27_47# input15/a_27_47# 5.3e-19
C836 VPWR _31_/a_285_297# 0.0174f
C837 _18_ _44_/a_93_21# 0.00485f
C838 _43_/a_193_413# _01_ 8.16e-19
C839 input5/a_841_47# net9 2.7e-19
C840 input2/a_27_47# _42_/a_209_311# 1e-22
C841 net10 _33_/a_296_53# 8.22e-20
C842 net11 net12 0.358f
C843 net8 _49_/a_75_199# 0.00214f
C844 _04_ _35_/a_226_47# 0.00551f
C845 _07_ _35_/a_489_413# 0.00429f
C846 _37_/a_27_47# input5/a_841_47# 4.64e-20
C847 net2 _42_/a_209_311# 5.1e-19
C848 net1 _09_ 5.26e-20
C849 _19_ _49_/a_75_199# 0.0206f
C850 _34_/a_47_47# _02_ 1.09e-19
C851 _45_/a_27_47# _17_ 1.16e-20
C852 _16_ p[11] 2.17e-20
C853 net5 _50_/a_223_47# 0.00202f
C854 _03_ _34_/a_47_47# 4.5e-20
C855 net10 _13_ 4.52e-21
C856 VPWR _32_/a_303_47# 6.03e-19
C857 net2 b[3] 0.311f
C858 net16 _13_ 0.0198f
C859 _10_ net7 6.22e-20
C860 _10_ _39_/a_285_47# 0.00289f
C861 _35_/a_489_413# _33_/a_209_311# 2.77e-20
C862 _47_/a_81_21# _20_ 0.0457f
C863 _29_/a_29_53# net3 1.68e-20
C864 net11 net17 3.19e-20
C865 _00_ _32_/a_27_47# 0.00228f
C866 _10_ _41_/a_59_75# 0.0172f
C867 _06_ _12_ 0.136f
C868 _27_/a_27_297# _20_ 3.14e-20
C869 _47_/a_384_47# _20_ 1.72e-19
C870 net1 net13 3.51e-19
C871 _48_/a_109_47# _07_ 3.01e-19
C872 input5/a_664_47# _02_ 0.00187f
C873 net5 net2 0.0616f
C874 _48_/a_27_47# _34_/a_47_47# 4.45e-21
C875 net19 _11_ 2.19e-19
C876 p[8] input6/a_27_47# 0.00139f
C877 net9 _36_/a_27_47# 0.00493f
C878 _41_/a_59_75# p[9] 1.02e-19
C879 _21_ _35_/a_556_47# 2.69e-19
C880 _37_/a_303_47# p[11] 1.04e-19
C881 _55_/a_80_21# net14 4.7e-19
C882 _30_/a_215_297# _33_/a_209_311# 1.56e-19
C883 _39_/a_377_297# _06_ 8.76e-20
C884 p[2] net9 1.4e-20
C885 _10_ _28_/a_109_297# 4.34e-19
C886 _06_ _52_/a_250_297# 0.0058f
C887 net9 p[7] 8.26e-19
C888 net10 _35_/a_226_47# 0.0159f
C889 _04_ _01_ 0.119f
C890 _18_ _12_ 0.0115f
C891 _50_/a_343_93# _12_ 5.63e-20
C892 _27_/a_109_297# _03_ 1.97e-20
C893 _40_/a_109_297# _17_ 9.67e-19
C894 _10_ VPWR 0.577f
C895 output16/a_27_47# net4 0.00706f
C896 _49_/a_315_47# _02_ 0.00134f
C897 _43_/a_27_47# _20_ 0.0124f
C898 _22_ _36_/a_27_47# 2.82e-20
C899 _21_ _12_ 7.99e-20
C900 _10_ _53_/a_183_297# 2.86e-19
C901 _49_/a_315_47# _03_ 9.22e-19
C902 _43_/a_369_47# net14 6.79e-21
C903 _33_/a_109_93# _52_/a_93_21# 2.89e-21
C904 _12_ _24_ 1.67e-19
C905 _34_/a_47_47# input12/a_27_47# 2.17e-19
C906 input2/a_27_47# _05_ 1.83e-19
C907 _26_/a_111_297# _06_ 9e-19
C908 VPWR p[3] 0.0874f
C909 net17 _42_/a_109_93# 3.1e-21
C910 _29_/a_29_53# net5 8.1e-20
C911 VPWR p[9] 0.374f
C912 _15_ _11_ 0.113f
C913 net17 _31_/a_285_47# 0.00134f
C914 net2 _05_ 4.03e-20
C915 net5 _31_/a_35_297# 2.04e-21
C916 _45_/a_109_297# _35_/a_226_47# 1.59e-21
C917 net18 _02_ 6.8e-20
C918 _03_ net18 2.07e-21
C919 _16_ _02_ 0.00564f
C920 _26_/a_29_53# net4 0.00412f
C921 input4/a_75_212# _41_/a_59_75# 0.00153f
C922 _18_ _52_/a_250_297# 1.77e-19
C923 net19 net3 0.611f
C924 _43_/a_193_413# _02_ 9.4e-21
C925 _10_ _55_/a_217_297# 1.43e-19
C926 _10_ net15 0.0101f
C927 net2 input2/a_27_47# 0.024f
C928 _44_/a_346_47# net3 8.04e-19
C929 p[12] _39_/a_47_47# 3.32e-19
C930 _30_/a_465_297# _03_ 7.72e-19
C931 _52_/a_250_297# _24_ 3.03e-19
C932 VPWR b[2] 0.262f
C933 _22_ _53_/a_111_297# 4.7e-20
C934 input14/a_27_47# p[9] 8.53e-21
C935 output18/a_27_47# _25_ 0.072f
C936 net15 p[9] 0.00306f
C937 net1 _35_/a_226_47# 1.3e-20
C938 VPWR _38_/a_197_47# -5.24e-19
C939 net19 _42_/a_209_311# 0.0766f
C940 _10_ _43_/a_469_47# 0.00124f
C941 _50_/a_27_47# _12_ 0.00354f
C942 _06_ _54_/a_75_212# 0.00727f
C943 _40_/a_191_297# _20_ 2.07e-20
C944 _39_/a_129_47# net6 6.91e-19
C945 _39_/a_285_47# net4 9.71e-19
C946 _29_/a_29_53# _50_/a_223_47# 1.45e-20
C947 p[4] net13 2.34e-20
C948 _29_/a_29_53# _05_ 3.79e-20
C949 net19 b[3] 0.0439f
C950 VPWR input4/a_75_212# 0.06f
C951 _31_/a_35_297# _05_ 0.00649f
C952 net6 _36_/a_27_47# 5.1e-19
C953 _41_/a_59_75# net4 1.76e-19
C954 _10_ _53_/a_29_53# 0.00779f
C955 _15_ net3 0.224f
C956 net11 _49_/a_75_199# 4.49e-19
C957 _15_ _55_/a_300_47# 1.42e-20
C958 _14_ _55_/a_472_297# 0.00192f
C959 _22_ _55_/a_80_21# 0.00926f
C960 _09_ p[7] 9.25e-21
C961 _00_ _44_/a_93_21# 4.54e-20
C962 b[1] _31_/a_285_297# 1.12e-19
C963 net12 _12_ 7.94e-21
C964 _32_/a_197_47# net5 5.61e-21
C965 net5 net19 0.00124f
C966 _31_/a_35_297# input2/a_27_47# 0.00136f
C967 _36_/a_27_47# net13 0.0488f
C968 input5/a_381_47# net1 1.27e-19
C969 _31_/a_35_297# net2 0.0635f
C970 _30_/a_297_297# net12 7.14e-21
C971 _14_ _42_/a_109_93# 0.00141f
C972 _15_ _42_/a_209_311# 0.0521f
C973 _04_ _02_ 0.0541f
C974 _16_ _17_ 0.242f
C975 p[8] net14 0.00868f
C976 _04_ input8/a_27_47# 2.36e-22
C977 p[7] net13 0.00809f
C978 _03_ _04_ 0.586f
C979 _09_ _53_/a_111_297# 3.4e-19
C980 VPWR net4 1.07f
C981 _43_/a_193_413# _17_ 0.0503f
C982 _15_ b[3] 0.00162f
C983 net1 _01_ 0.0509f
C984 _06_ _11_ 0.493f
C985 _44_/a_250_297# p[11] 1.13e-19
C986 _31_/a_285_297# net8 0.0215f
C987 _14_ _44_/a_93_21# 0.04f
C988 b[2] _53_/a_29_53# 6.22e-19
C989 _31_/a_285_297# _19_ 1.34e-19
C990 net17 p[1] 6.65e-20
C991 _42_/a_296_53# net3 1.81e-19
C992 _25_ _23_ 0.00465f
C993 _37_/a_27_47# input15/a_27_47# 3.27e-19
C994 net5 _15_ 0.0352f
C995 _32_/a_303_47# net8 2.22e-34
C996 VPWR _07_ 0.0728f
C997 net4 net15 8.68e-19
C998 _55_/a_217_297# net4 1.13e-19
C999 VPWR input6/a_27_47# 0.00162f
C1000 _29_/a_183_297# _04_ 0.0015f
C1001 _37_/a_303_47# _17_ 1.23e-20
C1002 p[10] net7 0.00481f
C1003 _18_ _11_ 0.484f
C1004 _50_/a_343_93# _11_ 0.0384f
C1005 _00_ _12_ 0.00396f
C1006 net11 _33_/a_109_93# 5.14e-19
C1007 VPWR _33_/a_209_311# -0.0131f
C1008 _21_ _11_ 9.98e-20
C1009 _21_ input9/a_75_212# 1.17e-21
C1010 input2/a_27_47# net19 2.9e-23
C1011 _24_ _11_ 7.29e-20
C1012 net10 _02_ 3.52e-19
C1013 net16 _02_ 8.94e-19
C1014 net2 net19 0.599f
C1015 _35_/a_76_199# net7 1.79e-20
C1016 net10 _03_ 0.32f
C1017 _43_/a_369_47# net6 3.62e-21
C1018 _06_ _55_/a_300_47# 2.5e-20
C1019 _06_ net3 0.0072f
C1020 VPWR _36_/a_303_47# -4.83e-19
C1021 net2 _44_/a_346_47# 1.64e-19
C1022 _10_ _39_/a_47_47# 0.00824f
C1023 p[3] _30_/a_109_53# 3.23e-20
C1024 net9 _30_/a_215_297# 0.0458f
C1025 VPWR _50_/a_515_93# -5.03e-19
C1026 input6/a_27_47# net15 0.00115f
C1027 _35_/a_489_413# _08_ 5.56e-19
C1028 _04_ _17_ 4.34e-19
C1029 _15_ _50_/a_223_47# 0.00698f
C1030 net4 _53_/a_29_53# 3.26e-19
C1031 p[8] _37_/a_27_47# 9.82e-21
C1032 _10_ _52_/a_93_21# 0.00534f
C1033 _45_/a_109_297# _02_ 8.44e-19
C1034 _06_ p[6] 2.62e-19
C1035 _27_/a_27_297# input5/a_664_47# 0.0116f
C1036 _34_/a_47_47# _25_ 1.08e-19
C1037 _43_/a_297_47# _17_ 5.72e-20
C1038 _10_ net8 5.86e-19
C1039 _14_ _12_ 1.98e-20
C1040 _35_/a_226_47# p[7] 2.82e-19
C1041 _48_/a_27_47# net10 8.4e-21
C1042 _26_/a_29_53# net14 1.33e-20
C1043 _38_/a_27_47# _06_ 0.0172f
C1044 VPWR p[10] 0.177f
C1045 _06_ _42_/a_209_311# 1.66e-19
C1046 _22_ _30_/a_215_297# 2.46e-21
C1047 input2/a_27_47# _15_ 3.18e-20
C1048 _38_/a_109_47# _12_ 0.00179f
C1049 p[3] net8 0.0015f
C1050 _00_ _26_/a_111_297# 3.7e-19
C1051 net2 _15_ 9.8e-19
C1052 _18_ net3 7.34e-20
C1053 _06_ b[3] 9.96e-21
C1054 _50_/a_27_47# _11_ 0.0592f
C1055 _27_/a_27_297# _27_/a_109_297# -3.68e-20
C1056 net6 input15/a_27_47# 0.146f
C1057 VPWR _35_/a_76_199# -0.00947f
C1058 _40_/a_109_297# _20_ 2.35e-20
C1059 net1 _02_ 0.00251f
C1060 net14 net7 2.23e-19
C1061 net1 _03_ 0.298f
C1062 net1 input8/a_27_47# 0.0347f
C1063 b[2] _52_/a_93_21# 1.63e-19
C1064 p[5] net12 0.00294f
C1065 _35_/a_489_413# _09_ 0.0296f
C1066 net5 _06_ 0.41f
C1067 p[10] net15 0.01f
C1068 input8/a_27_47# input7/a_27_47# 3.2e-20
C1069 net10 input12/a_27_47# 0.00182f
C1070 _21_ p[6] 0.00203f
C1071 _42_/a_209_311# _18_ 3.21e-19
C1072 net12 _11_ 3.82e-21
C1073 _21_ _38_/a_27_47# 3.87e-19
C1074 input4/a_75_212# _39_/a_47_47# 3.1e-19
C1075 _26_/a_183_297# _15_ 4.63e-36
C1076 p[2] _01_ 0.00164f
C1077 _27_/a_27_297# _16_ 3.74e-22
C1078 _06_ _52_/a_584_47# 0.00218f
C1079 _35_/a_489_413# net13 7.36e-20
C1080 p[8] net6 5.98e-19
C1081 net6 _30_/a_215_297# 3.3e-21
C1082 _34_/a_129_47# _08_ 3.29e-19
C1083 _45_/a_109_297# _17_ 4.29e-22
C1084 _26_/a_29_53# net9 0.00343f
C1085 VPWR _45_/a_193_297# -0.00859f
C1086 net5 _50_/a_343_93# 0.00124f
C1087 net5 _18_ 0.0426f
C1088 _05_ _33_/a_368_53# 9.2e-19
C1089 _21_ net5 0.00784f
C1090 _03_ _34_/a_377_297# 3.13e-20
C1091 _25_ net18 0.0594f
C1092 VPWR net14 0.182f
C1093 _06_ _50_/a_223_47# 0.0481f
C1094 input5/a_62_47# p[0] 1.39e-19
C1095 _06_ _05_ 0.00724f
C1096 _44_/a_250_297# _17_ 0.0336f
C1097 net5 _24_ 5.83e-20
C1098 _47_/a_299_297# _20_ 0.002f
C1099 _39_/a_47_47# net4 0.0202f
C1100 _10_ _32_/a_27_47# 0.00217f
C1101 _30_/a_215_297# net13 0.0246f
C1102 _16_ _43_/a_27_47# 2.47e-19
C1103 net4 _52_/a_93_21# 7.93e-20
C1104 _26_/a_29_53# _22_ 0.09f
C1105 _48_/a_181_47# _07_ 5.93e-19
C1106 net9 net7 0.00233f
C1107 net19 _44_/a_346_47# 0.00124f
C1108 net1 input12/a_27_47# 7.44e-20
C1109 input5/a_841_47# _02_ 0.00591f
C1110 _38_/a_27_47# _50_/a_27_47# 2.37e-20
C1111 _45_/a_27_47# _23_ 1.74e-19
C1112 input5/a_558_47# _04_ 1.25e-20
C1113 _33_/a_109_93# _12_ 9.75e-20
C1114 net2 _06_ 0.0108f
C1115 _00_ _11_ 0.238f
C1116 input14/a_27_47# net14 0.0232f
C1117 _55_/a_217_297# net14 2.1e-19
C1118 _55_/a_80_21# _01_ 0.0121f
C1119 net14 net15 1.07f
C1120 _50_/a_223_47# _18_ 0.0367f
C1121 net12 p[6] 0.0255f
C1122 net17 net3 3.72e-19
C1123 _21_ _50_/a_223_47# 2.91e-21
C1124 _22_ net7 2.73e-20
C1125 _21_ _05_ 0.0104f
C1126 _06_ _52_/a_256_47# 0.00157f
C1127 _27_/a_27_297# _04_ 0.0526f
C1128 _31_/a_35_297# _49_/a_201_297# 5.52e-20
C1129 _16_ _20_ 0.00271f
C1130 net5 _50_/a_27_47# 0.0169f
C1131 _10_ net11 0.0109f
C1132 net19 _15_ 0.166f
C1133 output16/a_27_47# net6 1.5e-19
C1134 _08_ net7 9.54e-25
C1135 _43_/a_193_413# _20_ 0.00161f
C1136 _22_ _41_/a_59_75# 6.24e-22
C1137 _33_/a_109_93# _52_/a_250_297# 5.17e-22
C1138 _43_/a_469_47# net14 1.44e-20
C1139 _14_ _44_/a_256_47# 0.00124f
C1140 _28_/a_109_297# net9 3.7e-19
C1141 net2 _50_/a_343_93# 1.25e-20
C1142 _26_/a_183_297# _06_ 3.16e-19
C1143 net2 _18_ 0.00181f
C1144 p[12] _12_ 2.08e-20
C1145 net17 _42_/a_209_311# 1.04e-21
C1146 _36_/a_27_47# _02_ 9.37e-20
C1147 VPWR net9 0.5f
C1148 _14_ _11_ 0.0415f
C1149 _07_ _34_/a_285_47# 0.00975f
C1150 b[1] p[10] 0.286f
C1151 _29_/a_29_53# _06_ 0.00111f
C1152 net5 net12 0.0674f
C1153 _37_/a_27_47# VPWR -0.0178f
C1154 _26_/a_29_53# net6 0.0032f
C1155 p[2] _02_ 7.08e-19
C1156 p[2] input8/a_27_47# 0.0159f
C1157 _10_ _55_/a_472_297# 7.35e-21
C1158 _00_ net3 2.12e-19
C1159 net11 b[2] 1.46e-19
C1160 VPWR _22_ 1.4f
C1161 _22_ _53_/a_183_297# 3.71e-20
C1162 p[12] _52_/a_250_297# 1.84e-20
C1163 net9 net15 8.49e-20
C1164 net5 net17 4.21e-21
C1165 _26_/a_29_53# net13 2.23e-20
C1166 _09_ net7 0.00258f
C1167 _50_/a_27_47# _50_/a_223_47# 5.68e-32
C1168 output18/a_27_47# net18 0.0106f
C1169 VPWR _08_ -0.0171f
C1170 VPWR _38_/a_303_47# -4.83e-19
C1171 net19 _42_/a_296_53# 2.71e-19
C1172 _40_/a_297_297# _20_ 9.18e-21
C1173 _39_/a_285_47# net6 1.53e-19
C1174 _02_ _53_/a_111_297# 9.57e-20
C1175 output16/a_27_47# _13_ 4.58e-19
C1176 _37_/a_27_47# net15 0.0541f
C1177 p[10] _19_ 0.00226f
C1178 p[10] net8 0.0097f
C1179 _44_/a_250_297# output19/a_27_47# 6.42e-20
C1180 input12/a_27_47# p[4] 8.26e-19
C1181 _27_/a_205_297# net14 3.63e-19
C1182 _21_ _29_/a_29_53# 0.0775f
C1183 _00_ b[3] 1.04e-19
C1184 _04_ _20_ 0.0677f
C1185 _41_/a_59_75# net6 0.0373f
C1186 _05_ net12 0.0414f
C1187 _52_/a_93_21# _35_/a_76_199# 6.83e-21
C1188 b[3] _44_/a_584_47# 0.00109f
C1189 _22_ net15 2.74e-19
C1190 _14_ net3 0.0295f
C1191 net7 net13 1.72e-19
C1192 _14_ _55_/a_300_47# 8.09e-19
C1193 _10_ _44_/a_93_21# 2.48e-19
C1194 _39_/a_129_47# _17_ 1.38e-20
C1195 net10 _25_ 2.02e-19
C1196 net16 _25_ 1.16e-19
C1197 _36_/a_109_47# net13 0.00126f
C1198 _30_/a_392_297# net12 2.19e-20
C1199 input5/a_558_47# net1 1.1e-19
C1200 _55_/a_80_21# _02_ 0.164f
C1201 _00_ net5 0.00954f
C1202 net17 _05_ 0.0111f
C1203 _29_/a_111_297# VPWR -5.85e-19
C1204 net19 _06_ 0.00522f
C1205 input5/a_558_47# input7/a_27_47# 1.22e-20
C1206 _14_ _42_/a_209_311# 0.00142f
C1207 _15_ _42_/a_296_53# 1.28e-19
C1208 VPWR _09_ 0.297f
C1209 _09_ _53_/a_183_297# 4.18e-19
C1210 input12/a_27_47# p[7] 3.2e-20
C1211 net3 _49_/a_75_199# 2.01e-19
C1212 net1 _47_/a_81_21# 1.58e-21
C1213 VPWR net6 0.999f
C1214 _14_ b[3] 1.92e-19
C1215 _27_/a_27_297# net1 6.05e-21
C1216 _22_ _53_/a_29_53# 0.00749f
C1217 _39_/a_47_47# _45_/a_193_297# 1.4e-20
C1218 input2/a_27_47# net17 0.0398f
C1219 p[10] output17/a_27_47# 0.118f
C1220 _39_/a_285_47# _13_ 0.00451f
C1221 net2 net17 0.261f
C1222 _29_/a_29_53# _50_/a_27_47# 1.44e-20
C1223 _52_/a_93_21# _45_/a_193_297# 6.01e-19
C1224 p[8] p[11] 0.0023f
C1225 _27_/a_27_297# input7/a_27_47# 0.00119f
C1226 _42_/a_368_53# net3 3.82e-19
C1227 VPWR net13 0.599f
C1228 net19 _18_ 4.89e-20
C1229 net10 _20_ 3.23e-19
C1230 net5 _14_ 3.89e-19
C1231 net14 net8 0.0516f
C1232 net11 _07_ 0.0206f
C1233 net14 _19_ 0.0512f
C1234 _00_ _50_/a_223_47# 0.00738f
C1235 _06_ _15_ 0.22f
C1236 net6 net15 0.0664f
C1237 _00_ _05_ 5.03e-22
C1238 _29_/a_29_53# net12 0.0132f
C1239 _10_ _12_ 0.19f
C1240 VPWR _33_/a_296_53# -1.15e-19
C1241 net11 _33_/a_209_311# 2.49e-19
C1242 _10_ _30_/a_297_297# 1.25e-20
C1243 input5/a_62_47# _04_ 0.00345f
C1244 net15 net13 8.84e-19
C1245 input5/a_558_47# input5/a_841_47# -4.44e-34
C1246 _43_/a_469_47# net6 4.85e-21
C1247 p[12] _11_ 3.51e-21
C1248 _35_/a_226_47# net7 2.93e-20
C1249 _55_/a_80_21# _17_ 7.64e-21
C1250 _00_ net2 0.00732f
C1251 VPWR _13_ 0.0804f
C1252 _31_/a_35_297# net17 0.0514f
C1253 net2 _44_/a_584_47# 0.0053f
C1254 p[14] input15/a_27_47# 6.15e-19
C1255 _36_/a_303_47# net11 7.63e-20
C1256 net9 _30_/a_109_53# 0.0193f
C1257 _10_ _39_/a_377_297# 7.42e-19
C1258 VPWR _50_/a_615_93# -5.34e-19
C1259 _09_ _53_/a_29_53# 0.00642f
C1260 input1/a_75_212# p[0] 0.0172f
C1261 _15_ _50_/a_343_93# 0.0098f
C1262 _15_ _18_ 0.042f
C1263 net6 _53_/a_29_53# 2.11e-20
C1264 _10_ _52_/a_250_297# 0.00368f
C1265 _35_/a_489_413# _02_ 3.86e-19
C1266 _21_ _15_ 1.13e-21
C1267 _03_ _35_/a_489_413# 0.0205f
C1268 net1 _20_ 0.363f
C1269 net16 output18/a_27_47# 3.45e-19
C1270 _43_/a_369_47# _17_ 5.87e-19
C1271 b[2] _12_ 3.89e-20
C1272 _49_/a_208_47# _09_ 5.43e-21
C1273 _22_ _30_/a_109_53# 3.67e-21
C1274 input5/a_381_47# net7 4.91e-19
C1275 _10_ _26_/a_111_297# 7.13e-20
C1276 _38_/a_197_47# _12_ 0.00173f
C1277 _00_ _26_/a_183_297# 4.53e-19
C1278 net9 net8 0.0605f
C1279 net2 _14_ 0.0104f
C1280 input4/a_75_212# _12_ 2.09e-20
C1281 net11 _35_/a_76_199# 4e-19
C1282 _30_/a_215_297# _02_ 3.58e-21
C1283 VPWR _35_/a_226_47# 0.00159f
C1284 input3/a_27_47# net14 3.47e-19
C1285 p[8] p[14] 0.226f
C1286 _37_/a_27_47# net8 6.66e-21
C1287 _03_ _30_/a_215_297# 0.0393f
C1288 input6/a_27_47# _44_/a_93_21# 8.53e-19
C1289 _01_ net7 0.233f
C1290 b[2] _52_/a_250_297# 1.6e-19
C1291 _22_ _52_/a_93_21# 0.0347f
C1292 _35_/a_226_297# _09_ 4.98e-19
C1293 _22_ net8 3.3e-20
C1294 _06_ _33_/a_368_53# 1.7e-19
C1295 b[0] b[2] 0.183f
C1296 net19 net17 8.84e-23
C1297 _50_/a_27_47# _15_ 5.65e-19
C1298 _13_ _53_/a_29_53# 9.05e-19
C1299 _17_ input15/a_27_47# 6.14e-19
C1300 _26_/a_183_297# _14_ 6.98e-22
C1301 input5/a_381_47# VPWR 8.33e-19
C1302 net16 _45_/a_27_47# 8.68e-19
C1303 input12/a_27_47# input10/a_27_47# 0.0154f
C1304 input5/a_62_47# _44_/a_250_297# 2.45e-20
C1305 net4 _12_ 0.105f
C1306 _35_/a_226_297# net13 6.88e-19
C1307 p[10] _42_/a_109_93# 1.82e-21
C1308 p[12] b[3] 7.54e-20
C1309 _07_ _35_/a_556_47# 0.00128f
C1310 _34_/a_285_47# _08_ 0.00414f
C1311 VPWR _45_/a_205_47# -1.62e-19
C1312 _36_/a_197_47# net5 0.00254f
C1313 _36_/a_27_47# _25_ 2.34e-20
C1314 net10 input13/a_27_47# 8.86e-20
C1315 _04_ _34_/a_47_47# 1.17e-20
C1316 net10 _23_ 7.53e-19
C1317 net11 net14 9.95e-19
C1318 VPWR _01_ 0.521f
C1319 _06_ _50_/a_343_93# 0.0376f
C1320 _06_ _18_ 0.54f
C1321 _39_/a_47_47# _09_ 7.7e-21
C1322 input5/a_62_47# net1 7.59e-20
C1323 _21_ _06_ 0.143f
C1324 _09_ _52_/a_93_21# 0.0227f
C1325 net5 p[12] 4.79e-20
C1326 _39_/a_377_297# net4 8.88e-19
C1327 _39_/a_47_47# net6 0.0249f
C1328 input5/a_381_47# net15 7.15e-19
C1329 _30_/a_109_53# net13 1.05e-19
C1330 _29_/a_29_53# _49_/a_75_199# 1.28e-19
C1331 _07_ _12_ 2.94e-23
C1332 _06_ _24_ 0.113f
C1333 p[13] p[10] 0.124f
C1334 _31_/a_35_297# _49_/a_75_199# 6.24e-19
C1335 _16_ _43_/a_193_413# 0.0261f
C1336 net4 _52_/a_250_297# 0.00136f
C1337 net6 _52_/a_93_21# 2.33e-19
C1338 _33_/a_109_93# _05_ 0.0206f
C1339 _09_ _19_ 4.8e-21
C1340 input5/a_664_47# _04_ 6.73e-21
C1341 b[0] net4 0.0024f
C1342 VPWR p[11] 0.247f
C1343 _32_/a_27_47# net9 0.0136f
C1344 _33_/a_209_311# _12_ 2.88e-20
C1345 _10_ _11_ 0.176f
C1346 _39_/a_129_47# _20_ 1.71e-20
C1347 _26_/a_29_53# _02_ 0.0466f
C1348 _01_ net15 0.0314f
C1349 input3/a_27_47# _22_ 5.13e-20
C1350 _26_/a_29_53# _03_ 7.93e-21
C1351 _10_ input9/a_75_212# 5.49e-21
C1352 _55_/a_217_297# _01_ 0.00112f
C1353 _52_/a_93_21# net13 7.21e-19
C1354 _50_/a_343_93# _18_ 0.0276f
C1355 _36_/a_27_47# _20_ 0.00148f
C1356 net8 net13 7.51e-20
C1357 p[9] _11_ 1.01e-19
C1358 _19_ net13 4.45e-20
C1359 input9/a_75_212# p[3] 0.0157f
C1360 _27_/a_109_297# _04_ 7.2e-20
C1361 _32_/a_27_47# _22_ 1.76e-19
C1362 input14/a_27_47# p[11] 0.00118f
C1363 _21_ _24_ 0.0388f
C1364 net19 _14_ 0.00714f
C1365 net1 input13/a_27_47# 1.9e-19
C1366 net10 _34_/a_47_47# 0.0507f
C1367 p[11] net15 3.83e-19
C1368 _02_ net7 0.445f
C1369 _00_ _15_ 0.207f
C1370 _49_/a_315_47# _04_ 7.71e-19
C1371 input8/a_27_47# net7 1.47e-19
C1372 _14_ _44_/a_346_47# 3.76e-19
C1373 _39_/a_285_47# _02_ 0.0019f
C1374 _42_/a_109_93# net14 0.00351f
C1375 _06_ _50_/a_27_47# 0.00972f
C1376 _34_/a_285_47# net13 4.11e-20
C1377 _03_ net7 0.078f
C1378 p[0] net1 0.00473f
C1379 net9 net11 0.136f
C1380 _39_/a_47_47# _13_ 0.00117f
C1381 _52_/a_93_21# _13_ 1.31e-19
C1382 net12 _33_/a_368_53# 2.63e-19
C1383 _43_/a_27_47# _55_/a_80_21# 1.56e-19
C1384 net14 _44_/a_93_21# 0.0646f
C1385 p[14] _41_/a_59_75# 5.13e-20
C1386 _37_/a_109_47# VPWR -4.38e-19
C1387 p[0] input7/a_27_47# 5.13e-20
C1388 _06_ net12 0.284f
C1389 _10_ net3 3.89e-19
C1390 _32_/a_303_47# net5 7.18e-21
C1391 p[13] net14 1.91e-19
C1392 net11 _22_ 6.82e-21
C1393 _04_ _43_/a_193_413# 5.67e-21
C1394 _35_/a_76_199# _12_ 6.84e-20
C1395 _01_ _49_/a_208_47# 2.13e-19
C1396 p[10] p[1] 9.52e-20
C1397 _50_/a_27_47# _18_ 0.0665f
C1398 _15_ _14_ 0.148f
C1399 net3 p[9] 1.63e-19
C1400 net11 _08_ 8.83e-19
C1401 _21_ _50_/a_27_47# 3.38e-21
C1402 net19 _42_/a_368_53# 5.12e-19
C1403 VPWR _02_ 0.33f
C1404 _10_ _38_/a_27_47# 0.0133f
C1405 VPWR input8/a_27_47# 0.0863f
C1406 _55_/a_80_21# _20_ 0.0291f
C1407 VPWR _03_ 0.845f
C1408 _02_ _53_/a_183_297# 4.14e-19
C1409 VPWR p[14] 0.0416f
C1410 _31_/a_285_297# _05_ 6.12e-19
C1411 _27_/a_277_297# net14 5.1e-19
C1412 _18_ net12 2.25e-21
C1413 _10_ b[3] 3.27e-20
C1414 _52_/a_250_297# _35_/a_76_199# 3.4e-21
C1415 _21_ net12 0.23f
C1416 _52_/a_93_21# _35_/a_226_47# 4.89e-20
C1417 _42_/a_209_311# p[9] 5.51e-21
C1418 p[8] output19/a_27_47# 0.0218f
C1419 net4 _11_ 0.0858f
C1420 _39_/a_285_47# _17_ 7.36e-21
C1421 _37_/a_27_47# _42_/a_109_93# 2.55e-20
C1422 b[3] p[9] 0.0898f
C1423 net16 net18 0.00585f
C1424 _48_/a_27_47# VPWR 0.0158f
C1425 input5/a_664_47# net1 2.41e-19
C1426 _12_ _45_/a_193_297# 0.0103f
C1427 _02_ net15 0.0806f
C1428 _03_ net15 4.26e-20
C1429 _55_/a_217_297# _02_ 6.01e-19
C1430 _10_ net5 0.199f
C1431 p[14] net15 0.00132f
C1432 _41_/a_59_75# _17_ 0.00149f
C1433 input5/a_664_47# input7/a_27_47# 1.08e-21
C1434 _29_/a_111_297# net11 8.27e-19
C1435 _29_/a_183_297# VPWR -8.13e-19
C1436 p[4] input13/a_27_47# 7.37e-20
C1437 _30_/a_465_297# net10 0.00106f
C1438 net11 _09_ 0.0262f
C1439 _37_/a_27_47# _44_/a_93_21# 3.19e-19
C1440 _22_ _42_/a_109_93# 1.21e-19
C1441 _00_ _06_ 0.1f
C1442 _25_ input10/a_27_47# 2.03e-20
C1443 net11 net6 1.08e-19
C1444 _14_ _49_/a_201_297# 4.76e-21
C1445 p[13] net9 1.72e-19
C1446 input5/a_381_47# net8 7.48e-19
C1447 net14 p[1] 0.0025f
C1448 _16_ _44_/a_250_297# 3.25e-19
C1449 b[1] p[11] 1.84e-20
C1450 _36_/a_27_47# _23_ 0.00118f
C1451 VPWR input12/a_27_47# 0.0646f
C1452 net11 net13 0.093f
C1453 _02_ _53_/a_29_53# 0.0388f
C1454 _50_/a_27_47# net12 7.99e-21
C1455 net5 b[2] 7.33e-20
C1456 VPWR _17_ 0.306f
C1457 _01_ net8 0.0802f
C1458 _00_ _50_/a_343_93# 0.102f
C1459 _00_ _18_ 0.157f
C1460 _10_ _50_/a_223_47# 0.0295f
C1461 _10_ _05_ 9.25e-21
C1462 net4 net3 9.28e-21
C1463 _01_ _19_ 0.031f
C1464 _06_ _14_ 0.0556f
C1465 _21_ _00_ 9.26e-20
C1466 p[7] input13/a_27_47# 0.0167f
C1467 _49_/a_208_47# _02_ 0.00193f
C1468 p[12] net19 6.8e-20
C1469 _03_ _49_/a_208_47# 3.86e-19
C1470 p[3] _05_ 5.83e-21
C1471 net5 input4/a_75_212# 0.0104f
C1472 _48_/a_27_47# _53_/a_29_53# 3.14e-21
C1473 net10 _04_ 0.121f
C1474 net11 _13_ 2.34e-19
C1475 net9 _12_ 4.39e-22
C1476 _10_ net2 2.65e-19
C1477 _17_ net15 0.195f
C1478 _38_/a_27_47# net4 0.0119f
C1479 _31_/a_117_297# net17 0.00149f
C1480 input5/a_381_47# output17/a_27_47# 6.6e-20
C1481 net9 _30_/a_297_297# 7.83e-19
C1482 input6/a_27_47# net3 2.52e-19
C1483 net17 net12 2.11e-21
C1484 input1/a_75_212# net1 0.00208f
C1485 _27_/a_205_297# _03_ 1.46e-20
C1486 _14_ _50_/a_343_93# 9.76e-19
C1487 _14_ _18_ 0.243f
C1488 _15_ _50_/a_429_93# 6.82e-19
C1489 _30_/a_215_297# _20_ 6.08e-19
C1490 _35_/a_556_47# _08_ 7.71e-19
C1491 _10_ _52_/a_256_47# 1.65e-19
C1492 net2 p[9] 0.00112f
C1493 net6 _44_/a_93_21# 1.08e-20
C1494 input1/a_75_212# input7/a_27_47# 3.2e-20
C1495 _03_ _35_/a_226_297# 0.00101f
C1496 _22_ _12_ 0.196f
C1497 _35_/a_76_199# _11_ 6.99e-22
C1498 _07_ p[6] 1.26e-19
C1499 _43_/a_469_47# _17_ 0.00177f
C1500 p[12] _15_ 0.0162f
C1501 net5 net4 0.0447f
C1502 input5/a_558_47# net7 0.00358f
C1503 _00_ _50_/a_27_47# 0.00197f
C1504 _38_/a_303_47# _12_ 0.00153f
C1505 _04_ _44_/a_250_297# 5.57e-21
C1506 _10_ _26_/a_183_297# 5.74e-19
C1507 _30_/a_109_53# _02_ 5.03e-22
C1508 b[1] _03_ 0.00143f
C1509 _48_/a_181_47# _02_ 3.9e-19
C1510 _10_ _29_/a_29_53# 5.17e-19
C1511 input6/a_27_47# b[3] 4.02e-19
C1512 _21_ _49_/a_75_199# 6.64e-19
C1513 net11 _35_/a_226_47# 3.21e-19
C1514 _03_ _30_/a_109_53# 0.0189f
C1515 _16_ input5/a_841_47# 8.62e-19
C1516 net1 _04_ 0.018f
C1517 _22_ _52_/a_250_297# 0.099f
C1518 _27_/a_27_297# net7 1.22e-19
C1519 _35_/a_556_47# _09_ 3.74e-19
C1520 p[10] net3 7.98e-19
C1521 _29_/a_29_53# p[3] 2.07e-19
C1522 _32_/a_27_47# _01_ 0.0266f
C1523 _47_/a_81_21# _41_/a_59_75# 1.5e-19
C1524 _39_/a_47_47# _02_ 0.0127f
C1525 _03_ _39_/a_47_47# 1.47e-19
C1526 input3/a_27_47# p[11] 0.0157f
C1527 _52_/a_93_21# _02_ 0.0957f
C1528 _44_/a_256_47# net14 0.00379f
C1529 _45_/a_193_297# _11_ 0.0292f
C1530 _03_ _52_/a_93_21# 0.00985f
C1531 _50_/a_223_47# net4 0.0107f
C1532 _26_/a_111_297# _22_ 0.00137f
C1533 net8 _02_ 0.334f
C1534 input8/a_27_47# net8 0.0181f
C1535 _02_ _19_ 0.213f
C1536 _03_ net8 0.0287f
C1537 _09_ _12_ 0.00509f
C1538 VPWR output19/a_27_47# 0.0229f
C1539 net14 _11_ 5e-19
C1540 _03_ _19_ 0.0019f
C1541 _06_ _33_/a_109_93# 9.13e-19
C1542 input5/a_558_47# VPWR 0.0083f
C1543 net16 _45_/a_109_297# 5.1e-20
C1544 net6 _12_ 0.0891f
C1545 p[10] _42_/a_209_311# 2.37e-20
C1546 _49_/a_315_47# p[2] 6.65e-20
C1547 p[10] b[3] 3.13e-20
C1548 _34_/a_285_47# _02_ 7.14e-19
C1549 _36_/a_303_47# net5 0.00256f
C1550 VPWR _45_/a_465_47# -5.05e-19
C1551 p[8] input5/a_62_47# 1.15e-19
C1552 _04_ _34_/a_377_297# 1.7e-20
C1553 _43_/a_27_47# net7 6.31e-19
C1554 _36_/a_109_47# _25_ 3.76e-21
C1555 VPWR _47_/a_81_21# 0.00889f
C1556 net11 _01_ 3.82e-20
C1557 _26_/a_29_53# _20_ 0.00447f
C1558 _36_/a_197_47# _06_ 6.18e-19
C1559 _06_ _50_/a_429_93# 0.00169f
C1560 _45_/a_27_47# _35_/a_489_413# 3.89e-21
C1561 _07_ _05_ 1.21e-19
C1562 _12_ net13 0.00632f
C1563 input14/a_27_47# output19/a_27_47# 0.0101f
C1564 _27_/a_27_297# VPWR 0.0329f
C1565 output19/a_27_47# net15 6.88e-19
C1566 _39_/a_377_297# net6 0.00143f
C1567 VPWR _47_/a_384_47# -1.45e-19
C1568 net1 net10 0.00388f
C1569 input5/a_558_47# net15 0.00672f
C1570 _09_ _52_/a_250_297# 1.97e-20
C1571 _30_/a_297_297# net13 3.27e-20
C1572 _14_ net17 2.4e-20
C1573 _10_ net19 0.00224f
C1574 net5 p[10] 5.12e-21
C1575 p[12] _06_ 0.0535f
C1576 net6 _52_/a_250_297# 0.00133f
C1577 _21_ _33_/a_109_93# 1.62e-20
C1578 _33_/a_209_311# _05_ 0.0311f
C1579 _10_ _44_/a_346_47# 9.13e-21
C1580 b[0] net6 2.52e-19
C1581 _48_/a_27_47# _34_/a_285_47# 6.66e-20
C1582 net7 _20_ 0.0257f
C1583 _32_/a_109_47# net9 6.44e-19
C1584 net19 p[9] 0.0729f
C1585 output16/a_27_47# output18/a_27_47# 7.85e-19
C1586 _47_/a_81_21# net15 0.00106f
C1587 _55_/a_472_297# _01_ 6.28e-19
C1588 _03_ output17/a_27_47# 1.95e-19
C1589 _39_/a_47_47# _17_ 1.47e-20
C1590 net5 _35_/a_76_199# 3.38e-19
C1591 VPWR _25_ 0.0829f
C1592 net14 net3 0.689f
C1593 _27_/a_27_297# net15 0.00888f
C1594 input5/a_381_47# _42_/a_109_93# 0.00763f
C1595 _26_/a_111_297# net6 1.12e-19
C1596 net2 input6/a_27_47# 0.0047f
C1597 _41_/a_59_75# _20_ 1.78e-20
C1598 _12_ _13_ 0.462f
C1599 net17 _49_/a_75_199# 0.00127f
C1600 net9 _11_ 5.39e-19
C1601 VPWR _43_/a_27_47# 0.0186f
C1602 input9/a_75_212# net9 0.0247f
C1603 _17_ net8 4.52e-20
C1604 _17_ _19_ 8.82e-21
C1605 p[12] _18_ 3.95e-21
C1606 _37_/a_27_47# _11_ 0.0018f
C1607 _10_ _15_ 0.479f
C1608 net10 _34_/a_377_297# 1.62e-19
C1609 _00_ _14_ 0.133f
C1610 _42_/a_209_311# net14 0.0238f
C1611 _01_ _31_/a_285_47# 3.36e-19
C1612 p[10] _05_ 6e-20
C1613 _32_/a_27_47# _02_ 0.00247f
C1614 input5/a_381_47# p[13] 0.00153f
C1615 _22_ _11_ 0.15f
C1616 b[3] net14 0.0172f
C1617 _04_ _36_/a_27_47# 0.00169f
C1618 _32_/a_27_47# _03_ 1.9e-19
C1619 _16_ _55_/a_80_21# 0.0143f
C1620 _28_/a_109_297# _20_ 0.00221f
C1621 _15_ p[9] 2.06e-19
C1622 _29_/a_29_53# _07_ 1.19e-20
C1623 _52_/a_250_297# _13_ 5.43e-19
C1624 _31_/a_285_297# _06_ 1.01e-20
C1625 net1 input7/a_27_47# 0.0383f
C1626 _43_/a_193_413# _55_/a_80_21# 2.54e-19
C1627 _43_/a_27_47# _55_/a_217_297# 2.18e-19
C1628 _37_/a_197_47# VPWR -3.27e-19
C1629 VPWR _20_ 0.342f
C1630 _05_ _35_/a_76_199# 0.00238f
C1631 p[11] _42_/a_109_93# 4.55e-21
C1632 b[0] _13_ 0.00299f
C1633 net5 _45_/a_193_297# 0.00935f
C1634 p[2] _04_ 1.83e-20
C1635 input2/a_27_47# p[10] 0.00924f
C1636 net2 p[10] 0.0632f
C1637 _35_/a_226_47# _12_ 8.38e-20
C1638 _04_ p[7] 0.00142f
C1639 p[13] _01_ 2.02e-20
C1640 net5 net14 0.0263f
C1641 net9 net3 5.09e-20
C1642 _33_/a_109_93# net12 0.0435f
C1643 VPWR _40_/a_191_297# -6.82e-19
C1644 _43_/a_369_47# _43_/a_193_413# -1.25e-19
C1645 net11 _02_ 0.0327f
C1646 _25_ _53_/a_29_53# 0.00146f
C1647 net10 p[4] 0.00268f
C1648 _37_/a_197_47# net15 1.78e-19
C1649 _55_/a_217_297# _20_ 0.0013f
C1650 _37_/a_27_47# net3 0.094f
C1651 net15 _20_ 0.0021f
C1652 input5/a_62_47# net7 2.04e-19
C1653 p[13] p[11] 0.00897f
C1654 _03_ net11 0.0952f
C1655 p[12] _50_/a_27_47# 1.34e-19
C1656 net19 net4 2.65e-20
C1657 _36_/a_197_47# net12 4.67e-20
C1658 _52_/a_250_297# _35_/a_226_47# 2.63e-20
C1659 _22_ net3 9.39e-20
C1660 _22_ _55_/a_300_47# 2.08e-19
C1661 _09_ _11_ 0.0665f
C1662 _05_ _45_/a_193_297# 4.84e-22
C1663 _14_ _49_/a_75_199# 6.79e-20
C1664 _40_/a_191_297# net15 8.41e-19
C1665 net10 _36_/a_27_47# 0.0366f
C1666 VPWR output18/a_27_47# 0.0689f
C1667 net6 _11_ 0.0257f
C1668 _48_/a_27_47# net11 0.0179f
C1669 _50_/a_223_47# net14 5.89e-21
C1670 _37_/a_27_47# _42_/a_209_311# 1.59e-20
C1671 _31_/a_35_297# p[10] 2.29e-19
C1672 input5/a_841_47# net1 1.33e-19
C1673 _55_/a_472_297# _02_ 1.25e-19
C1674 _12_ _45_/a_205_47# 7.46e-19
C1675 _16_ input15/a_27_47# 7.13e-19
C1676 p[5] net13 1.05e-19
C1677 _29_/a_183_297# net11 3.64e-19
C1678 net10 p[7] 4.96e-19
C1679 _22_ _42_/a_209_311# 1.72e-19
C1680 _38_/a_27_47# _22_ 2.86e-19
C1681 _43_/a_193_413# input15/a_27_47# 1.62e-20
C1682 _10_ _06_ 1.14f
C1683 _29_/a_29_53# _35_/a_76_199# 9.88e-19
C1684 net18 input10/a_27_47# 4.16e-20
C1685 net19 input6/a_27_47# 0.00586f
C1686 input9/a_75_212# net13 4.4e-19
C1687 net5 net9 0.0368f
C1688 _08_ p[6] 1.55e-19
C1689 input2/a_27_47# net14 0.0102f
C1690 _22_ b[3] 1.28e-19
C1691 _15_ net4 0.00427f
C1692 input5/a_558_47# net8 0.00357f
C1693 input5/a_62_47# VPWR 0.0601f
C1694 net2 net14 0.151f
C1695 _06_ p[9] 0.00205f
C1696 p[3] _06_ 1.59e-20
C1697 _39_/a_285_47# _23_ 1.9e-20
C1698 _37_/a_27_47# net5 1.13e-20
C1699 _03_ _31_/a_285_47# 8.54e-19
C1700 p[0] net7 1.36e-19
C1701 net11 input12/a_27_47# 0.00246f
C1702 _36_/a_109_47# _23_ 3.44e-19
C1703 net5 _22_ 0.405f
C1704 _47_/a_81_21# net8 2.08e-21
C1705 net1 _36_/a_27_47# 6.99e-20
C1706 p[14] _44_/a_93_21# 2.82e-20
C1707 net6 net3 0.00152f
C1708 _10_ _18_ 0.133f
C1709 _10_ _50_/a_343_93# 0.0284f
C1710 _27_/a_27_297# net8 0.0108f
C1711 _10_ _21_ 0.00421f
C1712 _06_ b[2] 0.0116f
C1713 _13_ _11_ 0.164f
C1714 _27_/a_27_297# _19_ 0.082f
C1715 _45_/a_27_47# VPWR -0.00418f
C1716 p[13] _02_ 7.58e-20
C1717 _15_ input6/a_27_47# 5.75e-19
C1718 _10_ _24_ 0.00484f
C1719 p[2] net1 0.0269f
C1720 _22_ _52_/a_584_47# 6.24e-19
C1721 _06_ _38_/a_197_47# 4.32e-19
C1722 net9 _05_ 0.124f
C1723 net9 _50_/a_223_47# 2e-19
C1724 output18/a_27_47# _53_/a_29_53# 9.46e-19
C1725 _21_ p[3] 3.95e-21
C1726 net1 p[7] 7.5e-20
C1727 p[10] net19 1.26e-21
C1728 _38_/a_27_47# _09_ 0.00195f
C1729 _29_/a_29_53# net14 1.61e-20
C1730 net3 net13 3.25e-21
C1731 p[2] input7/a_27_47# 0.0023f
C1732 VPWR input13/a_27_47# 0.0696f
C1733 _42_/a_209_311# net6 1.32e-20
C1734 VPWR _23_ -0.00374f
C1735 input4/a_75_212# _06_ 0.00205f
C1736 _52_/a_346_47# _02_ 0.00526f
C1737 net9 _30_/a_392_297# 9.92e-19
C1738 b[3] net6 7.68e-19
C1739 VPWR p[0] 0.0836f
C1740 _27_/a_277_297# _03_ 2.1e-20
C1741 _15_ _50_/a_515_93# 0.00147f
C1742 _22_ _50_/a_223_47# 0.031f
C1743 net2 net9 3.64e-20
C1744 _30_/a_109_53# _20_ 8.12e-19
C1745 _22_ _05_ 3.33e-21
C1746 _21_ b[2] 2.14e-19
C1747 input3/a_27_47# output19/a_27_47# 4.77e-21
C1748 net5 _09_ 5.18e-19
C1749 b[2] _24_ 1.85e-19
C1750 _08_ _05_ 0.00897f
C1751 _42_/a_109_93# _17_ 7.83e-20
C1752 _37_/a_27_47# net2 0.0692f
C1753 _10_ _50_/a_27_47# 0.0154f
C1754 net5 net6 0.722f
C1755 input5/a_664_47# net7 0.00199f
C1756 _39_/a_47_47# _20_ 2.3e-20
C1757 _02_ _12_ 0.265f
C1758 input4/a_75_212# _18_ 4.36e-19
C1759 net2 _22_ 1.93e-20
C1760 _03_ _12_ 2.76e-20
C1761 VPWR _40_/a_109_297# -4.23e-19
C1762 _06_ net4 0.281f
C1763 _17_ _44_/a_93_21# 0.0646f
C1764 net1 _55_/a_80_21# 1.8e-19
C1765 net8 _20_ 5.07e-19
C1766 _03_ _30_/a_297_297# 0.00117f
C1767 _04_ _30_/a_215_297# 0.00225f
C1768 _19_ _20_ 0.00734f
C1769 net5 net13 0.127f
C1770 _10_ net12 0.00257f
C1771 VPWR _34_/a_47_47# 0.0372f
C1772 _38_/a_27_47# _13_ 4.58e-19
C1773 _29_/a_29_53# net9 0.0205f
C1774 _32_/a_27_47# _47_/a_81_21# 5.06e-21
C1775 _26_/a_29_53# net18 2.57e-21
C1776 _32_/a_109_47# _01_ 0.00129f
C1777 _47_/a_299_297# _41_/a_59_75# 0.00146f
C1778 input8/a_27_47# p[1] 5.13e-20
C1779 _49_/a_315_47# net7 0.00706f
C1780 _06_ _07_ 0.185f
C1781 net19 net14 0.148f
C1782 _52_/a_250_297# _02_ 0.0128f
C1783 _40_/a_109_297# net15 0.0016f
C1784 _05_ _09_ 0.0683f
C1785 _44_/a_346_47# net14 0.00464f
C1786 _50_/a_343_93# net4 0.00124f
C1787 net4 _18_ 0.023f
C1788 _50_/a_223_47# net6 0.0194f
C1789 _06_ input6/a_27_47# 2.85e-19
C1790 net10 input10/a_27_47# 0.00321f
C1791 input11/a_27_47# p[4] 0.0646f
C1792 _26_/a_183_297# _22_ 0.00184f
C1793 _21_ net4 0.00535f
C1794 _29_/a_29_53# _22_ 2.24e-21
C1795 input5/a_664_47# VPWR 0.00488f
C1796 _06_ _33_/a_209_311# 0.0187f
C1797 p[4] p[7] 7.8e-20
C1798 _09_ _49_/a_544_297# 2.56e-20
C1799 net4 _24_ 8.65e-20
C1800 net5 _13_ 0.0352f
C1801 _16_ net7 7.5e-20
C1802 _43_/a_193_413# net7 3.49e-19
C1803 _05_ net13 0.192f
C1804 VPWR _47_/a_299_297# 0.0643f
C1805 p[11] _11_ 4.18e-20
C1806 _36_/a_303_47# _06_ 5.3e-19
C1807 _06_ _50_/a_515_93# 0.00244f
C1808 net2 net6 0.00139f
C1809 _27_/a_109_297# VPWR -2.45e-19
C1810 net10 _30_/a_215_297# 0.0512f
C1811 _27_/a_27_297# net11 1.58e-20
C1812 _21_ _07_ 0.133f
C1813 _32_/a_27_47# _43_/a_27_47# 2.01e-20
C1814 _15_ net14 0.225f
C1815 _17_ _12_ 0.0109f
C1816 _49_/a_544_297# net13 3.43e-19
C1817 input5/a_381_47# net3 0.0299f
C1818 input5/a_664_47# net15 0.0216f
C1819 _07_ _24_ 5.67e-19
C1820 _49_/a_315_47# VPWR 6.26e-19
C1821 _30_/a_392_297# net13 6.64e-20
C1822 input1/a_75_212# net7 3.77e-19
C1823 _10_ _00_ 0.301f
C1824 _33_/a_296_53# _05_ 4.53e-19
C1825 _10_ _44_/a_584_47# 1.14e-20
C1826 _34_/a_47_47# _53_/a_29_53# 5.88e-22
C1827 input5/a_62_47# net8 2.05e-19
C1828 _02_ _54_/a_75_212# 6.6e-20
C1829 _28_/a_109_297# _16_ 1.26e-19
C1830 _32_/a_197_47# net9 6.06e-19
C1831 _47_/a_299_297# net15 1.44e-20
C1832 _01_ net3 1.16e-19
C1833 input5/a_62_47# _19_ 0.00159f
C1834 _03_ _54_/a_75_212# 5.45e-21
C1835 _05_ _13_ 2.57e-20
C1836 _50_/a_223_47# _13_ 8.2e-20
C1837 _26_/a_29_53# _04_ 2.3e-21
C1838 net11 _25_ 0.0262f
C1839 _50_/a_27_47# net4 0.0239f
C1840 output19/a_27_47# _42_/a_109_93# 1.56e-20
C1841 _32_/a_27_47# _20_ 0.0069f
C1842 _55_/a_300_47# _01_ 0.00113f
C1843 VPWR net18 0.104f
C1844 _29_/a_29_53# _09_ 0.00488f
C1845 input5/a_558_47# _42_/a_109_93# 1.75e-19
C1846 input5/a_381_47# _42_/a_209_311# 3.88e-19
C1847 _16_ VPWR 0.126f
C1848 _37_/a_27_47# net19 0.0105f
C1849 _06_ _35_/a_76_199# 0.00425f
C1850 _29_/a_29_53# net6 1.4e-20
C1851 VPWR _43_/a_193_413# 0.0063f
C1852 _45_/a_27_47# _39_/a_47_47# 1.31e-19
C1853 VPWR _30_/a_465_297# -4.57e-19
C1854 net19 _22_ 2.17e-19
C1855 output19/a_27_47# _44_/a_93_21# 7.25e-20
C1856 net10 _34_/a_129_47# 0.003f
C1857 p[11] net3 0.00406f
C1858 input5/a_558_47# _44_/a_93_21# 2.71e-19
C1859 _10_ _14_ 0.0571f
C1860 net4 net12 2.57e-20
C1861 _45_/a_27_47# _52_/a_93_21# 1.18e-19
C1862 p[0] b[1] 0.00123f
C1863 _42_/a_296_53# net14 2.18e-19
C1864 _42_/a_209_311# _01_ 1.58e-19
C1865 net1 _30_/a_215_297# 0.00375f
C1866 _04_ net7 0.0602f
C1867 input1/a_75_212# VPWR 0.0786f
C1868 _29_/a_29_53# net13 0.00104f
C1869 _32_/a_109_47# _02_ 3.98e-19
C1870 _27_/a_27_297# _42_/a_109_93# 1.35e-20
C1871 _10_ _38_/a_109_47# 5.44e-19
C1872 _39_/a_47_47# _23_ 5.24e-21
C1873 net16 output16/a_27_47# 0.0101f
C1874 net14 _49_/a_201_297# 1.52e-19
C1875 _31_/a_35_297# net13 1.86e-20
C1876 input5/a_381_47# net5 0.0546f
C1877 input5/a_558_47# p[13] 0.00158f
C1878 b[3] _01_ 9.26e-20
C1879 _14_ p[9] 2.62e-21
C1880 _16_ _55_/a_217_297# 0.0017f
C1881 _16_ net15 0.214f
C1882 _04_ _36_/a_109_47# 2.39e-19
C1883 net9 _15_ 0.00113f
C1884 _52_/a_93_21# _23_ 0.0166f
C1885 net11 _20_ 0.00128f
C1886 _43_/a_193_413# net15 0.00169f
C1887 _37_/a_303_47# VPWR -3.13e-19
C1888 _18_ _35_/a_76_199# 6.82e-21
C1889 input5/a_62_47# output17/a_27_47# 1.02e-19
C1890 _05_ _35_/a_226_47# 0.0134f
C1891 _07_ net12 0.18f
C1892 _21_ _35_/a_76_199# 0.0175f
C1893 _37_/a_27_47# _15_ 1.11e-19
C1894 net5 _45_/a_205_47# 8.28e-20
C1895 _02_ _11_ 0.0621f
C1896 input8/a_27_47# input9/a_75_212# 3.09e-20
C1897 net5 _01_ 0.0779f
C1898 _06_ _45_/a_193_297# 0.00201f
C1899 _03_ input9/a_75_212# 9.32e-20
C1900 _26_/a_29_53# net10 3.48e-22
C1901 b[3] p[11] 0.243f
C1902 _15_ _22_ 0.0236f
C1903 VPWR _40_/a_297_297# -5.42e-19
C1904 _33_/a_209_311# net12 0.0769f
C1905 _06_ net14 1.94e-19
C1906 _41_/a_145_75# p[12] 0.00339f
C1907 input5/a_62_47# input3/a_27_47# 0.00179f
C1908 net18 _53_/a_29_53# 0.0118f
C1909 VPWR _04_ 0.456f
C1910 _37_/a_303_47# net15 0.00118f
C1911 _37_/a_109_47# net3 0.00212f
C1912 _55_/a_472_297# _20_ 0.00212f
C1913 net19 net6 0.00352f
C1914 _36_/a_303_47# net12 1.37e-19
C1915 _00_ net4 0.0166f
C1916 net17 _33_/a_209_311# 7.03e-21
C1917 _43_/a_297_47# VPWR -2.11e-19
C1918 net16 _39_/a_285_47# 1.29e-19
C1919 p[4] input10/a_27_47# 0.0215f
C1920 net11 output18/a_27_47# 6.84e-20
C1921 _40_/a_297_297# net15 4.08e-19
C1922 net14 _18_ 0.0147f
C1923 _50_/a_343_93# net14 1.07e-20
C1924 _12_ _45_/a_465_47# 0.00211f
C1925 _21_ net14 7.17e-21
C1926 _02_ net3 9.52e-20
C1927 _01_ _05_ 5.03e-19
C1928 _55_/a_300_47# _02_ 0.00371f
C1929 _04_ net15 0.0569f
C1930 _03_ net3 4.27e-20
C1931 input5/a_381_47# net2 0.0138f
C1932 p[14] net3 0.00446f
C1933 _47_/a_81_21# _12_ 0.00158f
C1934 p[5] input12/a_27_47# 0.00359f
C1935 p[0] output17/a_27_47# 0.00805f
C1936 input5/a_558_47# p[1] 1.61e-21
C1937 _12_ _47_/a_384_47# 9.51e-20
C1938 _01_ _49_/a_544_297# 0.00109f
C1939 _29_/a_29_53# _35_/a_226_47# 2.64e-19
C1940 input11/a_27_47# input10/a_27_47# 5.3e-19
C1941 _22_ _49_/a_201_297# 2.45e-20
C1942 _17_ _11_ 0.197f
C1943 net12 _35_/a_76_199# 0.0132f
C1944 _14_ net4 1.54e-20
C1945 _15_ net6 0.17f
C1946 input5/a_664_47# net8 0.0116f
C1947 net2 _01_ 2.72e-19
C1948 _42_/a_209_311# _02_ 9.92e-19
C1949 net9 _06_ 0.0505f
C1950 _38_/a_27_47# _02_ 0.00103f
C1951 p[10] net17 0.18f
C1952 input5/a_664_47# _19_ 2.19e-21
C1953 VPWR net10 0.362f
C1954 _38_/a_109_47# net4 7.32e-19
C1955 p[14] _42_/a_209_311# 3.45e-22
C1956 net16 VPWR 0.518f
C1957 _27_/a_27_297# p[1] 2.27e-19
C1958 b[3] _02_ 1.07e-19
C1959 _37_/a_27_47# _06_ 2.5e-20
C1960 _29_/a_183_297# net3 7.38e-21
C1961 net1 net7 0.0712f
C1962 _25_ _12_ 1.23e-20
C1963 p[14] b[3] 0.0645f
C1964 _36_/a_27_47# _30_/a_215_297# 7.13e-20
C1965 _10_ _36_/a_197_47# 1.54e-19
C1966 _10_ _50_/a_429_93# 0.00167f
C1967 net7 input7/a_27_47# 0.00318f
C1968 net2 p[11] 0.0204f
C1969 _06_ _22_ 0.124f
C1970 _48_/a_27_47# p[6] 2.22e-19
C1971 _43_/a_27_47# _12_ 2.33e-21
C1972 _27_/a_109_297# _19_ 7.54e-21
C1973 _08_ _33_/a_368_53# 5.04e-19
C1974 _45_/a_27_47# net11 3.64e-20
C1975 _45_/a_109_297# VPWR -0.011f
C1976 _14_ input6/a_27_47# 3.75e-21
C1977 net5 _02_ 0.233f
C1978 _49_/a_315_47# _19_ 1.33e-19
C1979 _06_ _08_ 0.0343f
C1980 net9 _50_/a_343_93# 6.64e-19
C1981 net9 _18_ 1.51e-19
C1982 net5 _03_ 1.04e-19
C1983 _10_ p[12] 0.0993f
C1984 VPWR _44_/a_250_297# 0.0231f
C1985 _29_/a_29_53# _01_ 8.33e-20
C1986 _21_ net9 0.0282f
C1987 _31_/a_35_297# _01_ 4.27e-19
C1988 net18 _52_/a_93_21# 8.21e-21
C1989 net11 _23_ 0.0461f
C1990 _37_/a_27_47# _18_ 3.31e-20
C1991 _17_ net3 0.0698f
C1992 p[12] p[9] 1.4e-19
C1993 input1/a_75_212# b[1] 4.16e-19
C1994 _09_ _49_/a_201_297# 1.74e-20
C1995 _15_ _13_ 3.69e-20
C1996 _52_/a_584_47# _02_ 0.00389f
C1997 _16_ net8 0.00624f
C1998 _07_ _49_/a_75_199# 4.05e-21
C1999 _12_ _20_ 3.9e-19
C2000 _27_/a_205_297# _04_ 6.42e-19
C2001 _15_ _50_/a_615_93# 0.00183f
C2002 VPWR net1 1.17f
C2003 _22_ _50_/a_343_93# 0.0597f
C2004 _22_ _18_ 0.0211f
C2005 _43_/a_193_413# net8 1.62e-20
C2006 input12/a_27_47# p[6] 0.0166f
C2007 _43_/a_193_413# _19_ 4.85e-21
C2008 _21_ _22_ 0.00314f
C2009 _10_ _41_/a_145_75# 5.18e-19
C2010 _04_ _35_/a_226_297# 4.51e-19
C2011 _22_ _24_ 0.0846f
C2012 input14/a_27_47# _44_/a_250_297# 8.25e-21
C2013 VPWR input7/a_27_47# 0.0768f
C2014 _44_/a_250_297# net15 8.86e-20
C2015 input5/a_62_47# _44_/a_93_21# 5.05e-20
C2016 net17 net14 5.43e-19
C2017 _21_ _08_ 0.00139f
C2018 _42_/a_209_311# _17_ 1.22e-19
C2019 _50_/a_223_47# _02_ 2.51e-20
C2020 net16 _53_/a_29_53# 2.04e-20
C2021 net10 _53_/a_29_53# 7.88e-22
C2022 _49_/a_201_297# net13 3.31e-19
C2023 _29_/a_111_297# _06_ 6.74e-20
C2024 _05_ _02_ 0.00163f
C2025 _03_ _50_/a_223_47# 1.41e-21
C2026 input8/a_27_47# _05_ 1.58e-19
C2027 _03_ _05_ 0.135f
C2028 b[3] _17_ 0.00637f
C2029 input5/a_841_47# net7 0.00193f
C2030 _06_ _09_ 0.0965f
C2031 input5/a_62_47# p[13] 0.0202f
C2032 _06_ net6 0.308f
C2033 net1 net15 7.44e-20
C2034 input5/a_381_47# net19 0.00173f
C2035 b[1] _04_ 5.79e-19
C2036 _03_ _49_/a_544_297# 0.00568f
C2037 _33_/a_368_53# net13 2.1e-20
C2038 _04_ _30_/a_109_53# 9.19e-21
C2039 _03_ _30_/a_392_297# 6.33e-19
C2040 input4/a_75_212# p[12] 0.02f
C2041 net15 input7/a_27_47# 1.88e-19
C2042 input2/a_27_47# _03_ 2.71e-19
C2043 _26_/a_29_53# _36_/a_27_47# 1.6e-19
C2044 net5 _17_ 0.00408f
C2045 VPWR _34_/a_377_297# -0.00192f
C2046 net2 _03_ 1.89e-19
C2047 net11 _34_/a_47_47# 0.0309f
C2048 _25_ _54_/a_75_212# 0.0247f
C2049 _00_ _45_/a_193_297# 4.38e-20
C2050 _06_ net13 0.0766f
C2051 net2 p[14] 1.38e-19
C2052 net19 _01_ 4.9e-19
C2053 _32_/a_197_47# _01_ 0.00156f
C2054 p[10] _49_/a_75_199# 2.29e-20
C2055 _00_ net14 4.11e-20
C2056 _18_ _09_ 7.01e-21
C2057 _44_/a_584_47# net14 7.2e-19
C2058 net9 net12 0.0596f
C2059 _50_/a_27_47# _22_ 0.0276f
C2060 _52_/a_256_47# _02_ 0.00344f
C2061 _04_ _52_/a_93_21# 2.35e-19
C2062 _50_/a_343_93# net6 0.00214f
C2063 _50_/a_429_93# net4 4.16e-19
C2064 _21_ _09_ 0.263f
C2065 net6 _18_ 0.166f
C2066 _47_/a_81_21# _11_ 0.0454f
C2067 net10 _35_/a_226_297# 2.48e-19
C2068 _21_ net6 2.92e-20
C2069 _06_ _33_/a_296_53# 1.11e-20
C2070 _04_ net8 0.02f
C2071 _07_ _33_/a_109_93# 3.2e-19
C2072 input5/a_841_47# VPWR 0.0775f
C2073 _09_ _24_ 0.0202f
C2074 _04_ _19_ 0.356f
C2075 net6 _24_ 0.00121f
C2076 _11_ _47_/a_384_47# 7.23e-20
C2077 net19 p[11] 0.00646f
C2078 input1/a_75_212# output17/a_27_47# 0.0101f
C2079 net9 net17 1.26e-20
C2080 p[12] net4 0.00758f
C2081 p[2] net7 0.00156f
C2082 _22_ net12 5.73e-20
C2083 _18_ net13 1.06e-20
C2084 _06_ _13_ 0.00188f
C2085 p[0] p[13] 1.88e-19
C2086 _29_/a_29_53# _02_ 6.76e-21
C2087 _31_/a_35_297# _02_ 0.00316f
C2088 _21_ net13 0.13f
C2089 _50_/a_223_47# _17_ 5.24e-20
C2090 _31_/a_35_297# _03_ 0.00749f
C2091 _31_/a_35_297# input8/a_27_47# 0.00955f
C2092 _08_ net12 0.0269f
C2093 _29_/a_29_53# _03_ 0.0414f
C2094 _06_ _50_/a_615_93# 0.00264f
C2095 p[8] input15/a_27_47# 7.57e-19
C2096 net10 _30_/a_109_53# 5.6e-20
C2097 VPWR p[4] 0.112f
C2098 _14_ net14 0.184f
C2099 _15_ _01_ 0.007f
C2100 _25_ _11_ 7.05e-19
C2101 output19/a_27_47# net3 0.00348f
C2102 _35_/a_226_47# _49_/a_201_297# 1.66e-20
C2103 input5/a_558_47# net3 0.0137f
C2104 input5/a_841_47# net15 0.00585f
C2105 _43_/a_27_47# _11_ 4.27e-19
C2106 VPWR _39_/a_129_47# -9.47e-19
C2107 net10 _39_/a_47_47# 4.72e-22
C2108 _45_/a_27_47# _12_ 0.0866f
C2109 p[12] input6/a_27_47# 2.78e-19
C2110 net16 _39_/a_47_47# 7.7e-20
C2111 _50_/a_27_47# _09_ 1.3e-19
C2112 net2 _17_ 0.181f
C2113 net10 _52_/a_93_21# 7.84e-20
C2114 _15_ p[11] 2.93e-19
C2115 VPWR _36_/a_27_47# -0.00832f
C2116 _50_/a_343_93# _13_ 5.63e-20
C2117 _18_ _13_ 0.019f
C2118 _47_/a_81_21# net3 6.66e-19
C2119 _10_ p[9] 0.00225f
C2120 _04_ output17/a_27_47# 0.027f
C2121 _10_ p[3] 1.37e-20
C2122 net11 net18 0.00221f
C2123 _00_ net9 0.00501f
C2124 _50_/a_27_47# net6 0.0428f
C2125 net10 net8 2.05e-21
C2126 VPWR input11/a_27_47# 0.0375f
C2127 net14 _49_/a_75_199# 3.67e-19
C2128 input5/a_558_47# _42_/a_209_311# 7.85e-20
C2129 _37_/a_109_47# net19 1.16e-20
C2130 _27_/a_27_297# net3 0.0166f
C2131 _21_ _13_ 1.69e-19
C2132 _12_ _23_ 0.00743f
C2133 _24_ _13_ 2.47e-19
C2134 VPWR p[2] 0.103f
C2135 _06_ _35_/a_226_47# 0.00487f
C2136 b[3] output19/a_27_47# 0.00809f
C2137 _37_/a_27_47# _00_ 6.15e-20
C2138 VPWR p[7] 0.0184f
C2139 _29_/a_111_297# net12 1.21e-19
C2140 net12 _09_ 0.0374f
C2141 _55_/a_80_21# net7 0.00163f
C2142 input3/a_27_47# _04_ 3.55e-19
C2143 net6 net12 0.00643f
C2144 _50_/a_27_47# net13 7.27e-21
C2145 output18/a_27_47# _54_/a_75_212# 2.28e-19
C2146 _11_ _20_ 0.268f
C2147 _33_/a_109_93# _35_/a_76_199# 3.08e-19
C2148 net10 _34_/a_285_47# 0.0454f
C2149 input5/a_664_47# _44_/a_93_21# 1.88e-20
C2150 _00_ _22_ 0.477f
C2151 net1 b[1] 1.78e-20
C2152 _42_/a_368_53# net14 7.39e-19
C2153 net1 _30_/a_109_53# 0.0297f
C2154 _27_/a_27_297# _42_/a_209_311# 4.7e-20
C2155 _01_ _49_/a_201_297# 0.0105f
C2156 input5/a_664_47# p[13] 8.06e-19
C2157 _32_/a_197_47# _02_ 3.78e-19
C2158 input5/a_558_47# net5 0.0597f
C2159 net19 _02_ 0.0474f
C2160 _10_ _38_/a_197_47# 6.29e-19
C2161 _32_/a_27_47# _04_ 1.43e-19
C2162 _16_ _55_/a_472_297# 3.71e-19
C2163 VPWR _53_/a_111_297# 1.11e-34
C2164 _52_/a_250_297# _23_ 3.17e-19
C2165 net19 p[14] 0.101f
C2166 _40_/a_191_297# _11_ 0.00207f
C2167 p[0] p[1] 0.187f
C2168 input5/a_381_47# _06_ 1.6e-19
C2169 net12 net13 0.363f
C2170 _37_/a_27_47# _14_ 0.00137f
C2171 _10_ input4/a_75_212# 0.00372f
C2172 _21_ _35_/a_226_47# 9.87e-19
C2173 net5 _47_/a_81_21# 4.59e-19
C2174 net10 output17/a_27_47# 1.31e-20
C2175 _50_/a_27_47# _13_ 0.00169f
C2176 _38_/a_27_47# _25_ 5.76e-19
C2177 _27_/a_27_297# net5 3.48e-19
C2178 _28_/a_109_297# _55_/a_80_21# 2.05e-20
C2179 net1 net8 0.381f
C2180 net5 _47_/a_384_47# 0.00129f
C2181 net1 _19_ 2.86e-19
C2182 net17 net13 5.21e-20
C2183 _14_ _22_ 0.00449f
C2184 _06_ _01_ 0.00157f
C2185 _33_/a_296_53# net12 1.23e-20
C2186 VPWR _55_/a_80_21# 0.0289f
C2187 net8 input7/a_27_47# 2.03e-21
C2188 net9 _49_/a_75_199# 0.00382f
C2189 _19_ input7/a_27_47# 3.12e-21
C2190 _37_/a_197_47# net3 0.0028f
C2191 net3 _20_ 4.07e-19
C2192 _04_ net11 0.078f
C2193 _15_ _02_ 0.101f
C2194 _16_ _44_/a_93_21# 0.00354f
C2195 _00_ _09_ 9.35e-21
C2196 _03_ _15_ 7.39e-20
C2197 p[14] _15_ 5.32e-19
C2198 net5 _25_ 6.42e-19
C2199 _43_/a_193_413# _44_/a_93_21# 0.0161f
C2200 _10_ net4 0.183f
C2201 _00_ net6 0.00178f
C2202 _43_/a_369_47# VPWR -3.75e-19
C2203 _32_/a_27_47# net10 2.76e-20
C2204 _22_ _49_/a_75_199# 9.85e-21
C2205 _40_/a_191_297# net3 1.89e-19
C2206 _55_/a_80_21# net15 0.00759f
C2207 _01_ _18_ 6.1e-20
C2208 input5/a_558_47# input2/a_27_47# 2.04e-20
C2209 _50_/a_429_93# net14 6.04e-21
C2210 _55_/a_80_21# _55_/a_217_297# 1.42e-32
C2211 _50_/a_343_93# _01_ 0.0131f
C2212 _42_/a_209_311# _20_ 1.66e-20
C2213 _41_/a_59_75# input15/a_27_47# 3.96e-20
C2214 net2 output19/a_27_47# 0.00168f
C2215 input5/a_558_47# net2 5.99e-21
C2216 net19 _17_ 0.0269f
C2217 _21_ _01_ 7.94e-19
C2218 _47_/a_299_297# _12_ 0.00805f
C2219 b[3] _20_ 1.37e-19
C2220 input5/a_664_47# p[1] 1.21e-20
C2221 net1 output17/a_27_47# 8.12e-19
C2222 input3/a_27_47# _44_/a_250_297# 2.07e-19
C2223 _10_ _07_ 2.19e-19
C2224 _44_/a_346_47# _17_ 7.2e-19
C2225 input1/a_75_212# p[13] 4.16e-19
C2226 _10_ input6/a_27_47# 4.57e-20
C2227 _14_ net6 2.11e-19
C2228 _27_/a_27_297# input2/a_27_47# 1.16e-19
C2229 net12 _35_/a_226_47# 8.29e-19
C2230 _47_/a_81_21# net2 4.95e-19
C2231 input5/a_841_47# net8 0.025f
C2232 net5 _20_ 0.0651f
C2233 _27_/a_27_297# net2 0.0131f
C2234 net16 net11 4.43e-22
C2235 net10 net11 0.592f
C2236 _04_ _42_/a_109_93# 5.77e-22
C2237 _45_/a_27_47# _11_ 0.0703f
C2238 input6/a_27_47# p[9] 0.0762f
C2239 _38_/a_197_47# net4 7.64e-19
C2240 VPWR input15/a_27_47# 0.0113f
C2241 input8/a_27_47# _49_/a_201_297# 2.46e-21
C2242 _03_ _49_/a_201_297# 0.00842f
C2243 _00_ _13_ 3.77e-20
C2244 net18 _12_ 8.24e-19
C2245 net9 _33_/a_109_93# 0.00211f
C2246 input4/a_75_212# net4 0.0189f
C2247 p[5] input13/a_27_47# 3.09e-19
C2248 _04_ _44_/a_93_21# 4.47e-21
C2249 _09_ _49_/a_75_199# 2.93e-19
C2250 _10_ _36_/a_303_47# 4.09e-19
C2251 _32_/a_27_47# net1 0.0211f
C2252 _10_ _50_/a_515_93# 0.00129f
C2253 _15_ _17_ 0.0752f
C2254 _11_ _23_ 2e-20
C2255 VPWR input10/a_27_47# 0.00986f
C2256 _43_/a_193_413# _12_ 7.94e-22
C2257 _38_/a_27_47# output18/a_27_47# 8.6e-19
C2258 _45_/a_109_297# net11 7.46e-20
C2259 VPWR _35_/a_489_413# -0.00725f
C2260 input9/a_75_212# input13/a_27_47# 0.00732f
C2261 input5/a_62_47# net3 0.00164f
C2262 net15 input15/a_27_47# 0.00325f
C2263 _22_ _33_/a_109_93# 1.34e-22
C2264 net2 _43_/a_27_47# 0.01f
C2265 _06_ _02_ 0.85f
C2266 _03_ _06_ 0.00635f
C2267 _06_ p[14] 1.04e-19
C2268 _36_/a_27_47# net8 1.52e-19
C2269 _49_/a_75_199# net13 3.2e-19
C2270 _05_ _20_ 6.79e-19
C2271 _50_/a_223_47# _20_ 1.71e-19
C2272 p[8] VPWR 0.208f
C2273 _14_ _13_ 1.47e-20
C2274 _01_ net12 1.67e-21
C2275 input5/a_381_47# net17 1.37e-20
C2276 VPWR _30_/a_215_297# -0.00472f
C2277 p[2] net8 0.00956f
C2278 _27_/a_277_297# _04_ 0.00113f
C2279 net1 net11 1.13e-19
C2280 _10_ _35_/a_76_199# 7.19e-20
C2281 input5/a_62_47# b[3] 0.00324f
C2282 _40_/a_109_297# _11_ 0.00522f
C2283 _48_/a_27_47# _06_ 0.0251f
C2284 input1/a_75_212# p[1] 0.0023f
C2285 net17 _01_ 0.0988f
C2286 _37_/a_197_47# net2 4.74e-20
C2287 _50_/a_343_93# _02_ 6.94e-19
C2288 _18_ _02_ 2.96e-20
C2289 p[12] _22_ 2.13e-21
C2290 net2 _20_ 8.83e-19
C2291 _03_ _18_ 7.25e-23
C2292 _21_ _02_ 0.397f
C2293 input14/a_27_47# p[8] 0.0159f
C2294 input5/a_62_47# net5 0.00329f
C2295 _21_ _03_ 0.0818f
C2296 p[8] net15 3.39e-19
C2297 _02_ _24_ 0.023f
C2298 net19 output19/a_27_47# 0.0279f
C2299 input5/a_558_47# net19 2.24e-20
C2300 _04_ _12_ 1.42e-19
C2301 _03_ _24_ 9.46e-20
C2302 _40_/a_191_297# net2 0.00143f
C2303 _33_/a_109_93# _09_ 7.36e-20
C2304 _44_/a_250_297# _42_/a_109_93# 6.38e-19
C2305 input13/a_27_47# p[6] 1.07e-19
C2306 VPWR _34_/a_129_47# -9.47e-19
C2307 _10_ _45_/a_193_297# 0.0047f
C2308 net18 _54_/a_75_212# 0.0143f
C2309 _06_ input12/a_27_47# 5.3e-22
C2310 _21_ _48_/a_27_47# 0.0121f
C2311 _04_ p[1] 1.74e-21
C2312 _44_/a_250_297# _44_/a_93_21# -6.97e-22
C2313 _06_ _17_ 0.0341f
C2314 VPWR output16/a_27_47# 0.122f
C2315 _55_/a_80_21# net8 1.84e-21
C2316 _29_/a_29_53# _20_ 0.0111f
C2317 _27_/a_27_297# net19 1.98e-19
C2318 _00_ _01_ 0.00124f
C2319 _10_ net14 2.4e-19
C2320 _40_/a_109_297# net3 3.14e-19
C2321 _45_/a_27_47# net5 0.0288f
C2322 _04_ _52_/a_250_297# 3.98e-21
C2323 _31_/a_35_297# _20_ 1.69e-19
C2324 _33_/a_109_93# net13 0.0254f
C2325 _36_/a_197_47# net6 6.94e-20
C2326 _50_/a_429_93# net6 6.18e-19
C2327 _47_/a_299_297# _11_ 0.00738f
C2328 p[13] _44_/a_250_297# 4.09e-20
C2329 _07_ _33_/a_209_311# 0.00859f
C2330 _32_/a_303_47# net9 0.00218f
C2331 net14 p[9] 1.05e-19
C2332 _35_/a_226_47# _49_/a_75_199# 8.73e-20
C2333 input5/a_558_47# _15_ 0.00166f
C2334 input5/a_381_47# _14_ 5.68e-20
C2335 net5 _23_ 0.0052f
C2336 _50_/a_27_47# _02_ 2.09e-19
C2337 _32_/a_27_47# _36_/a_27_47# 0.011f
C2338 p[12] net6 0.0941f
C2339 _26_/a_29_53# VPWR 0.0356f
C2340 _36_/a_197_47# net13 1.06e-19
C2341 net1 p[13] 2.13e-19
C2342 net10 _12_ 7.82e-20
C2343 _17_ _18_ 0.271f
C2344 net16 _12_ 0.131f
C2345 _21_ input12/a_27_47# 2.32e-19
C2346 _50_/a_343_93# _17_ 0.0015f
C2347 p[5] net18 1.98e-19
C2348 net11 p[4] 0.0557f
C2349 _31_/a_117_297# _03_ 5.32e-19
C2350 _47_/a_81_21# _15_ 0.00332f
C2351 _34_/a_47_47# p[6] 4.28e-19
C2352 net10 _30_/a_297_297# 1.68e-19
C2353 input5/a_62_47# net2 0.0197f
C2354 net12 _02_ 2.28e-19
C2355 _14_ _01_ 0.0193f
C2356 _03_ net12 0.0268f
C2357 input5/a_664_47# net3 0.00215f
C2358 _27_/a_27_297# _15_ 9.85e-20
C2359 _15_ _47_/a_384_47# 0.00112f
C2360 _45_/a_27_47# _05_ 9.34e-23
C2361 _16_ _11_ 4.42e-20
C2362 VPWR net7 0.784f
C2363 _26_/a_29_53# net15 9.06e-21
C2364 _45_/a_109_297# _12_ 0.00587f
C2365 _43_/a_193_413# _11_ 5.45e-19
C2366 VPWR _39_/a_285_47# -9.53e-19
C2367 net17 _02_ 0.0608f
C2368 net10 _52_/a_250_297# 2.86e-21
C2369 VPWR _36_/a_109_47# -4.66e-19
C2370 _14_ p[11] 7.85e-20
C2371 net11 _36_/a_27_47# 0.0717f
C2372 _03_ net17 5.1e-19
C2373 _10_ net9 0.0438f
C2374 _47_/a_299_297# net3 2.55e-19
C2375 VPWR _41_/a_59_75# 0.0179f
C2376 net11 input11/a_27_47# 0.00318f
C2377 _05_ input13/a_27_47# 3.93e-19
C2378 net16 b[0] 0.0306f
C2379 _48_/a_27_47# net12 0.0126f
C2380 input5/a_664_47# _42_/a_209_311# 0.0124f
C2381 _27_/a_109_297# net3 5.45e-19
C2382 net19 _20_ 1.29e-19
C2383 _01_ _49_/a_75_199# 0.009f
C2384 _07_ _35_/a_76_199# 0.00226f
C2385 net7 net15 2.91e-19
C2386 p[3] net9 0.0376f
C2387 _15_ _43_/a_27_47# 8.96e-20
C2388 _55_/a_217_297# net7 1.04e-19
C2389 _37_/a_27_47# p[9] 0.0117f
C2390 _10_ _22_ 0.0904f
C2391 _33_/a_109_93# _35_/a_226_47# 4.9e-19
C2392 _33_/a_209_311# _35_/a_76_199# 9.95e-21
C2393 _50_/a_27_47# _17_ 3.93e-20
C2394 net1 _30_/a_297_297# 7.34e-20
C2395 _28_/a_109_297# VPWR -1.71e-19
C2396 net4 _45_/a_193_297# 7.41e-19
C2397 _41_/a_59_75# net15 1.16e-20
C2398 input5/a_841_47# p[13] 1.73e-19
C2399 _16_ net3 1.77e-19
C2400 net4 net14 2.21e-21
C2401 input5/a_664_47# net5 0.0536f
C2402 _10_ _08_ 1.51e-19
C2403 _10_ _38_/a_303_47# 7.36e-19
C2404 _31_/a_285_297# net13 3.85e-20
C2405 _52_/a_256_47# _23_ 6.66e-19
C2406 _40_/a_297_297# _11_ 9.94e-19
C2407 _00_ _02_ 0.0269f
C2408 _00_ _03_ 2.31e-20
C2409 _06_ output19/a_27_47# 1.53e-19
C2410 net1 p[1] 0.0291f
C2411 input12/a_27_47# net12 0.0295f
C2412 input5/a_558_47# _06_ 3.55e-19
C2413 _43_/a_193_413# net3 5.65e-20
C2414 _37_/a_197_47# _15_ 3.02e-19
C2415 _15_ _20_ 0.691f
C2416 input7/a_27_47# p[1] 0.0164f
C2417 _30_/a_215_297# net8 8.14e-21
C2418 net5 _47_/a_299_297# 0.00198f
C2419 _04_ input9/a_75_212# 7.69e-22
C2420 _34_/a_47_47# _05_ 1.26e-20
C2421 net10 _54_/a_75_212# 6.24e-19
C2422 net16 _54_/a_75_212# 1.69e-21
C2423 _38_/a_27_47# net18 0.00997f
C2424 _16_ _42_/a_209_311# 0.00129f
C2425 input14/a_27_47# VPWR 0.0735f
C2426 _47_/a_81_21# _06_ 0.0388f
C2427 _22_ b[2] 0.0043f
C2428 _40_/a_109_297# net2 0.0011f
C2429 VPWR net15 0.61f
C2430 VPWR _55_/a_217_297# -0.00133f
C2431 _16_ b[3] 2.9e-19
C2432 input6/a_27_47# net14 7.05e-19
C2433 _49_/a_208_47# net7 0.00312f
C2434 _37_/a_303_47# net3 0.00133f
C2435 _14_ _02_ 0.0316f
C2436 _10_ _09_ 0.0222f
C2437 p[14] _14_ 1.66e-20
C2438 _10_ net6 0.0965f
C2439 _43_/a_469_47# VPWR -2.75e-19
C2440 _38_/a_109_47# _02_ 1.63e-19
C2441 _16_ net5 1.99e-20
C2442 _06_ _25_ 0.144f
C2443 _40_/a_297_297# net3 2.54e-19
C2444 net5 _43_/a_193_413# 1.39e-20
C2445 _55_/a_217_297# net15 7.79e-19
C2446 _47_/a_299_297# _50_/a_223_47# 2.74e-20
C2447 _47_/a_81_21# _18_ 7.96e-20
C2448 _47_/a_81_21# _50_/a_343_93# 0.00282f
C2449 input5/a_664_47# input2/a_27_47# 4.47e-21
C2450 net9 net4 1.99e-22
C2451 _50_/a_515_93# net14 1.39e-20
C2452 net6 p[9] 0.14f
C2453 net10 p[5] 0.00544f
C2454 VPWR _53_/a_29_53# 0.00821f
C2455 _02_ _49_/a_75_199# 0.0354f
C2456 _04_ net3 0.113f
C2457 _49_/a_201_297# _20_ 5.24e-21
C2458 _10_ net13 0.00151f
C2459 _06_ _43_/a_27_47# 0.0329f
C2460 input5/a_664_47# net2 8.11e-20
C2461 input8/a_27_47# _49_/a_75_199# 1.99e-20
C2462 _03_ _49_/a_75_199# 0.0849f
C2463 net16 _11_ 0.172f
C2464 _00_ _17_ 0.0851f
C2465 net10 input9/a_75_212# 0.00699f
C2466 _09_ b[2] 4.28e-20
C2467 p[3] net13 9.49e-19
C2468 _43_/a_469_47# net15 7.41e-19
C2469 p[10] net14 3.02e-19
C2470 VPWR _49_/a_208_47# -5.93e-19
C2471 _22_ net4 0.0866f
C2472 p[8] input3/a_27_47# 6.2e-19
C2473 _47_/a_299_297# net2 1.18e-19
C2474 _39_/a_129_47# _12_ 0.00175f
C2475 b[1] net7 0.005f
C2476 net9 _07_ 1.39e-20
C2477 _27_/a_109_297# net2 7.24e-20
C2478 _04_ _42_/a_209_311# 9.84e-22
C2479 _45_/a_109_297# _11_ 0.00168f
C2480 _38_/a_303_47# net4 5.95e-19
C2481 _36_/a_27_47# _12_ 0.00178f
C2482 _21_ _25_ 0.00164f
C2483 _06_ _20_ 0.133f
C2484 _10_ _13_ 0.0621f
C2485 net9 _33_/a_209_311# 4.33e-20
C2486 _43_/a_27_47# _18_ 0.0201f
C2487 _37_/a_27_47# input6/a_27_47# 9.35e-19
C2488 _27_/a_205_297# VPWR 1.05e-19
C2489 input4/a_75_212# net6 0.0273f
C2490 net11 input10/a_27_47# 0.112f
C2491 _10_ _50_/a_615_93# 8.82e-19
C2492 _14_ _17_ 0.489f
C2493 _07_ _22_ 1.19e-20
C2494 VPWR _35_/a_226_297# -8.54e-19
C2495 _40_/a_191_297# _06_ 5.84e-19
C2496 net8 net7 0.295f
C2497 _07_ _08_ 0.348f
C2498 _16_ net2 0.00654f
C2499 net5 _04_ 0.00476f
C2500 net7 _19_ 0.0458f
C2501 b[0] _39_/a_129_47# 2.6e-20
C2502 net1 input9/a_75_212# 0.002f
C2503 net2 _43_/a_193_413# 1.52e-19
C2504 p[2] p[1] 0.188f
C2505 _18_ _20_ 0.0151f
C2506 _50_/a_343_93# _20_ 0.00826f
C2507 _31_/a_285_297# _01_ 1.92e-19
C2508 _21_ _20_ 0.191f
C2509 input5/a_558_47# net17 2.88e-21
C2510 VPWR b[1] 0.396f
C2511 _08_ _33_/a_209_311# 0.0122f
C2512 _48_/a_181_47# VPWR -3.35e-19
C2513 _48_/a_109_47# net11 1.74e-19
C2514 net4 _09_ 0.00262f
C2515 _33_/a_109_93# _02_ 1.54e-21
C2516 _04_ _52_/a_584_47# 2.5e-19
C2517 net11 _30_/a_215_297# 1.04e-19
C2518 VPWR _30_/a_109_53# 0.0012f
C2519 net10 p[6] 0.0023f
C2520 _03_ _33_/a_109_93# 2.78e-19
C2521 net4 net6 0.713f
C2522 _10_ _35_/a_226_47# 1.25e-19
C2523 net16 _38_/a_27_47# 0.114f
C2524 _32_/a_303_47# _01_ 8.58e-19
C2525 _06_ output18/a_27_47# 0.0114f
C2526 _44_/a_250_297# net3 0.0088f
C2527 VPWR _39_/a_47_47# 0.0668f
C2528 _37_/a_303_47# net2 4.41e-19
C2529 _27_/a_27_297# net17 0.00181f
C2530 _04_ _50_/a_223_47# 7.89e-22
C2531 net4 net13 2.48e-19
C2532 VPWR _52_/a_93_21# -0.00838f
C2533 _04_ _05_ 0.0352f
C2534 _07_ _09_ 0.0405f
C2535 VPWR net8 0.703f
C2536 net12 _25_ 4.46e-20
C2537 VPWR _19_ 0.0335f
C2538 net1 net3 4.25e-20
C2539 output17/a_27_47# net7 0.00185f
C2540 input5/a_664_47# net19 1.38e-21
C2541 input6/a_27_47# net6 0.00208f
C2542 _40_/a_297_297# net2 0.00101f
C2543 net16 net5 0.00461f
C2544 net5 net10 0.0316f
C2545 _04_ _49_/a_544_297# 0.00204f
C2546 p[12] p[14] 0.00101f
C2547 _33_/a_209_311# _09_ 3.79e-20
C2548 input2/a_27_47# _04_ 4.5e-21
C2549 _22_ _35_/a_76_199# 6.58e-21
C2550 _39_/a_47_47# net15 9.44e-22
C2551 net11 _34_/a_129_47# 0.00242f
C2552 VPWR _34_/a_285_47# -0.00233f
C2553 _21_ output18/a_27_47# 0.00103f
C2554 b[3] _44_/a_250_297# 0.0112f
C2555 net2 _04_ 0.158f
C2556 _07_ net13 0.00686f
C2557 _10_ _45_/a_205_47# 6.19e-20
C2558 net1 p[6] 3.12e-20
C2559 _08_ _35_/a_76_199# 0.0061f
C2560 net8 net15 0.2f
C2561 _10_ _01_ 2.22e-19
C2562 _45_/a_109_297# net5 0.0184f
C2563 _00_ _47_/a_81_21# 0.0258f
C2564 net4 _13_ 0.212f
C2565 net15 _19_ 0.00628f
C2566 _50_/a_515_93# net6 4.7e-19
C2567 _36_/a_303_47# net6 1.25e-19
C2568 _00_ _47_/a_384_47# 5.15e-20
C2569 p[5] p[4] 0.385f
C2570 _33_/a_209_311# net13 0.0227f
C2571 _45_/a_27_47# _06_ 0.0021f
C2572 net5 _44_/a_250_297# 3.11e-20
C2573 _32_/a_27_47# net7 0.00559f
C2574 net12 _20_ 0.00437f
C2575 net9 net14 7.12e-20
C2576 _14_ output19/a_27_47# 1.43e-19
C2577 input5/a_664_47# _15_ 9.15e-22
C2578 net16 _50_/a_223_47# 4.77e-21
C2579 VPWR output17/a_27_47# 0.0263f
C2580 p[8] p[13] 0.00172f
C2581 _26_/a_29_53# net11 1.08e-20
C2582 net10 _05_ 0.457f
C2583 _06_ _23_ 0.218f
C2584 _37_/a_27_47# net14 0.0584f
C2585 _06_ input13/a_27_47# 7.75e-19
C2586 _07_ _13_ 3.22e-23
C2587 _36_/a_303_47# net13 5.5e-20
C2588 net17 _20_ 4e-20
C2589 _16_ net19 0.206f
C2590 _52_/a_93_21# _53_/a_29_53# 0.00116f
C2591 _22_ _45_/a_193_297# 0.0234f
C2592 net1 net5 0.0772f
C2593 p[11] p[9] 0.114f
C2594 _31_/a_285_297# _02_ 5.86e-20
C2595 _29_/a_29_53# _04_ 0.0408f
C2596 _47_/a_81_21# _14_ 6.24e-20
C2597 _47_/a_299_297# _15_ 0.0103f
C2598 _31_/a_285_297# input8/a_27_47# 1.04e-19
C2599 input11/a_27_47# p[5] 0.0433f
C2600 _31_/a_35_297# _04_ 1.89e-20
C2601 _31_/a_285_297# _03_ 0.00677f
C2602 net10 _30_/a_392_297# 3.4e-19
C2603 net19 _43_/a_193_413# 3.31e-19
C2604 _22_ net14 2.23e-19
C2605 _34_/a_377_297# p[6] 5.39e-19
C2606 net10 input2/a_27_47# 1.17e-20
C2607 _09_ _35_/a_76_199# 0.0374f
C2608 VPWR input3/a_27_47# 0.0687f
C2609 _00_ _43_/a_27_47# 0.0431f
C2610 net6 _35_/a_76_199# 4.6e-21
C2611 _27_/a_27_297# _14_ 1.66e-21
C2612 _45_/a_27_47# _18_ 0.00347f
C2613 p[5] p[7] 6.77e-20
C2614 net10 net2 2.05e-20
C2615 _45_/a_109_297# _05_ 2.79e-22
C2616 _21_ _45_/a_27_47# 1.18e-20
C2617 net11 net7 1.77e-19
C2618 _32_/a_303_47# _02_ 1.15e-20
C2619 p[2] input9/a_75_212# 5.13e-20
C2620 _45_/a_27_47# _24_ 4.57e-19
C2621 input9/a_75_212# p[7] 0.00102f
C2622 _49_/a_208_47# net8 1.4e-19
C2623 VPWR _32_/a_27_47# 0.0395f
C2624 _49_/a_208_47# _19_ 7.12e-20
C2625 net10 _52_/a_256_47# 8.13e-20
C2626 _40_/a_109_297# _06_ 0.00175f
C2627 _35_/a_76_199# net13 0.0337f
C2628 _21_ _23_ 0.0217f
C2629 input3/a_27_47# net15 6.19e-20
C2630 _24_ _23_ 0.012f
C2631 input14/a_27_47# input3/a_27_47# 5.08e-20
C2632 _27_/a_27_297# _49_/a_75_199# 0.011f
C2633 _07_ _35_/a_226_47# 8.96e-19
C2634 _16_ _15_ 0.0607f
C2635 _00_ _20_ 0.271f
C2636 net1 _05_ 0.151f
C2637 net2 _44_/a_250_297# 0.0169f
C2638 _14_ _43_/a_27_47# 0.00938f
C2639 _15_ _43_/a_193_413# 4.86e-19
C2640 _06_ _34_/a_47_47# 0.0391f
C2641 _09_ _45_/a_193_297# 0.00961f
C2642 p[4] p[6] 0.0051f
C2643 _30_/a_215_297# _30_/a_297_297# -8.88e-34
C2644 _29_/a_29_53# net10 1.77e-19
C2645 net1 _49_/a_544_297# 0.00175f
C2646 _33_/a_209_311# _35_/a_226_47# 1.31e-19
C2647 net10 _31_/a_35_297# 3.95e-20
C2648 net6 _45_/a_193_297# 9.84e-20
C2649 net1 input2/a_27_47# 4.81e-19
C2650 VPWR net11 0.996f
C2651 net6 net14 2.82e-21
C2652 input5/a_841_47# net5 0.0221f
C2653 _45_/a_27_47# _50_/a_27_47# 0.109f
C2654 _04_ net19 2.07e-20
C2655 net1 net2 1.64e-19
C2656 net9 _22_ 0.0023f
C2657 _35_/a_76_199# _13_ 3.01e-21
C2658 _10_ _02_ 0.0537f
C2659 input2/a_27_47# input7/a_27_47# 1.62e-19
C2660 input5/a_664_47# _06_ 3.21e-19
C2661 _10_ _03_ 0.00244f
C2662 _10_ p[14] 1.53e-19
C2663 _31_/a_285_47# net7 0.00132f
C2664 _14_ _20_ 0.144f
C2665 net2 input7/a_27_47# 3.24e-19
C2666 b[1] net8 0.00195f
C2667 net9 _08_ 7.71e-21
C2668 _30_/a_109_53# net8 1.76e-20
C2669 input8/a_27_47# p[3] 0.0023f
C2670 net14 net13 2.21e-21
C2671 p[14] p[9] 0.4f
C2672 _03_ p[3] 0.00348f
C2673 _21_ _34_/a_47_47# 8.93e-19
C2674 _47_/a_299_297# _06_ 0.0174f
C2675 _39_/a_47_47# _52_/a_93_21# 1.44e-20
C2676 p[7] p[6] 0.217f
C2677 _34_/a_47_47# _24_ 6.84e-21
C2678 _40_/a_191_297# _14_ 2.4e-19
C2679 VPWR _55_/a_472_297# 0.00488f
C2680 _10_ _48_/a_27_47# 4.55e-19
C2681 p[13] net7 1.91e-19
C2682 input10/a_27_47# _54_/a_75_212# 1.17e-22
C2683 _29_/a_183_297# _10_ 6.24e-20
C2684 net5 _39_/a_129_47# 0.00344f
C2685 net12 _23_ 2.28e-21
C2686 input5/a_664_47# _18_ 1.09e-20
C2687 net12 input13/a_27_47# 0.0163f
C2688 _20_ _49_/a_75_199# 0.0233f
C2689 b[2] _02_ 2.69e-19
C2690 _21_ input5/a_664_47# 9.42e-22
C2691 _29_/a_29_53# net1 9.76e-19
C2692 _04_ _15_ 3.61e-20
C2693 net5 _36_/a_27_47# 0.0163f
C2694 net8 _19_ 0.0322f
C2695 net1 _31_/a_35_297# 0.0111f
C2696 _29_/a_111_297# net9 8.06e-21
C2697 VPWR _42_/a_109_93# -0.00118f
C2698 p[12] output19/a_27_47# 1.78e-19
C2699 _04_ VGND 0.478f
C2700 _03_ VGND 0.481f
C2701 net10 VGND 0.909f
C2702 _30_/a_465_297# VGND 0.00105f
C2703 _30_/a_392_297# VGND 7.67e-19
C2704 _30_/a_297_297# VGND -4.43e-19
C2705 _30_/a_109_53# VGND 0.152f
C2706 _30_/a_215_297# VGND 0.158f
C2707 _05_ VGND 0.906f
C2708 net8 VGND 0.791f
C2709 _31_/a_285_297# VGND 1.12e-20
C2710 _31_/a_117_297# VGND -0.00177f
C2711 _31_/a_35_297# VGND 0.246f
C2712 _32_/a_303_47# VGND -4.83e-19
C2713 _32_/a_197_47# VGND 8.12e-20
C2714 _32_/a_109_47# VGND 1.05e-19
C2715 _32_/a_27_47# VGND 0.198f
C2716 _50_/a_615_93# VGND -5.19e-19
C2717 _50_/a_515_93# VGND -4.75e-19
C2718 _50_/a_429_93# VGND 4.71e-19
C2719 _50_/a_343_93# VGND 0.171f
C2720 _50_/a_223_47# VGND 0.157f
C2721 _50_/a_27_47# VGND 0.255f
C2722 _07_ VGND 0.483f
C2723 _06_ VGND 1.91f
C2724 net13 VGND 0.524f
C2725 _33_/a_368_53# VGND 2.38e-19
C2726 _33_/a_296_53# VGND -1.43e-19
C2727 _33_/a_209_311# VGND 0.136f
C2728 _33_/a_109_93# VGND 0.145f
C2729 _08_ VGND 0.293f
C2730 net12 VGND 0.874f
C2731 _34_/a_285_47# VGND 0.0144f
C2732 _34_/a_129_47# VGND -8.76e-20
C2733 _34_/a_377_297# VGND -9.51e-19
C2734 _34_/a_47_47# VGND 0.289f
C2735 _23_ VGND 0.266f
C2736 p[9] VGND 0.51f
C2737 input15/a_27_47# VGND 0.223f
C2738 _09_ VGND 0.544f
C2739 _35_/a_556_47# VGND 1.95e-19
C2740 _35_/a_226_297# VGND -4.55e-19
C2741 _35_/a_489_413# VGND 0.0246f
C2742 _35_/a_226_47# VGND 0.151f
C2743 _35_/a_76_199# VGND 0.137f
C2744 _24_ VGND 0.127f
C2745 _12_ VGND 1.2f
C2746 _52_/a_584_47# VGND -0.00112f
C2747 _52_/a_346_47# VGND -0.00175f
C2748 _52_/a_256_47# VGND -0.00161f
C2749 _52_/a_250_297# VGND 0.0246f
C2750 _52_/a_93_21# VGND 0.133f
C2751 _10_ VGND 1.75f
C2752 _36_/a_303_47# VGND 8.14e-19
C2753 _36_/a_197_47# VGND -3.75e-19
C2754 _36_/a_109_47# VGND 3.56e-19
C2755 _36_/a_27_47# VGND 0.196f
C2756 p[8] VGND 1.26f
C2757 input14/a_27_47# VGND 0.247f
C2758 _53_/a_183_297# VGND -4.34e-19
C2759 _53_/a_111_297# VGND -2.89e-19
C2760 _53_/a_29_53# VGND 0.163f
C2761 _11_ VGND 0.358f
C2762 _37_/a_303_47# VGND -1.63e-19
C2763 _37_/a_197_47# VGND -4.58e-19
C2764 _37_/a_109_47# VGND -7.9e-19
C2765 _37_/a_27_47# VGND 0.16f
C2766 p[7] VGND 0.887f
C2767 input13/a_27_47# VGND 0.255f
C2768 net18 VGND 0.463f
C2769 _25_ VGND 0.39f
C2770 _54_/a_75_212# VGND 0.263f
C2771 _38_/a_303_47# VGND 1.78e-19
C2772 _38_/a_197_47# VGND 2.29e-19
C2773 _38_/a_109_47# VGND 2.3e-19
C2774 _38_/a_27_47# VGND 0.183f
C2775 net19 VGND 0.31f
C2776 _22_ VGND 0.256f
C2777 _14_ VGND 0.454f
C2778 _15_ VGND 0.487f
C2779 _55_/a_300_47# VGND -0.00109f
C2780 _55_/a_472_297# VGND -0.00188f
C2781 _55_/a_217_297# VGND -0.00225f
C2782 _55_/a_80_21# VGND 0.213f
C2783 p[6] VGND 0.742f
C2784 input12/a_27_47# VGND 0.248f
C2785 net9 VGND 0.685f
C2786 p[3] VGND 0.825f
C2787 input9/a_75_212# VGND 0.276f
C2788 _39_/a_285_47# VGND 0.0128f
C2789 _39_/a_129_47# VGND -0.00126f
C2790 _39_/a_377_297# VGND -6.28e-19
C2791 _39_/a_47_47# VGND 0.266f
C2792 net11 VGND 1.25f
C2793 p[5] VGND 0.76f
C2794 input11/a_27_47# VGND 0.235f
C2795 p[2] VGND 0.769f
C2796 input8/a_27_47# VGND 0.265f
C2797 p[4] VGND 1.25f
C2798 input10/a_27_47# VGND 0.211f
C2799 net7 VGND 0.881f
C2800 p[1] VGND 0.772f
C2801 input7/a_27_47# VGND 0.265f
C2802 p[14] VGND 0.988f
C2803 input6/a_27_47# VGND 0.205f
C2804 net5 VGND 2.04f
C2805 p[13] VGND 0.557f
C2806 input5/a_841_47# VGND 0.187f
C2807 input5/a_664_47# VGND 0.144f
C2808 input5/a_558_47# VGND 0.163f
C2809 input5/a_381_47# VGND 0.107f
C2810 input5/a_62_47# VGND 0.218f
C2811 p[12] VGND 1.3f
C2812 input4/a_75_212# VGND 0.263f
C2813 p[11] VGND 0.865f
C2814 input3/a_27_47# VGND 0.249f
C2815 net2 VGND 1.5f
C2816 p[10] VGND 0.79f
C2817 input2/a_27_47# VGND 0.194f
C2818 net1 VGND 0.855f
C2819 p[0] VGND 1.01f
C2820 VPWR VGND 40.2f
C2821 input1/a_75_212# VGND 0.268f
C2822 b[3] VGND 0.546f
C2823 output19/a_27_47# VGND 0.534f
C2824 b[2] VGND 0.593f
C2825 output18/a_27_47# VGND 0.601f
C2826 _40_/a_297_297# VGND -5.1e-19
C2827 _40_/a_191_297# VGND -9.29e-19
C2828 _40_/a_109_297# VGND -0.00181f
C2829 b[1] VGND 0.526f
C2830 net17 VGND 0.385f
C2831 output17/a_27_47# VGND 0.545f
C2832 _41_/a_145_75# VGND 3.75e-19
C2833 _41_/a_59_75# VGND 0.191f
C2834 b[0] VGND 0.708f
C2835 output16/a_27_47# VGND 0.616f
C2836 _16_ VGND 0.119f
C2837 _42_/a_368_53# VGND -4.05e-19
C2838 _42_/a_209_311# VGND 0.135f
C2839 _42_/a_109_93# VGND 0.153f
C2840 _17_ VGND 0.563f
C2841 _00_ VGND 0.516f
C2842 _43_/a_369_47# VGND -8.43e-19
C2843 _43_/a_297_47# VGND -1.33e-19
C2844 _43_/a_193_413# VGND 0.122f
C2845 _43_/a_27_47# VGND 0.209f
C2846 net6 VGND 1f
C2847 net4 VGND 0.888f
C2848 _26_/a_183_297# VGND 2.42e-19
C2849 _26_/a_111_297# VGND -2.75e-19
C2850 _26_/a_29_53# VGND 0.218f
C2851 _01_ VGND 0.244f
C2852 net14 VGND 0.958f
C2853 net3 VGND 0.786f
C2854 net15 VGND 0.673f
C2855 _27_/a_277_297# VGND -4.65e-19
C2856 _27_/a_205_297# VGND -3.36e-19
C2857 _27_/a_109_297# VGND -6.15e-19
C2858 _27_/a_27_297# VGND 0.147f
C2859 _18_ VGND 0.159f
C2860 _44_/a_584_47# VGND -0.00145f
C2861 _44_/a_346_47# VGND -0.00198f
C2862 _44_/a_256_47# VGND -0.00184f
C2863 _44_/a_250_297# VGND 0.0219f
C2864 _44_/a_93_21# VGND 0.128f
C2865 net16 VGND 0.375f
C2866 _13_ VGND 0.496f
C2867 _45_/a_465_47# VGND -8.14e-19
C2868 _45_/a_205_47# VGND -2.47e-19
C2869 _45_/a_193_297# VGND -0.00131f
C2870 _45_/a_109_297# VGND -0.00108f
C2871 _45_/a_27_47# VGND 0.187f
C2872 _28_/a_109_297# VGND -9.87e-19
C2873 _29_/a_183_297# VGND 4.41e-19
C2874 _29_/a_111_297# VGND -1.9e-19
C2875 _29_/a_29_53# VGND 0.234f
C2876 _19_ VGND 0.497f
C2877 _47_/a_384_47# VGND -2.05e-19
C2878 _47_/a_299_297# VGND 0.0344f
C2879 _47_/a_81_21# VGND 0.136f
C2880 _48_/a_181_47# VGND 3.03e-19
C2881 _48_/a_109_47# VGND 9.44e-19
C2882 _48_/a_27_47# VGND 0.232f
C2883 _21_ VGND 0.586f
C2884 _20_ VGND 0.709f
C2885 _02_ VGND 2.08f
C2886 _49_/a_315_47# VGND -0.0034f
C2887 _49_/a_208_47# VGND -0.00164f
C2888 _49_/a_544_297# VGND -0.00256f
C2889 _49_/a_201_297# VGND -5.82e-19
C2890 _49_/a_75_199# VGND 0.205f
.ends

.subckt sky130_fd_pr__nfet_01v8_D7Y3TR a_n63_n101# a_n33_n75# a_n249_n145# a_63_n75#
+ a_n125_n75#
X0 a_63_n75# a_n63_n101# a_n33_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.233 pd=2.12 as=0.124 ps=1.08 w=0.75 l=0.15
X1 a_n33_n75# a_n63_n101# a_n125_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.08 as=0.233 ps=2.12 w=0.75 l=0.15
C0 a_n63_n101# a_63_n75# 0.0104f
C1 a_n33_n75# a_63_n75# 0.113f
C2 a_n63_n101# a_n125_n75# 0.00451f
C3 a_n33_n75# a_n125_n75# 0.113f
C4 a_n33_n75# a_n63_n101# 0.0186f
C5 a_63_n75# a_n249_n145# 0.0963f
C6 a_n33_n75# a_n249_n145# 0.0361f
C7 a_n125_n75# a_n249_n145# 0.105f
C8 a_n63_n101# a_n249_n145# 0.294f
.ends

.subckt sky130_fd_pr__pfet_01v8_2ZD99F w_n349_n261# a_n153_n139# a_n211_n42# a_153_n42#
+ VSUBS
X0 a_153_n42# a_n153_n139# a_n211_n42# w_n349_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.53
C0 a_n153_n139# a_153_n42# 0.0177f
C1 w_n349_n261# a_153_n42# 0.0179f
C2 a_n211_n42# a_153_n42# 0.0169f
C3 w_n349_n261# a_n153_n139# 0.388f
C4 a_n211_n42# a_n153_n139# 0.0177f
C5 a_n211_n42# w_n349_n261# 0.034f
C6 a_153_n42# VSUBS 0.0558f
C7 a_n211_n42# VSUBS 0.0456f
C8 a_n153_n139# VSUBS 0.556f
C9 w_n349_n261# VSUBS 1.16f
.ends

.subckt sky130_fd_pr__nfet_01v8_2BW22M a_154_n42# a_n154_n130# a_n314_n182# a_n212_n42#
X0 a_154_n42# a_n154_n130# a_n212_n42# a_n314_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.54
C0 a_n154_n130# a_n212_n42# 0.0178f
C1 a_154_n42# a_n212_n42# 0.0169f
C2 a_154_n42# a_n154_n130# 0.0178f
C3 a_154_n42# a_n314_n182# 0.0737f
C4 a_n212_n42# a_n314_n182# 0.0816f
C5 a_n154_n130# a_n314_n182# 0.924f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJP3BL a_15_n150# w_n211_n369# a_n73_n150# a_n33_n247#
+ VSUBS
X0 a_15_n150# a_n33_n247# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.15
C0 a_n33_n247# a_15_n150# 0.0267f
C1 w_n211_n369# a_15_n150# 0.0292f
C2 a_n73_n150# a_15_n150# 0.242f
C3 w_n211_n369# a_n33_n247# 0.19f
C4 a_n73_n150# a_n33_n247# 0.0267f
C5 a_n73_n150# w_n211_n369# 0.0292f
C6 a_15_n150# VSUBS 0.126f
C7 a_n73_n150# VSUBS 0.126f
C8 a_n33_n247# VSUBS 0.146f
C9 w_n211_n369# VSUBS 1.02f
.ends

.subckt sky130_fd_pr__nfet_01v8_LH5FDA a_n150_n130# a_276_n182# a_n208_n42# a_150_n42#
X0 a_150_n42# a_n150_n130# a_n208_n42# a_276_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.5
C0 a_n150_n130# a_n208_n42# 0.0176f
C1 a_150_n42# a_n208_n42# 0.0172f
C2 a_150_n42# a_n150_n130# 0.0176f
C3 a_150_n42# a_276_n182# 0.0815f
C4 a_n208_n42# a_276_n182# 0.0736f
C5 a_n150_n130# a_276_n182# 0.904f
.ends

.subckt th02 Vin V02 Vp m1_983_133# m1_571_144# Vn
XXM0 Vin Vn Vn m1_983_133# m1_983_133# sky130_fd_pr__nfet_01v8_D7Y3TR
XXM1 Vp Vin m1_571_144# m1_983_133# Vn sky130_fd_pr__pfet_01v8_2ZD99F
XXM2 m1_571_144# Vp Vn Vp sky130_fd_pr__nfet_01v8_2BW22M
XXM3 V02 Vp Vp m1_983_133# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_983_133# Vn V02 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 Vin Vn 0.0263f
C1 Vin Vp 0.25f
C2 Vin V02 0.00845f
C3 Vin m1_983_133# 0.279f
C4 m1_571_144# Vn 0.00115f
C5 Vp m1_571_144# 0.176f
C6 V02 m1_571_144# 0.011f
C7 Vp Vn 0.0235f
C8 m1_983_133# m1_571_144# 0.0183f
C9 V02 Vn 0.00239f
C10 Vp V02 0.118f
C11 m1_983_133# Vn 0.216f
C12 Vp m1_983_133# 0.366f
C13 Vin m1_571_144# 0.332f
C14 m1_983_133# V02 0.155f
C15 Vn 0 0.263f
C16 V02 0 0.334f
C17 m1_983_133# 0 1.44f
C18 Vp 0 3.16f
C19 m1_571_144# 0 0.252f
C20 Vin 0 0.949f
.ends

.subckt sky130_fd_pr__nfet_01v8_2V6S9N a_n216_n42# a_158_n42# a_n158_n130# a_n284_n216#
X0 a_158_n42# a_n158_n130# a_n216_n42# a_n284_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.58
C0 a_n216_n42# a_n158_n130# 0.018f
C1 a_158_n42# a_n158_n130# 0.018f
C2 a_158_n42# a_n216_n42# 0.0165f
C3 a_158_n42# a_n284_n216# 0.0746f
C4 a_n216_n42# a_n284_n216# 0.0746f
C5 a_n158_n130# a_n284_n216# 0.981f
.ends

.subckt sky130_fd_pr__pfet_01v8_XYZSMQ a_n33_n255# a_15_n158# w_n211_n377# a_n73_n158#
+ VSUBS
X0 a_15_n158# a_n33_n255# a_n73_n158# w_n211_n377# sky130_fd_pr__pfet_01v8 ad=0.458 pd=3.74 as=0.458 ps=3.74 w=1.58 l=0.15
C0 a_n33_n255# w_n211_n377# 0.191f
C1 a_15_n158# w_n211_n377# 0.0299f
C2 a_n73_n158# w_n211_n377# 0.0299f
C3 a_15_n158# a_n33_n255# 0.0271f
C4 a_n73_n158# a_n33_n255# 0.0271f
C5 a_n73_n158# a_15_n158# 0.254f
C6 a_15_n158# VSUBS 0.132f
C7 a_n73_n158# VSUBS 0.132f
C8 a_n33_n255# VSUBS 0.146f
C9 w_n211_n377# VSUBS 1.04f
.ends

.subckt sky130_fd_pr__pfet_01v8_AZD9DW w_n353_n261# a_n157_n139# a_n215_n42# a_157_n42#
+ VSUBS
X0 a_157_n42# a_n157_n139# a_n215_n42# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.57
C0 a_n157_n139# w_n353_n261# 0.396f
C1 a_157_n42# w_n353_n261# 0.0323f
C2 a_n215_n42# w_n353_n261# 0.0179f
C3 a_157_n42# a_n157_n139# 0.0179f
C4 a_n215_n42# a_n157_n139# 0.0179f
C5 a_n215_n42# a_157_n42# 0.0166f
C6 a_157_n42# VSUBS 0.0468f
C7 a_n215_n42# VSUBS 0.0559f
C8 a_n157_n139# VSUBS 0.569f
C9 w_n353_n261# VSUBS 1.17f
.ends

.subckt sky130_fd_pr__nfet_01v8_T8HSQ7 a_n175_n297# a_15_n157# a_n33_n245# a_n73_n157#
X0 a_15_n157# a_n33_n245# a_n73_n157# a_n175_n297# sky130_fd_pr__nfet_01v8 ad=0.455 pd=3.72 as=0.455 ps=3.72 w=1.57 l=0.15
C0 a_n73_n157# a_n33_n245# 0.0289f
C1 a_15_n157# a_n33_n245# 0.0289f
C2 a_15_n157# a_n73_n157# 0.253f
C3 a_15_n157# a_n175_n297# 0.161f
C4 a_n73_n157# a_n175_n297# 0.188f
C5 a_n33_n245# a_n175_n297# 0.322f
.ends

.subckt th09 V09 Vin Vn m1_485_n505# Vp m1_962_372#
XXM0 m1_485_n505# Vn Vin Vn sky130_fd_pr__nfet_01v8_2V6S9N
XXM1 Vin m1_485_n505# Vp Vp Vn sky130_fd_pr__pfet_01v8_XYZSMQ
XXM2 Vp m1_485_n505# Vp m1_962_372# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM3 Vp m1_485_n505# V09 m1_962_372# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM4 Vn V09 m1_485_n505# Vn sky130_fd_pr__nfet_01v8_T8HSQ7
C0 Vin V09 2.77e-19
C1 m1_485_n505# V09 0.104f
C2 Vp V09 0.0743f
C3 V09 m1_962_372# 0.00205f
C4 Vin m1_485_n505# 0.372f
C5 Vin Vp 0.187f
C6 Vp m1_485_n505# 0.372f
C7 V09 Vn 0.00364f
C8 Vin m1_962_372# 0.00821f
C9 m1_485_n505# m1_962_372# 0.0822f
C10 Vp m1_962_372# 0.0579f
C11 Vin Vn 0.0386f
C12 m1_485_n505# Vn 0.0846f
C13 Vp Vn 0.0176f
C14 Vn m1_962_372# 6.71e-21
C15 Vin 0 1.1f
C16 m1_485_n505# 0 1.18f
C17 V09 0 0.27f
C18 Vn 0 0.344f
C19 Vp 0 3.27f
C20 m1_962_372# 0 0.118f
.ends

.subckt sky130_fd_pr__pfet_01v8_HPNF99 a_n33_n147# a_23_n50# a_n81_n50# w_n219_n269#
+ VSUBS
X0 a_23_n50# a_n33_n147# a_n81_n50# w_n219_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.23
C0 w_n219_n269# a_n81_n50# 0.0419f
C1 a_23_n50# a_n81_n50# 0.07f
C2 a_n33_n147# a_n81_n50# 0.00814f
C3 a_23_n50# w_n219_n269# 0.0185f
C4 a_n33_n147# w_n219_n269# 0.173f
C5 a_n33_n147# a_23_n50# 0.00814f
C6 a_23_n50# VSUBS 0.0578f
C7 a_n81_n50# VSUBS 0.0428f
C8 a_n33_n147# VSUBS 0.157f
C9 w_n219_n269# VSUBS 0.779f
.ends

.subckt sky130_fd_pr__nfet_01v8_JZU22M a_n213_n42# a_155_n42# a_n155_n130# a_281_n238#
X0 a_155_n42# a_n155_n130# a_n213_n42# a_281_n238# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.55
C0 a_n155_n130# a_155_n42# 0.0178f
C1 a_n213_n42# a_155_n42# 0.0168f
C2 a_n213_n42# a_n155_n130# 0.0178f
C3 a_155_n42# a_281_n238# 0.0816f
C4 a_n213_n42# a_281_n238# 0.0737f
C5 a_n155_n130# a_281_n238# 0.928f
.ends

.subckt sky130_fd_pr__pfet_01v8_TM5S5A a_n80_n147# a_n138_n50# a_80_n50# w_n276_n269#
+ VSUBS
X0 a_80_n50# a_n80_n147# a_n138_n50# w_n276_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.8
C0 w_n276_n269# a_n138_n50# 0.0231f
C1 a_80_n50# a_n138_n50# 0.0335f
C2 a_n80_n147# a_n138_n50# 0.0141f
C3 a_80_n50# w_n276_n269# 0.0231f
C4 a_n80_n147# w_n276_n269# 0.297f
C5 a_n80_n147# a_80_n50# 0.0141f
C6 a_80_n50# VSUBS 0.0565f
C7 a_n138_n50# VSUBS 0.0565f
C8 a_n80_n147# VSUBS 0.296f
C9 w_n276_n269# VSUBS 1.01f
.ends

.subckt sky130_fd_pr__pfet_01v8_AM8GZ5 w_n526_n261# a_n330_n139# a_330_n42# a_n388_n42#
+ VSUBS
X0 a_330_n42# a_n330_n139# a_n388_n42# w_n526_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.3
C0 w_n526_n261# a_n388_n42# 0.0179f
C1 a_330_n42# a_n388_n42# 0.00853f
C2 a_n330_n139# a_n388_n42# 0.0223f
C3 a_330_n42# w_n526_n261# 0.0408f
C4 a_n330_n139# w_n526_n261# 0.719f
C5 a_n330_n139# a_330_n42# 0.0223f
C6 a_330_n42# VSUBS 0.0435f
C7 a_n388_n42# VSUBS 0.0585f
C8 a_n330_n139# VSUBS 1.13f
C9 w_n526_n261# VSUBS 1.76f
.ends

.subckt sky130_fd_pr__nfet_01v8_H7HSAV a_n73_n250# a_15_n250# a_n33_n338# a_n141_n424#
X0 a_15_n250# a_n33_n338# a_n73_n250# a_n141_n424# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.15
C0 a_n33_n338# a_15_n250# 0.0337f
C1 a_n73_n250# a_15_n250# 0.401f
C2 a_n73_n250# a_n33_n338# 0.0337f
C3 a_15_n250# a_n141_n424# 0.24f
C4 a_n73_n250# a_n141_n424# 0.24f
C5 a_n33_n338# a_n141_n424# 0.327f
.ends

.subckt th14 V14 Vin Vn m1_641_n318# Vp m1_891_419#
XXM0 Vn Vn m1_641_n318# Vp Vn sky130_fd_pr__pfet_01v8_HPNF99
XXM1 m1_641_n318# m1_891_419# Vin Vn sky130_fd_pr__nfet_01v8_JZU22M
XXM2 Vin Vp m1_891_419# Vp Vn sky130_fd_pr__pfet_01v8_TM5S5A
XXM3 Vp m1_891_419# V14 Vp Vn sky130_fd_pr__pfet_01v8_AM8GZ5
XXM4 Vn V14 m1_891_419# Vn sky130_fd_pr__nfet_01v8_H7HSAV
C0 Vin m1_891_419# 0.132f
C1 Vin Vp 0.201f
C2 m1_641_n318# m1_891_419# 0.00289f
C3 Vp m1_641_n318# 0.0629f
C4 V14 m1_891_419# 0.249f
C5 Vp V14 0.082f
C6 Vin m1_641_n318# 0.229f
C7 Vp m1_891_419# 0.227f
C8 Vin V14 0.00516f
C9 m1_891_419# Vn 1.7f
C10 V14 Vn 0.273f
C11 Vp Vn 3.39f
C12 Vin Vn 1.76f
C13 m1_641_n318# Vn 0.313f
.ends

.subckt sky130_fd_pr__nfet_01v8_VGVEGU a_n142_n216# a_n74_n42# a_n33_n130# a_16_n42#
X0 a_16_n42# a_n33_n130# a_n74_n42# a_n142_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.16
C0 a_n74_n42# a_16_n42# 0.0684f
C1 a_n74_n42# a_n33_n130# 0.0191f
C2 a_16_n42# a_n33_n130# 0.0191f
C3 a_16_n42# a_n142_n216# 0.0652f
C4 a_n74_n42# a_n142_n216# 0.0652f
C5 a_n33_n130# a_n142_n216# 0.317f
.ends

.subckt sky130_fd_pr__pfet_01v8_EDPLE3 a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n42# a_15_n42# 0.0699f
C1 w_n211_n261# a_15_n42# 0.0197f
C2 a_n33_n139# a_n73_n42# 0.0192f
C3 a_n33_n139# w_n211_n261# 0.187f
C4 a_n33_n139# a_15_n42# 0.0192f
C5 a_n73_n42# w_n211_n261# 0.0197f
C6 a_15_n42# VSUBS 0.0445f
C7 a_n73_n42# VSUBS 0.0445f
C8 a_n33_n139# VSUBS 0.143f
C9 w_n211_n261# VSUBS 0.749f
.ends

.subckt sky130_fd_pr__pfet_01v8_JM8GTH a_50_n42# w_n246_n261# a_n50_n139# a_n108_n42#
+ VSUBS
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 a_n108_n42# a_50_n42# 0.0391f
C1 w_n246_n261# a_50_n42# 0.0224f
C2 a_n50_n139# a_n108_n42# 0.00909f
C3 a_n50_n139# w_n246_n261# 0.223f
C4 a_n50_n139# a_50_n42# 0.00909f
C5 a_n108_n42# w_n246_n261# 0.0224f
C6 a_50_n42# VSUBS 0.0488f
C7 a_n108_n42# VSUBS 0.0488f
C8 a_n50_n139# VSUBS 0.209f
C9 w_n246_n261# VSUBS 0.88f
.ends

.subckt sky130_fd_pr__nfet_01v8_MYA4RC a_n73_n46# a_n33_n134# a_15_n46# a_n175_n186#
X0 a_15_n46# a_n33_n134# a_n73_n46# a_n175_n186# sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.5 as=0.133 ps=1.5 w=0.46 l=0.15
C0 a_n73_n46# a_15_n46# 0.0763f
C1 a_n73_n46# a_n33_n134# 0.0212f
C2 a_15_n46# a_n33_n134# 0.0212f
C3 a_15_n46# a_n175_n186# 0.0671f
C4 a_n73_n46# a_n175_n186# 0.0756f
C5 a_n33_n134# a_n175_n186# 0.314f
.ends

.subckt th07 Vin V07 Vp m1_808_n892# Vn
XXM0 Vn m1_808_n892# Vin Vn sky130_fd_pr__nfet_01v8_VGVEGU
XXM1 m1_808_n892# Vp Vin Vp Vn sky130_fd_pr__pfet_01v8_EDPLE3
XXM2 V07 Vp m1_808_n892# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM3 V07 m1_808_n892# Vn Vn sky130_fd_pr__nfet_01v8_MYA4RC
C0 m1_808_n892# Vin 0.365f
C1 V07 Vp 0.0569f
C2 m1_808_n892# Vp 0.209f
C3 m1_808_n892# V07 0.112f
C4 Vp Vin 0.157f
C5 V07 Vin 0.00135f
C6 Vin Vn 0.524f
C7 Vp Vn 1.57f
C8 m1_808_n892# Vn 0.596f
C9 V07 Vn 0.276f
.ends

.subckt sky130_fd_pr__pfet_01v8_P28Q2U a_n33_n232# a_15_n135# w_n211_n354# a_n73_n135#
+ VSUBS
X0 a_15_n135# a_n33_n232# a_n73_n135# w_n211_n354# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.28 as=0.391 ps=3.28 w=1.35 l=0.15
C0 a_n73_n135# a_n33_n232# 0.0258f
C1 a_15_n135# a_n33_n232# 0.0258f
C2 a_n73_n135# a_15_n135# 0.218f
C3 w_n211_n354# a_n33_n232# 0.19f
C4 w_n211_n354# a_n73_n135# 0.0279f
C5 w_n211_n354# a_15_n135# 0.0279f
C6 a_15_n135# VSUBS 0.115f
C7 a_n73_n135# VSUBS 0.115f
C8 a_n33_n232# VSUBS 0.146f
C9 w_n211_n354# VSUBS 0.983f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZMY3VB a_n348_n42# a_n290_n130# a_n450_n182# a_290_n42#
X0 a_290_n42# a_n290_n130# a_n348_n42# a_n450_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.9
C0 a_290_n42# a_n348_n42# 0.00961f
C1 a_n290_n130# a_n348_n42# 0.0217f
C2 a_n290_n130# a_290_n42# 0.0217f
C3 a_290_n42# a_n450_n182# 0.076f
C4 a_n348_n42# a_n450_n182# 0.0839f
C5 a_n290_n130# a_n450_n182# 1.6f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n73_n100# a_n33_n197# 0.0236f
C1 a_15_n100# a_n33_n197# 0.0236f
C2 a_n73_n100# a_15_n100# 0.162f
C3 w_n211_n319# a_n33_n197# 0.189f
C4 w_n211_n319# a_n73_n100# 0.0248f
C5 w_n211_n319# a_15_n100# 0.0248f
C6 a_15_n100# VSUBS 0.0885f
C7 a_n73_n100# VSUBS 0.0885f
C8 a_n33_n197# VSUBS 0.145f
C9 w_n211_n319# VSUBS 0.894f
.ends

.subckt sky130_fd_pr__pfet_01v8_WV9GCW a_n158_n42# w_n296_n261# a_n100_n139# a_100_n42#
+ VSUBS
X0 a_100_n42# a_n100_n139# a_n158_n42# w_n296_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1
C0 a_n158_n42# a_n100_n139# 0.0144f
C1 a_100_n42# a_n100_n139# 0.0144f
C2 a_n158_n42# a_100_n42# 0.024f
C3 w_n296_n261# a_n100_n139# 0.346f
C4 w_n296_n261# a_n158_n42# 0.0224f
C5 w_n296_n261# a_100_n42# 0.0224f
C6 a_100_n42# VSUBS 0.0504f
C7 a_n158_n42# VSUBS 0.0504f
C8 a_n100_n139# VSUBS 0.353f
C9 w_n296_n261# VSUBS 1.06f
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n141_240# a_n33_n188# a_15_n100#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n141_240# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_15_n100# a_n73_n100# 0.162f
C1 a_n33_n188# a_n73_n100# 0.0254f
C2 a_n33_n188# a_15_n100# 0.0254f
C3 a_15_n100# a_n141_240# 0.113f
C4 a_n73_n100# a_n141_240# 0.113f
C5 a_n33_n188# a_n141_240# 0.322f
.ends

.subckt th12 Vp V12 Vin m1_529_n42# m1_394_n856# Vn
XXM0 Vn Vn Vp m1_394_n856# Vn sky130_fd_pr__pfet_01v8_P28Q2U
XXM1 m1_529_n42# Vin Vn m1_394_n856# sky130_fd_pr__nfet_01v8_ZMY3VB
XXM2 m1_529_n42# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM3 Vp Vp m1_529_n42# V12 Vn sky130_fd_pr__pfet_01v8_WV9GCW
XXM4 V12 Vn m1_529_n42# Vn sky130_fd_pr__nfet_01v8_648S5X
C0 Vin m1_394_n856# 0.321f
C1 Vn Vp 0.132f
C2 Vn Vin 0.135f
C3 Vp m1_529_n42# 0.322f
C4 Vin m1_529_n42# 0.0965f
C5 Vp Vin 0.238f
C6 m1_394_n856# V12 4.74e-19
C7 Vn V12 0.0234f
C8 Vn m1_394_n856# 0.0338f
C9 m1_529_n42# V12 0.0929f
C10 m1_529_n42# m1_394_n856# 0.0134f
C11 Vn m1_529_n42# 0.254f
C12 Vp V12 0.0454f
C13 Vin V12 0.00205f
C14 Vp m1_394_n856# 0.04f
C15 Vn 0 0.29f
C16 Vp 0 2.88f
C17 m1_529_n42# 0 0.861f
C18 V12 0 0.359f
C19 Vin 0 1.9f
C20 m1_394_n856# 0 0.215f
.ends

.subckt sky130_fd_pr__nfet_01v8_Q7AWK3 a_n180_n340# a_20_n200# a_n78_n200# a_n33_n288#
X0 a_20_n200# a_n33_n288# a_n78_n200# a_n180_n340# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
C0 a_20_n200# a_n78_n200# 0.288f
C1 a_n33_n288# a_n78_n200# 0.024f
C2 a_n33_n288# a_20_n200# 0.024f
C3 a_20_n200# a_n180_n340# 0.202f
C4 a_n78_n200# a_n180_n340# 0.237f
C5 a_n33_n288# a_n180_n340# 0.325f
.ends

.subckt sky130_fd_pr__pfet_01v8_EXJYQP w_n359_n261# a_n163_n139# a_n221_n42# a_163_n42#
+ VSUBS
X0 a_163_n42# a_n163_n139# a_n221_n42# w_n359_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.63
C0 a_n221_n42# a_n163_n139# 0.0182f
C1 a_163_n42# a_n163_n139# 0.0182f
C2 a_163_n42# a_n221_n42# 0.0161f
C3 w_n359_n261# a_n163_n139# 0.413f
C4 w_n359_n261# a_n221_n42# 0.0179f
C5 w_n359_n261# a_163_n42# 0.0408f
C6 a_163_n42# VSUBS 0.041f
C7 a_n221_n42# VSUBS 0.056f
C8 a_n163_n139# VSUBS 0.584f
C9 w_n359_n261# VSUBS 1.24f
.ends

.subckt sky130_fd_pr__pfet_01v8_HJHF6N a_n170_n50# w_n308_n269# a_n112_n147# a_112_n50#
+ VSUBS
X0 a_112_n50# a_n112_n147# a_n170_n50# w_n308_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1.12
C0 a_n170_n50# a_n112_n147# 0.0172f
C1 a_112_n50# a_n112_n147# 0.0172f
C2 a_112_n50# a_n170_n50# 0.0259f
C3 w_n308_n269# a_n112_n147# 0.378f
C4 w_n308_n269# a_n170_n50# 0.0232f
C5 w_n308_n269# a_112_n50# 0.0232f
C6 a_112_n50# VSUBS 0.0577f
C7 a_n170_n50# VSUBS 0.0577f
C8 a_n112_n147# VSUBS 0.389f
C9 w_n308_n269# VSUBS 1.14f
.ends

.subckt sky130_fd_pr__nfet_01v8_N39H2X a_n76_n100# a_n33_n188# a_18_n100# a_144_n240#
X0 a_18_n100# a_n33_n188# a_n76_n100# a_144_n240# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.18
C0 a_18_n100# a_n76_n100# 0.152f
C1 a_n33_n188# a_n76_n100# 0.0205f
C2 a_n33_n188# a_18_n100# 0.0205f
C3 a_18_n100# a_144_n240# 0.133f
C4 a_n76_n100# a_144_n240# 0.115f
C5 a_n33_n188# a_144_n240# 0.32f
.ends

.subckt th05 Vp V05 Vin m1_752_n794# Vn
XXM0 Vn m1_752_n794# Vn Vin sky130_fd_pr__nfet_01v8_Q7AWK3
XXM1 Vp Vin m1_752_n794# Vp Vn sky130_fd_pr__pfet_01v8_EXJYQP
XXM2 Vp Vp m1_752_n794# V05 Vn sky130_fd_pr__pfet_01v8_HJHF6N
XXM3 Vn m1_752_n794# V05 Vn sky130_fd_pr__nfet_01v8_N39H2X
C0 V05 m1_752_n794# 0.0855f
C1 V05 Vp 0.0548f
C2 V05 Vin 0.00406f
C3 Vp m1_752_n794# 0.198f
C4 Vin m1_752_n794# 0.2f
C5 Vin Vp 0.139f
C6 V05 Vn 0.0364f
C7 m1_752_n794# Vn 0.136f
C8 Vp Vn 0.0115f
C9 Vin Vn 0.041f
C10 m1_752_n794# 0 0.788f
C11 Vp 0 2.28f
C12 V05 0 0.314f
C13 Vin 0 0.905f
C14 Vn 0 0.547f
.ends

.subckt sky130_fd_pr__nfet_01v8_4L9AWD a_n206_n182# a_n46_n130# a_n104_n42# a_46_n42#
X0 a_46_n42# a_n46_n130# a_n104_n42# a_n206_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.46
C0 a_46_n42# a_n46_n130# 0.00852f
C1 a_n104_n42# a_n46_n130# 0.00852f
C2 a_n104_n42# a_46_n42# 0.0412f
C3 a_46_n42# a_n206_n182# 0.0705f
C4 a_n104_n42# a_n206_n182# 0.0784f
C5 a_n46_n130# a_n206_n182# 0.388f
.ends

.subckt sky130_fd_pr__pfet_01v8_EZD9Q7 w_n224_n261# a_28_n42# a_n33_n139# a_n86_n42#
+ VSUBS
X0 a_28_n42# a_n33_n139# a_n86_n42# w_n224_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.28
C0 a_n86_n42# a_28_n42# 0.0541f
C1 a_n33_n139# a_28_n42# 0.00625f
C2 a_n86_n42# w_n224_n261# 0.0224f
C3 a_n33_n139# w_n224_n261# 0.183f
C4 w_n224_n261# a_28_n42# 0.0224f
C5 a_n33_n139# a_n86_n42# 0.00625f
C6 a_28_n42# VSUBS 0.0479f
C7 a_n86_n42# VSUBS 0.0479f
C8 a_n33_n139# VSUBS 0.155f
C9 w_n224_n261# VSUBS 0.799f
.ends

.subckt sky130_fd_pr__pfet_01v8_M479BZ a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n42# a_15_n42# 0.0699f
C1 a_n33_n139# a_15_n42# 0.0192f
C2 a_n73_n42# w_n211_n261# 0.016f
C3 a_n33_n139# w_n211_n261# 0.182f
C4 w_n211_n261# a_15_n42# 0.0389f
C5 a_n33_n139# a_n73_n42# 0.0192f
C6 a_15_n42# VSUBS 0.0328f
C7 a_n73_n42# VSUBS 0.0478f
C8 a_n33_n139# VSUBS 0.145f
C9 w_n211_n261# VSUBS 0.785f
.ends

.subckt sky130_fd_pr__nfet_01v8_4BNSKG a_n144_n216# a_18_n42# a_n33_n130# a_n76_n42#
X0 a_18_n42# a_n33_n130# a_n76_n42# a_n144_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.18
C0 a_18_n42# a_n33_n130# 0.0154f
C1 a_n76_n42# a_n33_n130# 0.0154f
C2 a_n76_n42# a_18_n42# 0.0655f
C3 a_18_n42# a_n144_n216# 0.0668f
C4 a_n76_n42# a_n144_n216# 0.0668f
C5 a_n33_n130# a_n144_n216# 0.319f
.ends

.subckt th10 Vp V10 Vin Vn m1_502_n495# m1_536_174#
XXM0 m1_502_n495# Vn Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vn Vin m1_536_174# m1_502_n495# sky130_fd_pr__nfet_01v8_4L9AWD
XXM2 Vp m1_536_174# Vin Vp Vn sky130_fd_pr__pfet_01v8_EZD9Q7
XXM3 Vp Vp m1_536_174# V10 Vn sky130_fd_pr__pfet_01v8_M479BZ
XXM4 Vn V10 m1_536_174# Vn sky130_fd_pr__nfet_01v8_4BNSKG
C0 V10 Vp 0.0702f
C1 Vn m1_502_n495# 0.0348f
C2 Vin m1_502_n495# 0.0207f
C3 m1_536_174# m1_502_n495# 0.00612f
C4 Vp m1_502_n495# 0.0256f
C5 Vn Vin 0.114f
C6 V10 m1_502_n495# 0.042f
C7 Vn m1_536_174# 0.233f
C8 m1_536_174# Vin 0.0971f
C9 Vn Vp 0.102f
C10 Vp Vin 0.175f
C11 m1_536_174# Vp 0.172f
C12 V10 Vn 0.0577f
C13 V10 Vin 0.0187f
C14 V10 m1_536_174# 0.177f
C15 Vin 0 0.664f
C16 m1_536_174# 0 0.825f
C17 Vp 0 2.17f
C18 V10 0 0.249f
C19 Vn 0 0.463f
C20 m1_502_n495# 0 0.146f
.ends

.subckt sky130_fd_pr__nfet_01v8_X33H33 a_n73_n110# a_n175_n250# a_n33_n198# a_15_n110#
X0 a_15_n110# a_n33_n198# a_n73_n110# a_n175_n250# sky130_fd_pr__nfet_01v8 ad=0.319 pd=2.78 as=0.319 ps=2.78 w=1.1 l=0.15
C0 a_15_n110# a_n33_n198# 0.0261f
C1 a_15_n110# a_n73_n110# 0.178f
C2 a_n73_n110# a_n33_n198# 0.0261f
C3 a_15_n110# a_n175_n250# 0.121f
C4 a_n73_n110# a_n175_n250# 0.141f
C5 a_n33_n198# a_n175_n250# 0.32f
.ends

.subckt sky130_fd_pr__pfet_01v8_AMA9E4 a_n194_n44# a_n136_n141# w_n332_n263# a_136_n44#
+ VSUBS
X0 a_136_n44# a_n136_n141# a_n194_n44# w_n332_n263# sky130_fd_pr__pfet_01v8 ad=0.128 pd=1.46 as=0.128 ps=1.46 w=0.44 l=1.36
C0 a_136_n44# a_n136_n141# 0.0174f
C1 a_n194_n44# w_n332_n263# 0.0226f
C2 a_n194_n44# a_n136_n141# 0.0174f
C3 a_n194_n44# a_136_n44# 0.0196f
C4 a_n136_n141# w_n332_n263# 0.434f
C5 a_136_n44# w_n332_n263# 0.0226f
C6 a_136_n44# VSUBS 0.0532f
C7 a_n194_n44# VSUBS 0.0532f
C8 a_n136_n141# VSUBS 0.457f
C9 w_n332_n263# VSUBS 1.2f
.ends

.subckt sky130_fd_pr__pfet_01v8_8DZSNJ a_n74_n100# a_16_n100# w_n212_n319# a_n33_n197#
+ VSUBS
X0 a_16_n100# a_n33_n197# a_n74_n100# w_n212_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.16
C0 a_16_n100# a_n33_n197# 0.0223f
C1 a_n74_n100# w_n212_n319# 0.0252f
C2 a_n74_n100# a_n33_n197# 0.0223f
C3 a_n74_n100# a_16_n100# 0.159f
C4 a_n33_n197# w_n212_n319# 0.189f
C5 a_16_n100# w_n212_n319# 0.0252f
C6 a_16_n100# VSUBS 0.089f
C7 a_n74_n100# VSUBS 0.089f
C8 a_n33_n197# VSUBS 0.146f
C9 w_n212_n319# VSUBS 0.899f
.ends

.subckt th03 V03 Vin Vp m1_890_n844# m1_638_n591# Vn
XXM0 Vn Vn Vin m1_890_n844# sky130_fd_pr__nfet_01v8_X33H33
XXM1 m1_638_n591# Vin Vp m1_890_n844# Vn sky130_fd_pr__pfet_01v8_AMA9E4
XXM2 Vp Vn Vp m1_638_n591# sky130_fd_pr__nfet_01v8_LH5FDA
XXM3 Vp V03 Vp m1_890_n844# Vn sky130_fd_pr__pfet_01v8_8DZSNJ
XXM4 m1_890_n844# Vn Vn V03 sky130_fd_pr__nfet_01v8_LH5FDA
C0 Vn m1_890_n844# 0.183f
C1 Vin Vp 0.313f
C2 V03 Vp 0.0492f
C3 Vin V03 0.0036f
C4 Vn m1_638_n591# 0.0097f
C5 m1_890_n844# Vp 0.459f
C6 Vin m1_890_n844# 0.188f
C7 m1_890_n844# V03 0.129f
C8 m1_638_n591# Vp 0.169f
C9 Vin m1_638_n591# 0.0439f
C10 m1_890_n844# m1_638_n591# 0.0187f
C11 Vn Vp 0.023f
C12 Vn Vin 0.105f
C13 Vn V03 0.0337f
C14 Vp 0 3.07f
C15 V03 0 0.308f
C16 Vn 0 0.446f
C17 m1_890_n844# 0 1.05f
C18 m1_638_n591# 0 0.224f
C19 Vin 0 0.924f
.ends

.subckt sky130_fd_pr__nfet_01v8_SHU4BF a_n73_n353# a_n141_493# a_15_n353# a_n33_n441#
X0 a_15_n353# a_n33_n441# a_n73_n353# a_n141_493# sky130_fd_pr__nfet_01v8 ad=1.02 pd=7.64 as=1.02 ps=7.64 w=3.53 l=0.15
C0 a_15_n353# a_n73_n353# 0.564f
C1 a_n33_n441# a_15_n353# 0.0384f
C2 a_n33_n441# a_n73_n353# 0.0384f
C3 a_15_n353# a_n141_493# 0.327f
C4 a_n73_n353# a_n141_493# 0.327f
C5 a_n33_n441# a_n141_493# 0.329f
.ends

.subckt sky130_fd_pr__pfet_01v8_HE9GT9 a_n408_n42# a_350_n42# w_n546_n261# a_n350_n139#
+ VSUBS
X0 a_350_n42# a_n350_n139# a_n408_n42# w_n546_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 a_n408_n42# a_350_n42# 0.00807f
C1 a_350_n42# a_n350_n139# 0.0226f
C2 a_n408_n42# a_n350_n139# 0.0226f
C3 w_n546_n261# a_350_n42# 0.0179f
C4 w_n546_n261# a_n408_n42# 0.0408f
C5 w_n546_n261# a_n350_n139# 0.756f
C6 a_350_n42# VSUBS 0.0587f
C7 a_n408_n42# VSUBS 0.0437f
C8 a_n350_n139# VSUBS 1.19f
C9 w_n546_n261# VSUBS 1.83f
.ends

.subckt sky130_fd_pr__nfet_01v8_LHD8GA a_n408_n42# a_350_n42# a_n350_n130# a_n510_n182#
X0 a_350_n42# a_n350_n130# a_n408_n42# a_n510_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 a_350_n42# a_n408_n42# 0.00807f
C1 a_n350_n130# a_350_n42# 0.0226f
C2 a_n350_n130# a_n408_n42# 0.0226f
C3 a_350_n42# a_n510_n182# 0.0766f
C4 a_n408_n42# a_n510_n182# 0.0845f
C5 a_n350_n130# a_n510_n182# 1.9f
.ends

.subckt th01 Vp Vin V01 m1_991_n1219# Vn m1_571_n501#
XXM0 Vn Vn m1_991_n1219# Vin sky130_fd_pr__nfet_01v8_SHU4BF
XXM1 m1_571_n501# m1_991_n1219# Vp Vin Vn sky130_fd_pr__pfet_01v8_HE9GT9
XXM2 Vp m1_571_n501# Vp Vn sky130_fd_pr__nfet_01v8_LHD8GA
XXM3 Vp Vp V01 m1_991_n1219# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_991_n1219# Vn V01 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 Vn V01 0.0149f
C1 Vp V01 0.0684f
C2 m1_571_n501# Vin 0.274f
C3 m1_991_n1219# Vin 0.208f
C4 Vin Vn 0.0582f
C5 Vp Vin 0.354f
C6 m1_571_n501# m1_991_n1219# 0.0899f
C7 m1_571_n501# Vn 2.57e-20
C8 Vp m1_571_n501# 0.32f
C9 m1_991_n1219# Vn 0.0569f
C10 Vp m1_991_n1219# 0.423f
C11 Vin V01 0.00412f
C12 Vp Vn 0.0233f
C13 m1_571_n501# V01 2.16e-20
C14 m1_991_n1219# V01 0.0901f
C15 Vn 0 0.633f
C16 m1_991_n1219# 0 1.24f
C17 V01 0 0.373f
C18 Vp 0 4.41f
C19 m1_571_n501# 0 0.194f
C20 Vin 0 1.87f
.ends

.subckt sky130_fd_pr__pfet_01v8_MWHFPY a_n73_n63# a_n33_n160# w_n211_n282# a_15_n63#
+ VSUBS
X0 a_15_n63# a_n33_n160# a_n73_n63# w_n211_n282# sky130_fd_pr__pfet_01v8 ad=0.183 pd=1.84 as=0.183 ps=1.84 w=0.63 l=0.15
C0 w_n211_n282# a_n33_n160# 0.237f
C1 a_n73_n63# w_n211_n282# 0.0591f
C2 a_n73_n63# a_n33_n160# 0.021f
C3 a_15_n63# w_n211_n282# 0.0591f
C4 a_15_n63# a_n33_n160# 0.021f
C5 a_15_n63# a_n73_n63# 0.103f
C6 a_15_n63# VSUBS 0.0348f
C7 a_n73_n63# VSUBS 0.0348f
C8 a_n33_n160# VSUBS 0.116f
C9 w_n211_n282# VSUBS 1.1f
.ends

.subckt sky130_fd_pr__nfet_01v8_DPSGWY a_350_n100# a_n408_n100# a_n350_n188# a_n510_n274#
X0 a_350_n100# a_n350_n188# a_n408_n100# a_n510_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3.5
C0 a_n350_n188# a_n408_n100# 0.0439f
C1 a_350_n100# a_n350_n188# 0.0439f
C2 a_350_n100# a_n408_n100# 0.0188f
C3 a_350_n100# a_n510_n274# 0.159f
C4 a_n408_n100# a_n510_n274# 0.159f
C5 a_n350_n188# a_n510_n274# 2.13f
.ends

.subckt preamp Vp Vin Vpamp Vn
XXM0 Vn Vin Vp Vpamp Vn sky130_fd_pr__pfet_01v8_MWHFPY
XXM1 Vpamp Vp Vin Vn sky130_fd_pr__nfet_01v8_DPSGWY
C0 Vp Vin 0.324f
C1 Vp Vn 0.297f
C2 Vpamp Vin 0.0777f
C3 Vpamp Vn 0.047f
C4 Vp Vpamp 0.0552f
C5 Vin Vn 0.29f
C6 Vn 0 0.193f
C7 Vpamp 0 0.444f
C8 Vp 0 1.53f
C9 Vin 0 2.21f
.ends

.subckt sky130_fd_pr__pfet_01v8_LDQF7K a_n33_n147# a_29_n50# a_n87_n50# w_n225_n269#
+ VSUBS
X0 a_29_n50# a_n33_n147# a_n87_n50# w_n225_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.29
C0 a_29_n50# a_n33_n147# 0.00691f
C1 w_n225_n269# a_n87_n50# 0.0457f
C2 a_n33_n147# w_n225_n269# 0.176f
C3 a_29_n50# w_n225_n269# 0.0186f
C4 a_n33_n147# a_n87_n50# 0.00691f
C5 a_29_n50# a_n87_n50# 0.0628f
C6 a_29_n50# VSUBS 0.0581f
C7 a_n87_n50# VSUBS 0.0403f
C8 a_n33_n147# VSUBS 0.158f
C9 w_n225_n269# VSUBS 0.854f
.ends

.subckt sky130_fd_pr__nfet_01v8_HZA4VB a_326_n230# a_n200_n130# a_200_n42# li_n360_158#
+ a_n258_n42#
X0 a_200_n42# a_n200_n130# a_n258_n42# a_326_n230# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_n200_n130# a_200_n42# 0.0196f
C1 a_n258_n42# a_n200_n130# 0.0196f
C2 a_n258_n42# a_200_n42# 0.0134f
C3 li_n360_158# a_326_n230# 0.0244f
C4 a_200_n42# a_326_n230# 0.0748f
C5 a_n258_n42# a_326_n230# 0.0746f
C6 a_n200_n130# a_326_n230# 1.15f
.ends

.subckt sky130_fd_pr__pfet_01v8_GEY2B5 w_n275_n270# a_n137_n51# a_79_n51# a_n79_n148#
+ VSUBS
X0 a_79_n51# a_n79_n148# a_n137_n51# w_n275_n270# sky130_fd_pr__pfet_01v8 ad=0.148 pd=1.6 as=0.148 ps=1.6 w=0.51 l=0.79
C0 a_79_n51# a_n79_n148# 0.0141f
C1 w_n275_n270# a_n137_n51# 0.0232f
C2 a_n79_n148# w_n275_n270# 0.294f
C3 a_79_n51# w_n275_n270# 0.0232f
C4 a_n79_n148# a_n137_n51# 0.0141f
C5 a_79_n51# a_n137_n51# 0.0345f
C6 a_79_n51# VSUBS 0.0573f
C7 a_n137_n51# VSUBS 0.0573f
C8 a_n79_n148# VSUBS 0.294f
C9 w_n275_n270# VSUBS 1.01f
.ends

.subckt sky130_fd_pr__pfet_01v8_KQKFM4 w_n526_n261# a_n330_n139# a_330_n42# a_n388_n42#
+ VSUBS
X0 a_330_n42# a_n330_n139# a_n388_n42# w_n526_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.3
C0 a_330_n42# a_n330_n139# 0.0223f
C1 w_n526_n261# a_n388_n42# 0.0224f
C2 a_n330_n139# w_n526_n261# 0.911f
C3 a_330_n42# w_n526_n261# 0.0224f
C4 a_n330_n139# a_n388_n42# 0.0223f
C5 a_330_n42# a_n388_n42# 0.00853f
C6 a_330_n42# VSUBS 0.0545f
C7 a_n388_n42# VSUBS 0.0545f
C8 a_n330_n139# VSUBS 1.02f
C9 w_n526_n261# VSUBS 1.89f
.ends

.subckt sky130_fd_pr__nfet_01v8_5NW376 a_n73_n251# a_n141_391# a_15_n251# a_n33_n339#
X0 a_15_n251# a_n33_n339# a_n73_n251# a_n141_391# sky130_fd_pr__nfet_01v8 ad=0.728 pd=5.6 as=0.728 ps=5.6 w=2.51 l=0.15
C0 a_n33_n339# a_15_n251# 0.0337f
C1 a_n73_n251# a_n33_n339# 0.0337f
C2 a_n73_n251# a_15_n251# 0.402f
C3 a_15_n251# a_n141_391# 0.241f
C4 a_n73_n251# a_n141_391# 0.241f
C5 a_n33_n339# a_n141_391# 0.327f
.ends

.subckt th15 V15 Vin m1_597_n912# Vp m1_849_n157# Vn
XXM0 Vn Vn m1_597_n912# Vp Vn sky130_fd_pr__pfet_01v8_LDQF7K
XXM1 Vn Vin m1_849_n157# Vn m1_597_n912# sky130_fd_pr__nfet_01v8_HZA4VB
XXM2 Vp Vp m1_849_n157# Vin Vn sky130_fd_pr__pfet_01v8_GEY2B5
XXM3 Vp m1_849_n157# V15 Vp Vn sky130_fd_pr__pfet_01v8_KQKFM4
XXM4 Vn Vn V15 m1_849_n157# sky130_fd_pr__nfet_01v8_5NW376
C0 V15 Vp 0.0762f
C1 V15 m1_849_n157# 0.202f
C2 m1_597_n912# Vp 0.0557f
C3 m1_597_n912# m1_849_n157# 0.00715f
C4 Vp m1_849_n157# 0.226f
C5 V15 Vn 2.72e-19
C6 m1_597_n912# Vn 0.175f
C7 Vin V15 0.00573f
C8 Vp Vn 0.0678f
C9 Vin m1_597_n912# 0.211f
C10 m1_849_n157# Vn 0.171f
C11 Vin Vp 0.166f
C12 Vin m1_849_n157# 0.0977f
C13 Vin Vn 0.38f
C14 V15 0 0.332f
C15 Vn 0 0.276f
C16 m1_849_n157# 0 1.28f
C17 Vp 0 3.52f
C18 Vin 0 1.58f
C19 m1_597_n912# 0 0.19f
.ends

.subckt sky130_fd_pr__nfet_01v8_JSJ4VK a_113_n42# a_n239_n216# a_n171_n42# a_n113_n130#
X0 a_113_n42# a_n113_n130# a_n171_n42# a_n239_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.13
C0 a_n171_n42# a_113_n42# 0.0218f
C1 a_n113_n130# a_113_n42# 0.0154f
C2 a_n113_n130# a_n171_n42# 0.0154f
C3 a_113_n42# a_n239_n216# 0.0734f
C4 a_n171_n42# a_n239_n216# 0.0734f
C5 a_n113_n130# a_n239_n216# 0.746f
.ends

.subckt sky130_fd_pr__pfet_01v8_EVXEQ2 a_16_n67# a_n33_n164# a_n74_n67# w_n212_n286#
+ VSUBS
X0 a_16_n67# a_n33_n164# a_n74_n67# w_n212_n286# sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.92 as=0.194 ps=1.92 w=0.67 l=0.16
C0 a_n33_n164# a_n74_n67# 0.0198f
C1 w_n212_n286# a_16_n67# 0.0544f
C2 a_n74_n67# a_16_n67# 0.107f
C3 a_n33_n164# a_16_n67# 0.0198f
C4 w_n212_n286# a_n74_n67# 0.0184f
C5 w_n212_n286# a_n33_n164# 0.183f
C6 a_16_n67# VSUBS 0.0435f
C7 a_n74_n67# VSUBS 0.0673f
C8 a_n33_n164# VSUBS 0.147f
C9 w_n212_n286# VSUBS 0.864f
.ends

.subckt sky130_fd_pr__pfet_01v8_BBE9QE w_n244_n262# a_n106_n43# a_48_n43# a_n48_n140#
+ VSUBS
X0 a_48_n43# a_n48_n140# a_n106_n43# w_n244_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.48
C0 a_n48_n140# a_n106_n43# 0.00893f
C1 w_n244_n262# a_48_n43# 0.0225f
C2 a_n106_n43# a_48_n43# 0.041f
C3 a_n48_n140# a_48_n43# 0.00893f
C4 w_n244_n262# a_n106_n43# 0.0225f
C5 w_n244_n262# a_n48_n140# 0.218f
C6 a_48_n43# VSUBS 0.0495f
C7 a_n106_n43# VSUBS 0.0495f
C8 a_n48_n140# VSUBS 0.203f
C9 w_n244_n262# VSUBS 0.876f
.ends

.subckt sky130_fd_pr__nfet_01v8_NCP4B2 a_n73_n47# a_n141_n221# a_n33_n135# a_15_n47#
X0 a_15_n47# a_n33_n135# a_n73_n47# a_n141_n221# sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.52 as=0.136 ps=1.52 w=0.47 l=0.15
C0 a_n73_n47# a_15_n47# 0.0779f
C1 a_n33_n135# a_15_n47# 0.0213f
C2 a_n33_n135# a_n73_n47# 0.0213f
C3 a_15_n47# a_n141_n221# 0.0686f
C4 a_n73_n47# a_n141_n221# 0.0686f
C5 a_n33_n135# a_n141_n221# 0.317f
.ends

.subckt th08 Vin V08 m1_477_n803# Vp Vn
XXM0 Vn Vn m1_477_n803# Vin sky130_fd_pr__nfet_01v8_JSJ4VK
XXM1 Vp Vin m1_477_n803# Vp Vn sky130_fd_pr__pfet_01v8_EVXEQ2
XXM2 Vp Vp V08 m1_477_n803# Vn sky130_fd_pr__pfet_01v8_BBE9QE
XXM3 Vn Vn m1_477_n803# V08 sky130_fd_pr__nfet_01v8_NCP4B2
C0 m1_477_n803# Vin 0.356f
C1 Vp V08 0.0461f
C2 m1_477_n803# Vp 0.154f
C3 Vin Vp 0.0933f
C4 m1_477_n803# V08 0.108f
C5 Vin V08 0.00163f
C6 m1_477_n803# Vn 0.656f
C7 Vin Vn 1.02f
C8 V08 Vn 0.271f
C9 Vp Vn 1.66f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFRTVB a_n410_n216# a_n250_n130# a_n308_n42# a_250_n42#
X0 a_250_n42# a_n250_n130# a_n308_n42# a_n410_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.5
C0 a_n308_n42# a_n250_n130# 0.0209f
C1 a_250_n42# a_n250_n130# 0.0209f
C2 a_250_n42# a_n308_n42# 0.011f
C3 a_250_n42# a_n410_n216# 0.0852f
C4 a_n308_n42# a_n410_n216# 0.0853f
C5 a_n250_n130# a_n410_n216# 1.48f
.ends

.subckt sky130_fd_pr__pfet_01v8_XQZLDL a_15_n240# w_n211_n459# a_n73_n240# a_n33_n337#
+ VSUBS
X0 a_15_n240# a_n33_n337# a_n73_n240# w_n211_n459# sky130_fd_pr__pfet_01v8 ad=0.696 pd=5.38 as=0.696 ps=5.38 w=2.4 l=0.15
C0 a_n33_n337# w_n211_n459# 0.206f
C1 a_n73_n240# a_15_n240# 0.385f
C2 a_15_n240# w_n211_n459# 0.163f
C3 a_n33_n337# a_15_n240# 0.0313f
C4 a_n73_n240# w_n211_n459# 0.0371f
C5 a_n73_n240# a_n33_n337# 0.0313f
C6 a_15_n240# VSUBS 0.11f
C7 a_n73_n240# VSUBS 0.195f
C8 a_n33_n337# VSUBS 0.139f
C9 w_n211_n459# VSUBS 1.47f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GC6 a_200_n42# w_n396_n261# a_n200_n139# a_n258_n42#
+ VSUBS
X0 a_200_n42# a_n200_n139# a_n258_n42# w_n396_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_n200_n139# w_n396_n261# 0.73f
C1 a_n258_n42# a_200_n42# 0.0134f
C2 a_200_n42# w_n396_n261# 0.0498f
C3 a_n200_n139# a_200_n42# 0.0196f
C4 a_n258_n42# w_n396_n261# 0.0269f
C5 a_n258_n42# a_n200_n139# 0.0196f
C6 a_200_n42# VSUBS 0.0338f
C7 a_n258_n42# VSUBS 0.0488f
C8 a_n200_n139# VSUBS 0.563f
C9 w_n396_n261# VSUBS 1.69f
.ends

.subckt sky130_fd_pr__nfet_01v8_ATLS57 a_15_n200# a_n73_n200# a_n33_n288# a_n141_n374#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n141_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n73_n200# a_n33_n288# 0.0312f
C1 a_15_n200# a_n33_n288# 0.0312f
C2 a_15_n200# a_n73_n200# 0.321f
C3 a_15_n200# a_n141_n374# 0.233f
C4 a_n73_n200# a_n141_n374# 0.199f
C5 a_n33_n288# a_n141_n374# 0.341f
.ends

.subckt th13 V13 Vin m1_831_275# Vn Vp m1_559_n458#
XXM0 Vn m1_559_n458# Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vn Vin m1_559_n458# m1_831_275# sky130_fd_pr__nfet_01v8_ZFRTVB
XXM2 Vp Vp m1_831_275# Vin Vn sky130_fd_pr__pfet_01v8_XQZLDL
XXM3 V13 Vp m1_831_275# Vp Vn sky130_fd_pr__pfet_01v8_VZ9GC6
XXM4 V13 Vn m1_831_275# Vn sky130_fd_pr__nfet_01v8_ATLS57
C0 Vn m1_559_n458# 0.152f
C1 Vn Vin 0.347f
C2 Vn Vp 0.206f
C3 m1_559_n458# m1_831_275# 0.0183f
C4 Vin m1_831_275# 0.197f
C5 m1_831_275# Vp 0.215f
C6 V13 Vn 0.0706f
C7 V13 m1_831_275# 0.184f
C8 m1_559_n458# Vin 0.181f
C9 m1_559_n458# Vp 0.0628f
C10 Vn m1_831_275# 0.232f
C11 Vin Vp 0.176f
C12 V13 Vin 0.0076f
C13 V13 Vp 0.135f
C14 m1_831_275# 0 1.05f
C15 Vin 0 1.79f
C16 V13 0 0.365f
C17 Vn 0 0.117f
C18 Vp 0 3.98f
C19 m1_559_n458# 0 0.286f
.ends

.subckt sky130_fd_pr__nfet_01v8_DD6SHA a_n33_n130# a_15_n42# a_n175_n182# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_15_n42# a_n73_n42# 0.0699f
C1 a_n73_n42# a_n33_n130# 0.0209f
C2 a_15_n42# a_n33_n130# 0.0209f
C3 a_15_n42# a_n175_n182# 0.0637f
C4 a_n73_n42# a_n175_n182# 0.0716f
C5 a_n33_n130# a_n175_n182# 0.314f
.ends

.subckt sky130_fd_pr__pfet_01v8_7DPLFP w_n245_n261# a_n107_n42# a_n49_n139# a_49_n42#
+ VSUBS
X0 a_49_n42# a_n49_n139# a_n107_n42# w_n245_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.49
C0 a_n107_n42# a_n49_n139# 0.00895f
C1 a_n49_n139# w_n245_n261# 0.221f
C2 a_n107_n42# w_n245_n261# 0.0224f
C3 a_n107_n42# a_49_n42# 0.0396f
C4 a_n49_n139# a_49_n42# 0.00895f
C5 a_49_n42# w_n245_n261# 0.0224f
C6 a_49_n42# VSUBS 0.0487f
C7 a_n107_n42# VSUBS 0.0487f
C8 a_n49_n139# VSUBS 0.206f
C9 w_n245_n261# VSUBS 0.876f
.ends

.subckt sky130_fd_pr__pfet_01v8_MDPZBH a_n102_n42# a_44_n42# a_n44_n139# w_n240_n261#
+ VSUBS
X0 a_44_n42# a_n44_n139# a_n102_n42# w_n240_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.44
C0 a_n102_n42# a_n44_n139# 0.00823f
C1 a_n44_n139# w_n240_n261# 0.208f
C2 a_n102_n42# w_n240_n261# 0.0224f
C3 a_n102_n42# a_44_n42# 0.0423f
C4 a_n44_n139# a_44_n42# 0.00823f
C5 a_44_n42# w_n240_n261# 0.0224f
C6 a_44_n42# VSUBS 0.0485f
C7 a_n102_n42# VSUBS 0.0485f
C8 a_n44_n139# VSUBS 0.191f
C9 w_n240_n261# VSUBS 0.858f
.ends

.subckt th06 Vp Vin V06 Vn m1_904_n796#
XXM0 Vin m1_904_n796# Vn Vn sky130_fd_pr__nfet_01v8_DD6SHA
XXM1 Vp Vp Vin m1_904_n796# Vn sky130_fd_pr__pfet_01v8_7DPLFP
XXM2 Vp V06 m1_904_n796# Vp Vn sky130_fd_pr__pfet_01v8_MDPZBH
XXM3 Vn m1_904_n796# V06 Vn sky130_fd_pr__nfet_01v8_MYA4RC
C0 V06 Vn 0.00141f
C1 Vin m1_904_n796# 0.203f
C2 Vp Vn 0.0214f
C3 V06 Vp 0.06f
C4 m1_904_n796# Vn 0.0382f
C5 Vin Vn 0.0188f
C6 V06 m1_904_n796# 0.157f
C7 Vp m1_904_n796# 0.197f
C8 Vin Vp 0.113f
C9 Vp 0 1.69f
C10 V06 0 0.217f
C11 Vn 0 0.286f
C12 m1_904_n796# 0 0.495f
C13 Vin 0 0.524f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGAKDL a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
+ VSUBS
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n33_n297# a_n73_n200# 0.0293f
C1 a_n33_n297# w_n211_n419# 0.191f
C2 a_15_n200# a_n73_n200# 0.321f
C3 a_15_n200# w_n211_n419# 0.0336f
C4 w_n211_n419# a_n73_n200# 0.0336f
C5 a_n33_n297# a_15_n200# 0.0293f
C6 a_15_n200# VSUBS 0.164f
C7 a_n73_n200# VSUBS 0.164f
C8 a_n33_n297# VSUBS 0.147f
C9 w_n211_n419# VSUBS 1.14f
.ends

.subckt sky130_fd_pr__nfet_01v8_4X3CDA a_n306_n216# a_n180_n130# a_n238_n42# a_180_n42#
X0 a_180_n42# a_n180_n130# a_n238_n42# a_n306_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.8
C0 a_n238_n42# a_180_n42# 0.0147f
C1 a_n238_n42# a_n180_n130# 0.0189f
C2 a_n180_n130# a_180_n42# 0.0189f
C3 a_180_n42# a_n306_n216# 0.075f
C4 a_n238_n42# a_n306_n216# 0.075f
C5 a_n180_n130# a_n306_n216# 1.1f
.ends

.subckt sky130_fd_pr__pfet_01v8_MWB9BZ a_15_n43# w_n211_n262# a_n73_n43# a_n33_n140#
+ VSUBS
X0 a_15_n43# a_n33_n140# a_n73_n43# w_n211_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.15
C0 a_n33_n140# a_n73_n43# 0.0193f
C1 a_n33_n140# w_n211_n262# 0.187f
C2 a_15_n43# a_n73_n43# 0.0715f
C3 a_15_n43# w_n211_n262# 0.0198f
C4 w_n211_n262# a_n73_n43# 0.0198f
C5 a_n33_n140# a_15_n43# 0.0193f
C6 a_15_n43# VSUBS 0.0453f
C7 a_n73_n43# VSUBS 0.0453f
C8 a_n33_n140# VSUBS 0.143f
C9 w_n211_n262# VSUBS 0.752f
.ends

.subckt sky130_fd_pr__nfet_01v8_L9ESAD a_n175_n190# a_n73_n50# a_n33_n138# a_15_n50#
X0 a_15_n50# a_n33_n138# a_n73_n50# a_n175_n190# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_n73_n50# a_15_n50# 0.0826f
C1 a_n73_n50# a_n33_n138# 0.0216f
C2 a_n33_n138# a_15_n50# 0.0216f
C3 a_15_n50# a_n175_n190# 0.0704f
C4 a_n73_n50# a_n175_n190# 0.0797f
C5 a_n33_n138# a_n175_n190# 0.315f
.ends

.subckt th11 V11 Vin Vn m1_577_n654# Vp m1_705_187#
XXM0 Vn Vp Vn m1_577_n654# Vn sky130_fd_pr__pfet_01v8_XGAKDL
XXM1 Vn Vin m1_577_n654# m1_705_187# sky130_fd_pr__nfet_01v8_4X3CDA
XXM2 m1_705_187# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_MWB9BZ
XXM3 V11 Vp m1_705_187# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM4 Vn Vn m1_705_187# V11 sky130_fd_pr__nfet_01v8_L9ESAD
C0 Vn V11 0.00327f
C1 m1_577_n654# V11 6.11e-19
C2 Vin V11 2.69e-19
C3 Vn m1_705_187# 0.463f
C4 m1_577_n654# m1_705_187# 0.0258f
C5 Vp Vn 0.0775f
C6 Vin m1_705_187# 0.0649f
C7 m1_577_n654# Vp 0.0405f
C8 Vin Vp 0.285f
C9 m1_705_187# V11 0.376f
C10 Vp V11 0.026f
C11 Vp m1_705_187# 0.286f
C12 m1_577_n654# Vn 0.0457f
C13 Vin Vn 0.135f
C14 Vin m1_577_n654# 0.213f
C15 Vp 0 2.61f
C16 m1_705_187# 0 0.602f
C17 V11 0 0.404f
C18 Vn 0 0.355f
C19 Vin 0 1.27f
C20 m1_577_n654# 0 0.286f
.ends

.subckt sky130_fd_pr__nfet_01v8_42G4RD a_n80_n42# a_n148_n216# a_n33_n130# a_22_n42#
X0 a_22_n42# a_n33_n130# a_n80_n42# a_n148_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_n33_n130# a_22_n42# 0.00866f
C1 a_n80_n42# a_22_n42# 0.0604f
C2 a_n33_n130# a_n80_n42# 0.00866f
C3 a_22_n42# a_n148_n216# 0.0698f
C4 a_n80_n42# a_n148_n216# 0.0698f
C5 a_n33_n130# a_n148_n216# 0.321f
.ends

.subckt sky130_fd_pr__pfet_01v8_DDPLQ8 a_n77_n42# w_n215_n261# a_n33_n139# a_19_n42#
+ VSUBS
X0 a_19_n42# a_n33_n139# a_n77_n42# w_n215_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 w_n215_n261# a_n77_n42# 0.017f
C1 a_n33_n139# a_n77_n42# 0.0127f
C2 a_19_n42# a_n77_n42# 0.0641f
C3 w_n215_n261# a_n33_n139# 0.181f
C4 w_n215_n261# a_19_n42# 0.0399f
C5 a_19_n42# a_n33_n139# 0.0127f
C6 a_19_n42# VSUBS 0.035f
C7 a_n77_n42# VSUBS 0.05f
C8 a_n33_n139# VSUBS 0.149f
C9 w_n215_n261# VSUBS 0.797f
.ends

.subckt sky130_fd_pr__nfet_01v8_VWP3K3 a_n33_n130# a_15_n42# a_n141_182# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n141_182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n33_n130# a_15_n42# 0.0209f
C1 a_n73_n42# a_15_n42# 0.0699f
C2 a_n33_n130# a_n73_n42# 0.0209f
C3 a_15_n42# a_n141_182# 0.0643f
C4 a_n73_n42# a_n141_182# 0.0643f
C5 a_n33_n130# a_n141_182# 0.317f
.ends

.subckt sky130_fd_pr__pfet_01v8_LZD9A4 a_n80_n42# a_22_n42# a_n33_n139# w_n218_n261#
+ VSUBS
X0 a_22_n42# a_n33_n139# a_n80_n42# w_n218_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 w_n218_n261# a_n80_n42# 0.0222f
C1 a_n33_n139# a_n80_n42# 0.0084f
C2 a_22_n42# a_n80_n42# 0.0604f
C3 w_n218_n261# a_n33_n139# 0.185f
C4 w_n218_n261# a_22_n42# 0.0222f
C5 a_22_n42# a_n33_n139# 0.0084f
C6 a_22_n42# VSUBS 0.0474f
C7 a_n80_n42# VSUBS 0.0474f
C8 a_n33_n139# VSUBS 0.149f
C9 w_n218_n261# VSUBS 0.775f
.ends

.subckt sky130_fd_pr__nfet_01v8_VRD6K3 a_n77_n42# a_n145_n214# a_n33_n130# a_19_n42#
X0 a_19_n42# a_n33_n130# a_n77_n42# a_n145_n214# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_n33_n130# a_19_n42# 0.0136f
C1 a_n77_n42# a_19_n42# 0.0641f
C2 a_n33_n130# a_n77_n42# 0.0136f
C3 a_19_n42# a_n145_n214# 0.0677f
C4 a_n77_n42# a_n145_n214# 0.0677f
C5 a_n33_n130# a_n145_n214# 0.32f
.ends

.subckt th04 Vp V04 Vin Vn m1_620_n488# m1_892_n998#
XXM0 m1_892_n998# Vn Vin Vn sky130_fd_pr__nfet_01v8_42G4RD
XXM1 m1_620_n488# Vp Vin m1_892_n998# Vn sky130_fd_pr__pfet_01v8_DDPLQ8
XXM2 Vp m1_620_n488# Vn Vp sky130_fd_pr__nfet_01v8_VWP3K3
XXM3 Vp V04 m1_892_n998# Vp Vn sky130_fd_pr__pfet_01v8_LZD9A4
XXM4 Vn Vn m1_892_n998# V04 sky130_fd_pr__nfet_01v8_VRD6K3
C0 m1_620_n488# m1_892_n998# 0.0117f
C1 m1_620_n488# V04 0.00264f
C2 m1_620_n488# Vin 0.0346f
C3 m1_892_n998# V04 0.13f
C4 m1_620_n488# Vp 0.17f
C5 m1_892_n998# Vin 0.463f
C6 V04 Vin 0.00141f
C7 m1_620_n488# Vn 2.16e-19
C8 m1_892_n998# Vp 0.383f
C9 V04 Vp 0.0462f
C10 Vn m1_892_n998# 0.1f
C11 Vp Vin 0.14f
C12 Vn V04 0.0639f
C13 Vn Vin 0.0468f
C14 Vn Vp 0.0386f
C15 Vin 0 0.679f
C16 V04 0 0.287f
C17 Vn 0 0.259f
C18 m1_892_n998# 0 0.832f
C19 Vp 0 2.13f
C20 m1_620_n488# 0 0.0632f
.ends

.subckt Analog Vin V01 V02 V03 V04 V08 V07 V06 V09 V10 V11 V12 V13 V14 V15 V05 th01_0/m1_991_n1219#
+ th10_0/m1_502_n495# th15_0/m1_597_n912# th13_0/m1_831_275# th15_0/m1_849_n157# th15_0/Vin
+ th07_0/m1_808_n892# th02_0/m1_571_144# th14_0/m1_891_419# th12_0/m1_529_n42# th09_0/m1_962_372#
+ th13_0/m1_559_n458# th02_0/m1_983_133# th04_0/m1_892_n998# th11_0/m1_577_n654# th04_0/m1_620_n488#
+ th12_0/m1_394_n856# th05_0/m1_752_n794# th09_0/m1_485_n505# th03_0/m1_890_n844#
+ th03_0/m1_638_n591# th06_0/m1_904_n796# th14_0/m1_641_n318# th10_0/m1_536_174# th11_0/m1_705_187#
+ th08_0/m1_477_n803# Vp th01_0/m1_571_n501# Vn
Xth02_0 th15_0/Vin V02 Vp th02_0/m1_983_133# th02_0/m1_571_144# Vn th02
Xth09_0 V09 Vin Vn th09_0/m1_485_n505# Vp th09_0/m1_962_372# th09
Xth14_0 V14 th15_0/Vin Vn th14_0/m1_641_n318# Vp th14_0/m1_891_419# th14
Xth07_0 Vin V07 Vp th07_0/m1_808_n892# Vn th07
Xth12_0 Vp V12 Vin th12_0/m1_529_n42# th12_0/m1_394_n856# Vn th12
Xth05_0 Vp V05 Vin th05_0/m1_752_n794# Vn th05
Xth10_0 Vp V10 Vin Vn th10_0/m1_502_n495# th10_0/m1_536_174# th10
Xth03_0 V03 Vin Vp th03_0/m1_890_n844# th03_0/m1_638_n591# Vn th03
Xth01_0 Vp th15_0/Vin V01 th01_0/m1_991_n1219# Vn th01_0/m1_571_n501# th01
Xpreamp_0 Vp Vin th15_0/Vin Vn preamp
Xth15_0 V15 th15_0/Vin th15_0/m1_597_n912# Vp th15_0/m1_849_n157# Vn th15
Xth08_0 Vin V08 th08_0/m1_477_n803# Vp Vn th08
Xth13_0 V13 Vin th13_0/m1_831_275# Vn Vp th13_0/m1_559_n458# th13
Xth06_0 Vp Vin V06 Vn th06_0/m1_904_n796# th06
Xth11_0 V11 Vin Vn th11_0/m1_577_n654# Vp th11_0/m1_705_187# th11
Xth04_0 Vp V04 Vin Vn th04_0/m1_620_n488# th04_0/m1_892_n998# th04
C0 th10_0/m1_536_174# th12_0/m1_529_n42# 0.002f
C1 th09_0/m1_962_372# V09 8.77e-19
C2 Vp th02_0/m1_983_133# 0.0442f
C3 th01_0/m1_991_n1219# Vn 0.00203f
C4 Vp th06_0/m1_904_n796# 0.0232f
C5 th14_0/m1_641_n318# th09_0/m1_485_n505# 6.8e-20
C6 th15_0/m1_849_n157# V15 0.0154f
C7 th12_0/m1_529_n42# V14 1.86e-19
C8 th06_0/m1_904_n796# th08_0/m1_477_n803# 2.84e-21
C9 V06 th07_0/m1_808_n892# 5.69e-20
C10 th09_0/m1_962_372# th02_0/m1_571_144# 0.0112f
C11 V13 th15_0/m1_849_n157# 0.0171f
C12 Vin th10_0/m1_502_n495# 1.09e-19
C13 V06 Vn 5.44e-19
C14 Vp th11_0/m1_577_n654# 0.0262f
C15 th03_0/m1_638_n591# Vn 0.0534f
C16 Vn V02 0.00543f
C17 Vp th12_0/m1_529_n42# 0.0641f
C18 Vp V11 0.0406f
C19 V07 Vin 0.0909f
C20 th12_0/m1_529_n42# th14_0/m1_891_419# 0.0381f
C21 th15_0/Vin Vn 1.48f
C22 V11 th14_0/m1_891_419# 0.0143f
C23 th03_0/m1_890_n844# th02_0/m1_983_133# 0.00411f
C24 th12_0/m1_529_n42# th12_0/m1_394_n856# 1.78e-33
C25 th13_0/m1_831_275# th09_0/m1_485_n505# 2.23e-19
C26 V09 th14_0/m1_641_n318# 6.83e-21
C27 V13 th13_0/m1_831_275# 0.0112f
C28 V05 th05_0/m1_752_n794# 1.39e-19
C29 th15_0/Vin th01_0/m1_991_n1219# 0.00291f
C30 th01_0/m1_991_n1219# th04_0/m1_620_n488# 7.52e-20
C31 Vp th10_0/m1_502_n495# 0.035f
C32 V07 V08 6.64e-21
C33 V03 th02_0/m1_983_133# 2.47e-20
C34 Vn V15 2.4e-20
C35 Vp V07 0.0372f
C36 th15_0/Vin th03_0/m1_638_n591# 0.0177f
C37 th15_0/Vin V02 0.00312f
C38 th08_0/m1_477_n803# V07 9.47e-21
C39 Vn th09_0/m1_485_n505# 0.0537f
C40 th13_0/m1_559_n458# Vn 0.017f
C41 V04 Vin 0.175f
C42 th15_0/Vin th04_0/m1_620_n488# 2.61e-19
C43 th06_0/m1_904_n796# V05 1.38e-20
C44 V13 Vn 0.0182f
C45 th02_0/m1_571_144# th11_0/m1_705_187# 1.03e-19
C46 th10_0/m1_536_174# Vin 0.0133f
C47 Vn V10 0.0168f
C48 V04 th04_0/m1_892_n998# 1.47e-19
C49 V04 V08 2.69e-20
C50 th07_0/m1_808_n892# th05_0/m1_752_n794# 1.42e-20
C51 Vn V09 0.0232f
C52 V14 Vin 0.00129f
C53 th15_0/Vin V15 1.81e-19
C54 Vp V04 0.00153f
C55 Vn th05_0/m1_752_n794# 0.00258f
C56 th04_0/m1_892_n998# Vin 0.111f
C57 th15_0/Vin th09_0/m1_485_n505# 0.113f
C58 th13_0/m1_559_n458# th15_0/Vin 0.11f
C59 Vin V08 0.164f
C60 V04 th08_0/m1_477_n803# 4.48e-19
C61 Vn th02_0/m1_571_144# 0.0142f
C62 th15_0/Vin V13 1e-23
C63 Vp Vin 1.96f
C64 V11 th11_0/m1_705_187# 5.77e-19
C65 th08_0/m1_477_n803# Vin 0.055f
C66 th14_0/m1_891_419# Vin 0.0347f
C67 Vn V12 0.0372f
C68 th12_0/m1_529_n42# th13_0/m1_831_275# 1.36e-20
C69 th12_0/m1_394_n856# Vin 0.0013f
C70 Vp th10_0/m1_536_174# 0.0514f
C71 th06_0/m1_904_n796# th07_0/m1_808_n892# 2e-19
C72 th04_0/m1_892_n998# V08 3.48e-19
C73 V06 th05_0/m1_752_n794# 0.001f
C74 Vn th02_0/m1_983_133# 0.157f
C75 th06_0/m1_904_n796# Vn 0.00332f
C76 Vp V14 0.0751f
C77 th15_0/Vin V09 0.0644f
C78 Vp th04_0/m1_892_n998# 0.0374f
C79 V14 th14_0/m1_891_419# 0.0202f
C80 th03_0/m1_890_n844# Vin 4.79e-20
C81 Vp V08 0.0346f
C82 th01_0/m1_571_n501# Vin 6.06e-19
C83 th13_0/m1_559_n458# th09_0/m1_485_n505# 0.00612f
C84 V13 V15 0.00246f
C85 th08_0/m1_477_n803# th04_0/m1_892_n998# 0.00506f
C86 th08_0/m1_477_n803# V08 0.00927f
C87 th15_0/Vin th02_0/m1_571_144# 0.00185f
C88 th09_0/m1_962_372# Vin 6.36e-19
C89 Vn th11_0/m1_577_n654# 0.0365f
C90 Vn th12_0/m1_529_n42# 0.0621f
C91 V11 Vn 0.0184f
C92 V04 V01 1.84e-20
C93 Vp th08_0/m1_477_n803# 0.0268f
C94 Vp th14_0/m1_891_419# 0.0102f
C95 Vp th12_0/m1_394_n856# 0.0145f
C96 th15_0/Vin V12 1.05e-21
C97 th06_0/m1_904_n796# V06 -1.42e-32
C98 th12_0/m1_394_n856# th14_0/m1_891_419# 5.71e-20
C99 th02_0/m1_983_133# V02 0.0161f
C100 th03_0/m1_638_n591# th02_0/m1_983_133# 0.0193f
C101 V01 Vin 0.00532f
C102 th15_0/m1_597_n912# Vin 3.87e-19
C103 V03 Vin 4.84e-19
C104 th15_0/Vin th02_0/m1_983_133# 0.0246f
C105 V09 th09_0/m1_485_n505# 0.0182f
C106 th13_0/m1_559_n458# V09 0.00378f
C107 Vp th03_0/m1_890_n844# 0.0291f
C108 Vp th01_0/m1_571_n501# 0.0265f
C109 Vn th10_0/m1_502_n495# 0.00962f
C110 V05 Vin 0.00116f
C111 V07 th07_0/m1_808_n892# 0.00298f
C112 th14_0/m1_641_n318# Vin 0.0621f
C113 th11_0/m1_577_n654# V02 3.56e-21
C114 Vp th09_0/m1_962_372# 0.0369f
C115 th02_0/m1_571_144# th09_0/m1_485_n505# 0.00503f
C116 th15_0/m1_849_n157# Vin 0.00238f
C117 th15_0/Vin th11_0/m1_577_n654# 0.016f
C118 Vn V07 0.00179f
C119 th04_0/m1_892_n998# V01 0.0123f
C120 th15_0/Vin th12_0/m1_529_n42# 0.0262f
C121 V11 th15_0/Vin 0.00172f
C122 Vp V01 0.116f
C123 th03_0/m1_890_n844# th01_0/m1_571_n501# 0.00797f
C124 Vp th15_0/m1_597_n912# -2.84e-32
C125 Vp V03 0.011f
C126 th11_0/m1_705_187# Vin 0.278f
C127 th08_0/m1_477_n803# V01 4.9e-21
C128 th02_0/m1_983_133# th09_0/m1_485_n505# 0.00736f
C129 Vin th13_0/m1_831_275# 0.0149f
C130 Vp V05 0.00375f
C131 V09 th02_0/m1_571_144# 3.21e-19
C132 V06 V07 5.71e-22
C133 Vp th14_0/m1_641_n318# 0.0569f
C134 V04 th07_0/m1_808_n892# 6.58e-21
C135 Vp th15_0/m1_849_n157# 0.0962f
C136 th14_0/m1_641_n318# th12_0/m1_394_n856# 0.00861f
C137 th13_0/m1_559_n458# th12_0/m1_529_n42# 9.14e-21
C138 th03_0/m1_890_n844# V03 7.56e-19
C139 V04 Vn 0.00815f
C140 th07_0/m1_808_n892# Vin 0.0324f
C141 Vp th11_0/m1_705_187# 0.0213f
C142 Vn Vin 1.97f
C143 V04 th01_0/m1_991_n1219# 2.28e-19
C144 th06_0/m1_904_n796# th05_0/m1_752_n794# 0.00251f
C145 th11_0/m1_705_187# th14_0/m1_891_419# 0.00195f
C146 Vp th13_0/m1_831_275# 0.0414f
C147 th11_0/m1_705_187# th12_0/m1_394_n856# 6.45e-22
C148 V10 th12_0/m1_529_n42# 2.39e-20
C149 th10_0/m1_536_174# Vn 0.0537f
C150 th12_0/m1_394_n856# th13_0/m1_831_275# 4.06e-20
C151 th01_0/m1_991_n1219# Vin 0.0315f
C152 th04_0/m1_892_n998# th07_0/m1_808_n892# 1.1e-19
C153 th07_0/m1_808_n892# V08 0.0102f
C154 Vn V14 0.0201f
C155 Vn th04_0/m1_892_n998# 4.09e-20
C156 th01_0/m1_571_n501# th11_0/m1_705_187# 9.49e-20
C157 Vn V08 7.17e-19
C158 th11_0/m1_577_n654# th02_0/m1_571_144# 0.0183f
C159 Vp th07_0/m1_808_n892# 0.0183f
C160 V06 Vin 0.094f
C161 V11 th02_0/m1_571_144# 4.75e-20
C162 th08_0/m1_477_n803# th07_0/m1_808_n892# 4.41e-19
C163 Vin V02 0.292f
C164 Vp Vn 1.69f
C165 th12_0/m1_529_n42# V12 3.26e-19
C166 th15_0/Vin Vin 0.87f
C167 th01_0/m1_991_n1219# th04_0/m1_892_n998# 0.0226f
C168 th04_0/m1_620_n488# Vin 0.00123f
C169 Vn th08_0/m1_477_n803# 0.00115f
C170 Vn th14_0/m1_891_419# 0.0525f
C171 Vn th12_0/m1_394_n856# 0.0035f
C172 th15_0/Vin th10_0/m1_536_174# 3.79e-20
C173 th11_0/m1_577_n654# th02_0/m1_983_133# 1.64e-19
C174 Vp th01_0/m1_991_n1219# 0.0315f
C175 th01_0/m1_991_n1219# th14_0/m1_891_419# 0.0018f
C176 th15_0/Vin V14 6.88e-20
C177 V07 th05_0/m1_752_n794# 4.77e-21
C178 th03_0/m1_890_n844# Vn 0.0101f
C179 th01_0/m1_571_n501# Vn 0.00241f
C180 th15_0/Vin th04_0/m1_892_n998# 0.00125f
C181 Vp V06 0.025f
C182 th04_0/m1_620_n488# V08 3.51e-21
C183 th14_0/m1_641_n318# th11_0/m1_705_187# 5.69e-22
C184 Vp th03_0/m1_638_n591# 0.0167f
C185 Vp V02 0.00255f
C186 th09_0/m1_962_372# Vn 0.00557f
C187 V11 th11_0/m1_577_n654# 1.77e-19
C188 Vp th15_0/Vin 1.24f
C189 Vp th04_0/m1_620_n488# 0.00246f
C190 Vin th09_0/m1_485_n505# 0.0287f
C191 th15_0/m1_849_n157# th13_0/m1_831_275# 0.0859f
C192 th13_0/m1_559_n458# Vin 0.0257f
C193 th15_0/Vin th14_0/m1_891_419# 0.00394f
C194 th04_0/m1_620_n488# th08_0/m1_477_n803# 6.18e-20
C195 th15_0/Vin th12_0/m1_394_n856# 0.0129f
C196 V13 Vin 0.00669f
C197 Vn V01 0.00263f
C198 Vn th15_0/m1_597_n912# 0.106f
C199 Vn V03 2.75e-19
C200 th06_0/m1_904_n796# V07 0.00384f
C201 th03_0/m1_890_n844# V02 0.00134f
C202 V10 Vin 0.00422f
C203 th12_0/m1_529_n42# th10_0/m1_502_n495# 8.5e-20
C204 th03_0/m1_890_n844# th15_0/Vin 0.00307f
C205 th15_0/Vin th01_0/m1_571_n501# -5.68e-32
C206 Vn V05 6.36e-19
C207 th01_0/m1_991_n1219# V01 0.00159f
C208 Vn th14_0/m1_641_n318# 0.0401f
C209 Vp V15 0.00307f
C210 V09 Vin 0.00465f
C211 th15_0/Vin th09_0/m1_962_372# 0.0637f
C212 Vn th15_0/m1_849_n157# 0.0342f
C213 th10_0/m1_536_174# V10 0.0035f
C214 Vp th09_0/m1_485_n505# 0.0355f
C215 Vp th13_0/m1_559_n458# 0.0105f
C216 th05_0/m1_752_n794# Vin 0.00963f
C217 th14_0/m1_891_419# th09_0/m1_485_n505# 3.27e-19
C218 Vp V13 0.00713f
C219 th02_0/m1_571_144# Vin 0.00869f
C220 th13_0/m1_559_n458# th12_0/m1_394_n856# 3.47e-20
C221 th15_0/Vin V01 3.18e-19
C222 th04_0/m1_620_n488# V01 0.00118f
C223 Vn th11_0/m1_705_187# -0.0527f
C224 th15_0/Vin V03 1.39e-20
C225 th15_0/Vin th15_0/m1_597_n912# 0.0049f
C226 Vin V12 1.77e-19
C227 Vn th13_0/m1_831_275# 0.0355f
C228 Vp V10 0.0332f
C229 th10_0/m1_536_174# V12 9.23e-19
C230 th01_0/m1_991_n1219# th11_0/m1_705_187# 0.00184f
C231 th02_0/m1_983_133# Vin 0.0835f
C232 th15_0/Vin th14_0/m1_641_n318# 0.0354f
C233 Vp V09 0.00542f
C234 th06_0/m1_904_n796# Vin 0.0348f
C235 V09 th14_0/m1_891_419# 3.7e-19
C236 th15_0/Vin th15_0/m1_849_n157# 6.18e-19
C237 Vp th05_0/m1_752_n794# 8.03e-19
C238 Vp th02_0/m1_571_144# 0.026f
C239 Vn th07_0/m1_808_n892# 0.00532f
C240 th11_0/m1_577_n654# Vin 0.0113f
C241 th12_0/m1_529_n42# Vin 0.0104f
C242 V11 Vin 0.0579f
C243 Vp V12 0.0535f
C244 th15_0/Vin th11_0/m1_705_187# 0.0359f
C245 th14_0/m1_891_419# V12 2.97e-19
C246 th06_0/m1_904_n796# V08 9.74e-22
C247 th15_0/Vin th13_0/m1_831_275# 0.0168f
C248 th12_0/m1_394_n856# V12 2.12e-19
C249 V04 0 0.191f
C250 th04_0/m1_892_n998# 0 0.832f
C251 th04_0/m1_620_n488# 0 0.0632f
C252 th11_0/m1_705_187# 0 0.602f
C253 V11 0 0.349f
C254 Vin 0 15f
C255 th11_0/m1_577_n654# 0 0.286f
C256 V06 0 0.132f
C257 th06_0/m1_904_n796# 0 0.495f
C258 th13_0/m1_831_275# 0 1.05f
C259 V13 0 0.371f
C260 th13_0/m1_559_n458# 0 0.286f
C261 th08_0/m1_477_n803# 0 0.577f
C262 V08 0 0.139f
C263 V15 0 0.356f
C264 th15_0/m1_849_n157# 0 1.28f
C265 th15_0/m1_597_n912# 0 0.19f
C266 Vn 0 6.57f
C267 th01_0/m1_991_n1219# 0 1.24f
C268 V01 0 0.241f
C269 th01_0/m1_571_n501# 0 0.194f
C270 th15_0/Vin 0 5.76f
C271 Vp 0 43.6f
C272 V03 0 0.303f
C273 th03_0/m1_890_n844# 0 1.05f
C274 th03_0/m1_638_n591# 0 0.224f
C275 th10_0/m1_536_174# 0 0.825f
C276 V10 0 0.269f
C277 th10_0/m1_502_n495# 0 0.146f
C278 th05_0/m1_752_n794# 0 0.788f
C279 V05 0 0.321f
C280 th12_0/m1_529_n42# 0 0.861f
C281 V12 0 0.468f
C282 th12_0/m1_394_n856# 0 0.215f
C283 th07_0/m1_808_n892# 0 0.511f
C284 V07 0 0.159f
C285 th14_0/m1_891_419# 0 1.48f
C286 V14 0 0.233f
C287 th14_0/m1_641_n318# 0 0.241f
C288 th09_0/m1_485_n505# 0 1.18f
C289 V09 0 0.213f
C290 th09_0/m1_962_372# 0 0.118f
C291 V02 0 0.211f
C292 th02_0/m1_983_133# 0 1.44f
C293 th02_0/m1_571_144# 0 0.252f
.ends

.subckt analog_therm Vp Vin Vn
Xtherm_raw_0 therm_raw_0/b[0] therm_raw_0/b[2] therm_raw_0/b[3] Analog_0/V12 Analog_0/V13
+ Analog_0/V14 Analog_0/V15 Analog_0/V02 Analog_0/V03 Analog_0/V05 Analog_0/V06 Analog_0/V09
+ Analog_0/V10 therm_raw_0/input3/a_27_47# therm_raw_0/net7 therm_raw_0/input13/a_27_47#
+ therm_raw_0/net3 therm_raw_0/net15 therm_raw_0/net14 therm_raw_0/input7/a_27_47#
+ therm_raw_0/_04_ therm_raw_0/input9/a_75_212# therm_raw_0/b[1] therm_raw_0/_27_/a_27_297#
+ therm_raw_0/input1/a_75_212# therm_raw_0/input5/a_62_47# therm_raw_0/net2 Analog_0/V01
+ therm_raw_0/input5/a_381_47# therm_raw_0/_19_ therm_raw_0/net8 therm_raw_0/input8/a_27_47#
+ Analog_0/V08 therm_raw_0/output17/a_27_47# therm_raw_0/_01_ therm_raw_0/_02_ therm_raw_0/input15/a_27_47#
+ therm_raw_0/input5/a_558_47# therm_raw_0/_15_ Analog_0/V04 therm_raw_0/input5/a_664_47#
+ therm_raw_0/_08_ therm_raw_0/input6/a_27_47# therm_raw_0/net17 therm_raw_0/net5
+ Vp Analog_0/V11 Vn Analog_0/V07 therm_raw
XAnalog_0 Vin Analog_0/V01 Analog_0/V02 Analog_0/V03 Analog_0/V04 Analog_0/V08 Analog_0/V07
+ Analog_0/V06 Analog_0/V09 Analog_0/V10 Analog_0/V11 Analog_0/V12 Analog_0/V13 Analog_0/V14
+ Analog_0/V15 Analog_0/V05 Analog_0/th01_0/m1_991_n1219# Analog_0/th10_0/m1_502_n495#
+ Analog_0/th15_0/m1_597_n912# Analog_0/th13_0/m1_831_275# Analog_0/th15_0/m1_849_n157#
+ Analog_0/th15_0/Vin Analog_0/th07_0/m1_808_n892# Analog_0/th02_0/m1_571_144# Analog_0/th14_0/m1_891_419#
+ Analog_0/th12_0/m1_529_n42# Analog_0/th09_0/m1_962_372# Analog_0/th13_0/m1_559_n458#
+ Analog_0/th02_0/m1_983_133# Analog_0/th04_0/m1_892_n998# Analog_0/th11_0/m1_577_n654#
+ Analog_0/th04_0/m1_620_n488# Analog_0/th12_0/m1_394_n856# Analog_0/th05_0/m1_752_n794#
+ Analog_0/th09_0/m1_485_n505# Analog_0/th03_0/m1_890_n844# Analog_0/th03_0/m1_638_n591#
+ Analog_0/th06_0/m1_904_n796# Analog_0/th14_0/m1_641_n318# Analog_0/th10_0/m1_536_174#
+ Analog_0/th11_0/m1_705_187# Analog_0/th08_0/m1_477_n803# Vp Analog_0/th01_0/m1_571_n501#
+ Vn Analog
C0 Analog_0/th04_0/m1_620_n488# Analog_0/V03 1.36e-19
C1 Analog_0/th04_0/m1_892_n998# Analog_0/th01_0/m1_991_n1219# -0.0169f
C2 Analog_0/th15_0/Vin Analog_0/V03 0.132f
C3 Analog_0/th14_0/m1_891_419# Analog_0/V01 1.15e-19
C4 Analog_0/V02 Vp 0.374f
C5 Analog_0/th15_0/Vin Analog_0/V01 0.00129f
C6 Analog_0/V07 therm_raw_0/input8/a_27_47# 5.01e-21
C7 Analog_0/V12 Analog_0/th12_0/m1_529_n42# 0.00558f
C8 Analog_0/V09 Analog_0/th02_0/m1_571_144# 0.00844f
C9 Analog_0/V11 Analog_0/th12_0/m1_529_n42# 0.00638f
C10 therm_raw_0/input1/a_75_212# Analog_0/V11 1.77e-19
C11 Analog_0/th11_0/m1_577_n654# Analog_0/V01 5.35e-20
C12 Vin Analog_0/th05_0/m1_752_n794# -1.94e-20
C13 Analog_0/th02_0/m1_571_144# Vin -5.88e-21
C14 Analog_0/th01_0/m1_991_n1219# Analog_0/V03 0.0286f
C15 Analog_0/V08 Analog_0/V02 0.148f
C16 therm_raw_0/net2 Analog_0/V11 -8.67e-21
C17 Analog_0/th01_0/m1_991_n1219# Analog_0/V01 0.0525f
C18 Analog_0/th14_0/m1_891_419# Vp -9.9e-20
C19 Analog_0/th15_0/Vin Vp -2.28e-19
C20 Analog_0/th06_0/m1_904_n796# Analog_0/V02 0.00793f
C21 Analog_0/V07 Analog_0/th08_0/m1_477_n803# 4.51e-21
C22 Analog_0/V09 Vin 0.17f
C23 Analog_0/V15 Analog_0/th15_0/Vin 0.0318f
C24 Analog_0/V10 Analog_0/th10_0/m1_536_174# 0.0602f
C25 Analog_0/V07 Analog_0/V06 0.0777f
C26 Analog_0/th07_0/m1_808_n892# Analog_0/V02 0.0224f
C27 Analog_0/th01_0/m1_991_n1219# Vp -0.00523f
C28 Vin Analog_0/V12 4.62e-19
C29 therm_raw_0/input5/a_62_47# Analog_0/V14 0.00136f
C30 Vin Analog_0/V11 0.159f
C31 Analog_0/V10 Analog_0/V14 0.00199f
C32 Analog_0/V04 Vin 0.0574f
C33 Analog_0/V12 Analog_0/V11 0.121f
C34 therm_raw_0/_15_ therm_raw_0/input3/a_27_47# 2.22e-34
C35 Analog_0/V14 Analog_0/V01 0.0181f
C36 therm_raw_0/_15_ Vp -4.97e-32
C37 therm_raw_0/b[3] Analog_0/V12 0.0305f
C38 Analog_0/th10_0/m1_536_174# Vp -1.52e-21
C39 Analog_0/V05 Vp 0.00767f
C40 Analog_0/V09 Analog_0/th13_0/m1_559_n458# 3.18e-19
C41 therm_raw_0/output17/a_27_47# Analog_0/V11 5.42e-20
C42 Vin Analog_0/th11_0/m1_705_187# -1.09e-19
C43 Analog_0/V14 Vp 0.315f
C44 Analog_0/V07 Analog_0/V02 0.365f
C45 Analog_0/V10 therm_raw_0/input15/a_27_47# -5.55e-35
C46 Analog_0/th08_0/m1_477_n803# Analog_0/V02 0.0044f
C47 therm_raw_0/b[1] Analog_0/V01 0.00918f
C48 Analog_0/th11_0/m1_705_187# Analog_0/V11 0.00493f
C49 Analog_0/th06_0/m1_904_n796# Analog_0/V05 1.32e-20
C50 Analog_0/th01_0/m1_571_n501# Analog_0/V02 8.31e-19
C51 Analog_0/th15_0/Vin Analog_0/th09_0/m1_485_n505# -4.22e-20
C52 Analog_0/V06 Analog_0/V02 0.0412f
C53 Analog_0/V15 Analog_0/th15_0/m1_849_n157# 0.0256f
C54 Analog_0/th15_0/m1_597_n912# Analog_0/V15 0.00155f
C55 Analog_0/V13 Analog_0/th15_0/Vin 0.0338f
C56 Analog_0/th03_0/m1_638_n591# Analog_0/V02 6.44e-19
C57 therm_raw_0/net3 Vp 7.13e-20
C58 therm_raw_0/_04_ Analog_0/V14 2.04e-19
C59 Analog_0/V14 Analog_0/th10_0/m1_502_n495# 1.06e-19
C60 Vp therm_raw_0/b[1] 4.71e-19
C61 therm_raw_0/input1/a_75_212# Analog_0/V01 7.39e-20
C62 Analog_0/V09 Analog_0/th02_0/m1_983_133# 0.00361f
C63 Analog_0/th04_0/m1_892_n998# Vin -1.97e-19
C64 Vin Analog_0/th02_0/m1_983_133# -5.51e-19
C65 Analog_0/V09 Analog_0/V10 7.52e-19
C66 Vp Analog_0/th12_0/m1_529_n42# 1.14e-31
C67 therm_raw_0/input6/a_27_47# Analog_0/V10 1.11e-34
C68 Analog_0/V04 Analog_0/th04_0/m1_892_n998# 0.00165f
C69 Analog_0/th02_0/m1_571_144# Analog_0/th09_0/m1_962_372# 4.44e-34
C70 Analog_0/V10 Vin 1.81e-19
C71 Analog_0/V07 Analog_0/V05 2.33e-20
C72 Analog_0/V14 Analog_0/th14_0/m1_641_n318# 5.9e-20
C73 therm_raw_0/net2 Vp 0.00947f
C74 therm_raw_0/input5/a_62_47# Analog_0/V12 2.93e-19
C75 Vin Analog_0/V03 0.209f
C76 Analog_0/V10 Analog_0/V12 0.0944f
C77 Vin Analog_0/V01 0.0602f
C78 Analog_0/th02_0/m1_571_144# Vp 1.42e-32
C79 Analog_0/V09 Analog_0/th09_0/m1_962_372# 3.51e-19
C80 Analog_0/th04_0/m1_620_n488# Analog_0/V02 7.54e-20
C81 Analog_0/V06 Analog_0/V05 0.0587f
C82 Analog_0/V10 therm_raw_0/b[3] 0.00686f
C83 Analog_0/V13 Analog_0/th15_0/m1_849_n157# 0.0154f
C84 Analog_0/V13 Analog_0/th15_0/m1_597_n912# 1.93e-19
C85 Analog_0/V03 Analog_0/V11 1.2e-20
C86 Analog_0/th15_0/Vin Analog_0/V02 0.0561f
C87 Analog_0/V11 Analog_0/V01 0.0855f
C88 Analog_0/V04 Analog_0/V03 0.703f
C89 Analog_0/V14 therm_raw_0/_19_ 1.88e-19
C90 Analog_0/V04 Analog_0/V01 0.0664f
C91 Analog_0/V09 Vp 0.169f
C92 therm_raw_0/net2 therm_raw_0/_04_ -4.44e-34
C93 Analog_0/V14 therm_raw_0/input5/a_381_47# 1.06e-19
C94 Analog_0/V09 Analog_0/V15 0.743f
C95 Vin Vp 0.0115f
C96 therm_raw_0/input3/a_27_47# Analog_0/V12 1.58e-19
C97 Analog_0/V15 Vin 4.43e-19
C98 Analog_0/th01_0/m1_991_n1219# Analog_0/V02 0.00345f
C99 Analog_0/V12 Vp 0.284f
C100 Analog_0/V11 Vp 0.58f
C101 Analog_0/V04 Vp 0.0117f
C102 therm_raw_0/_27_/a_27_297# Vp 1.85e-19
C103 therm_raw_0/b[3] Vp 1.12e-19
C104 Analog_0/V08 Vin 0.181f
C105 Analog_0/V07 therm_raw_0/net7 4.14e-20
C106 Analog_0/th11_0/m1_705_187# Analog_0/V03 2.36e-19
C107 Analog_0/th11_0/m1_705_187# Analog_0/V01 0.00398f
C108 Analog_0/V14 therm_raw_0/net5 6.93e-19
C109 Analog_0/th12_0/m1_394_n856# Analog_0/V14 0.0145f
C110 Analog_0/th06_0/m1_904_n796# Vin -0.00189f
C111 therm_raw_0/net8 Vp 3.95e-20
C112 Analog_0/V09 Analog_0/th13_0/m1_831_275# 0.0253f
C113 Analog_0/V08 Analog_0/V04 0.426f
C114 therm_raw_0/_04_ Analog_0/V12 6.13e-20
C115 Analog_0/th07_0/m1_808_n892# Vin -8.48e-19
C116 Vin Analog_0/th10_0/m1_502_n495# 0.025f
C117 therm_raw_0/_04_ Analog_0/V11 -1.56e-20
C118 Analog_0/th06_0/m1_904_n796# Analog_0/V04 0.0012f
C119 Analog_0/th03_0/m1_890_n844# Analog_0/V03 0.0091f
C120 therm_raw_0/net17 Vp -1.42e-32
C121 Analog_0/th07_0/m1_808_n892# Analog_0/V04 5.62e-20
C122 therm_raw_0/net15 Vp 0.00128f
C123 Analog_0/th02_0/m1_571_144# Analog_0/th09_0/m1_485_n505# -1.12e-19
C124 Analog_0/V07 Analog_0/th05_0/m1_752_n794# 7.58e-20
C125 Analog_0/th12_0/m1_394_n856# therm_raw_0/b[1] 5.17e-20
C126 therm_raw_0/net2 therm_raw_0/_19_ -8.88e-34
C127 Analog_0/V09 Analog_0/th09_0/m1_485_n505# 0.152f
C128 Analog_0/V09 Analog_0/th14_0/m1_641_n318# 9.22e-20
C129 Analog_0/V13 Analog_0/V09 0.487f
C130 Analog_0/V14 Analog_0/th14_0/m1_891_419# 0.0676f
C131 Analog_0/V14 Analog_0/th15_0/Vin 0.0061f
C132 Analog_0/th04_0/m1_892_n998# Analog_0/V03 0.0726f
C133 Vin Analog_0/th09_0/m1_485_n505# -5.64e-19
C134 Analog_0/V06 Analog_0/th05_0/m1_752_n794# 0.0128f
C135 Analog_0/th04_0/m1_892_n998# Analog_0/V01 -0.00984f
C136 Analog_0/V13 Vin 0.0124f
C137 Analog_0/V07 Vin 0.0546f
C138 Analog_0/th14_0/m1_641_n318# Analog_0/V11 0.00195f
C139 Vin Analog_0/th08_0/m1_477_n803# -1.26e-19
C140 therm_raw_0/net2 therm_raw_0/net5 7.11e-33
C141 Analog_0/V06 Vin 0.188f
C142 Analog_0/th04_0/m1_892_n998# Vp 0.00896f
C143 Analog_0/V03 Analog_0/V01 0.66f
C144 Analog_0/V07 Analog_0/V04 0.0925f
C145 therm_raw_0/_19_ Analog_0/V12 6.25e-21
C146 therm_raw_0/input5/a_558_47# Vp -2.84e-32
C147 Analog_0/V04 Analog_0/th08_0/m1_477_n803# 4.31e-20
C148 Analog_0/V14 Analog_0/th10_0/m1_536_174# 0.00621f
C149 therm_raw_0/input5/a_664_47# Vp -2.84e-32
C150 Analog_0/V04 Analog_0/V06 0.0364f
C151 Analog_0/V10 Vp 0.00425f
C152 Analog_0/V08 Analog_0/th04_0/m1_892_n998# 3.24e-19
C153 Analog_0/V10 Analog_0/V15 0.0185f
C154 Analog_0/V03 Vp 0.563f
C155 Analog_0/V02 Analog_0/th05_0/m1_752_n794# 1.1e-19
C156 Vp Analog_0/V01 0.0753f
C157 Analog_0/th12_0/m1_394_n856# Analog_0/V11 5.23e-22
C158 Analog_0/V09 Analog_0/V02 5.38e-19
C159 Analog_0/V08 Analog_0/V03 0.0991f
C160 Analog_0/V08 Analog_0/V01 0.21f
C161 Analog_0/th06_0/m1_904_n796# Analog_0/V03 2.01e-19
C162 Vin Analog_0/V02 0.399f
C163 therm_raw_0/_02_ Vp 3.51e-20
C164 Analog_0/th07_0/m1_808_n892# Analog_0/V03 0.00405f
C165 Analog_0/V15 Vp 0.0118f
C166 Analog_0/V14 therm_raw_0/b[1] 0.0162f
C167 Analog_0/V04 Analog_0/V02 0.0476f
C168 Analog_0/V09 Analog_0/th15_0/Vin 0.0131f
C169 Analog_0/V08 Vp 0.00655f
C170 Analog_0/V07 therm_raw_0/input9/a_75_212# 5.01e-21
C171 Vin Analog_0/th14_0/m1_891_419# -0.015f
C172 Analog_0/th09_0/m1_485_n505# Analog_0/th02_0/m1_983_133# -1.49e-20
C173 therm_raw_0/_04_ Vp 7.33e-19
C174 Vin Analog_0/th15_0/Vin -3.32e-19
C175 Analog_0/th10_0/m1_502_n495# Vp -0.012f
C176 Analog_0/th14_0/m1_891_419# Analog_0/V11 0.068f
C177 Analog_0/th15_0/Vin Analog_0/V11 0.0102f
C178 Vp Analog_0/th13_0/m1_831_275# -1.78e-19
C179 therm_raw_0/input1/a_75_212# Analog_0/V14 6.76e-20
C180 Analog_0/V14 Analog_0/th12_0/m1_529_n42# 0.0164f
C181 Vin Analog_0/th01_0/m1_991_n1219# -0.0112f
C182 Analog_0/th06_0/m1_904_n796# Analog_0/V08 0.00229f
C183 Analog_0/V05 Analog_0/th05_0/m1_752_n794# 8.69e-19
C184 Analog_0/V11 Analog_0/th11_0/m1_577_n654# 1.23e-19
C185 Analog_0/V07 therm_raw_0/input7/a_27_47# 4.62e-20
C186 Analog_0/V08 Analog_0/th07_0/m1_808_n892# 0.00506f
C187 therm_raw_0/net2 Analog_0/V14 0.00832f
C188 Analog_0/th01_0/m1_991_n1219# Analog_0/V11 4.41e-20
C189 Analog_0/V07 Analog_0/V03 0.21f
C190 Analog_0/V04 Analog_0/th01_0/m1_991_n1219# 3.84e-19
C191 therm_raw_0/input13/a_27_47# Analog_0/V07 1.72e-20
C192 Analog_0/V07 Analog_0/V01 1.12e-19
C193 therm_raw_0/net14 Vp 5.27e-20
C194 Analog_0/th08_0/m1_477_n803# Analog_0/V03 0.00463f
C195 Analog_0/th10_0/m1_536_174# Vin 1.1e-19
C196 Analog_0/th08_0/m1_477_n803# Analog_0/V01 2.53e-21
C197 Analog_0/V03 Analog_0/th01_0/m1_571_n501# 0.00963f
C198 Analog_0/th03_0/m1_890_n844# Analog_0/V02 0.0277f
C199 Vin Analog_0/V05 0.00184f
C200 Analog_0/th01_0/m1_571_n501# Analog_0/V01 1.33e-20
C201 Analog_0/th10_0/m1_536_174# Analog_0/V12 8.6e-19
C202 therm_raw_0/net2 therm_raw_0/net3 -1.42e-32
C203 therm_raw_0/_15_ therm_raw_0/b[3] -2.22e-34
C204 therm_raw_0/b[1] Analog_0/th12_0/m1_529_n42# 0.00163f
C205 Analog_0/V13 Vp 0.0659f
C206 therm_raw_0/b[3] Analog_0/th10_0/m1_536_174# 7.88e-21
C207 Analog_0/V14 Vin 0.0125f
C208 Analog_0/V09 Analog_0/th15_0/m1_849_n157# 0.0503f
C209 Analog_0/V07 Vp 8.84e-19
C210 Analog_0/V13 Analog_0/V15 0.154f
C211 Analog_0/V09 Analog_0/th15_0/m1_597_n912# 2.88e-21
C212 Analog_0/V14 Analog_0/V12 0.108f
C213 therm_raw_0/_19_ Vp 4.88e-19
C214 Analog_0/V14 Analog_0/V11 0.308f
C215 Analog_0/V06 Vp 0.0293f
C216 therm_raw_0/b[3] Analog_0/V14 1.02e-19
C217 therm_raw_0/input5/a_381_47# Vp -2.84e-32
C218 Analog_0/th04_0/m1_892_n998# Analog_0/V02 0.0341f
C219 Analog_0/V02 Analog_0/th02_0/m1_983_133# 0.0567f
C220 Analog_0/V07 Analog_0/V08 0.46f
C221 Analog_0/th06_0/m1_904_n796# Analog_0/V07 9.64e-20
C222 Analog_0/V08 Analog_0/th08_0/m1_477_n803# 0.00722f
C223 therm_raw_0/_01_ Vp 1.29e-19
C224 therm_raw_0/net3 Analog_0/V12 7.96e-21
C225 Analog_0/V08 Analog_0/V06 0.0717f
C226 Analog_0/V13 Analog_0/th13_0/m1_831_275# 0.0128f
C227 Analog_0/V07 Analog_0/th07_0/m1_808_n892# 0.0154f
C228 Analog_0/th06_0/m1_904_n796# Analog_0/V06 0.0113f
C229 Analog_0/V03 Analog_0/V02 0.0621f
C230 Vp therm_raw_0/net5 5.68e-32
C231 Analog_0/V12 therm_raw_0/b[1] 0.00221f
C232 Analog_0/V02 Analog_0/V01 -0.0388f
C233 Analog_0/V11 therm_raw_0/b[1] 0.0644f
C234 Analog_0/th07_0/m1_808_n892# Analog_0/V06 9.18e-20
C235 Analog_0/V04 Vn 1.72f
C236 Analog_0/th04_0/m1_892_n998# Vn 0.832f
C237 Analog_0/th04_0/m1_620_n488# Vn 0.0632f
C238 Analog_0/th11_0/m1_705_187# Vn 0.602f
C239 Analog_0/V11 Vn 2.18f
C240 Vin Vn 15f
C241 Analog_0/th11_0/m1_577_n654# Vn 0.286f
C242 Analog_0/V06 Vn 1.67f
C243 Analog_0/th06_0/m1_904_n796# Vn 0.495f
C244 Analog_0/th13_0/m1_831_275# Vn 1.05f
C245 Analog_0/V13 Vn 2.83f
C246 Analog_0/th13_0/m1_559_n458# Vn 0.286f
C247 Analog_0/th08_0/m1_477_n803# Vn 0.577f
C248 Analog_0/V08 Vn 1.72f
C249 Analog_0/V15 Vn 2.68f
C250 Analog_0/th15_0/m1_849_n157# Vn 1.28f
C251 Analog_0/th15_0/m1_597_n912# Vn 0.19f
C252 Analog_0/th01_0/m1_991_n1219# Vn 1.24f
C253 Analog_0/V01 Vn 2.54f
C254 Analog_0/th01_0/m1_571_n501# Vn 0.194f
C255 Analog_0/th15_0/Vin Vn 5.76f
C256 Analog_0/V03 Vn 2.11f
C257 Analog_0/th03_0/m1_890_n844# Vn 1.05f
C258 Analog_0/th03_0/m1_638_n591# Vn 0.224f
C259 Analog_0/th10_0/m1_536_174# Vn 0.825f
C260 Analog_0/V10 Vn 1.54f
C261 Analog_0/th10_0/m1_502_n495# Vn 0.145f
C262 Analog_0/th05_0/m1_752_n794# Vn 0.788f
C263 Analog_0/V05 Vn 2.13f
C264 Analog_0/th12_0/m1_529_n42# Vn 0.861f
C265 Analog_0/V12 Vn 1.91f
C266 Analog_0/th12_0/m1_394_n856# Vn 0.215f
C267 Analog_0/th07_0/m1_808_n892# Vn 0.506f
C268 Analog_0/V07 Vn 2.1f
C269 Analog_0/th14_0/m1_891_419# Vn 1.47f
C270 Analog_0/V14 Vn 1.56f
C271 Analog_0/th14_0/m1_641_n318# Vn 0.241f
C272 Analog_0/th09_0/m1_485_n505# Vn 1.18f
C273 Analog_0/V09 Vn 5.22f
C274 Analog_0/th09_0/m1_962_372# Vn 0.118f
C275 Analog_0/V02 Vn 3.73f
C276 Analog_0/th02_0/m1_983_133# Vn 1.44f
C277 Analog_0/th02_0/m1_571_144# Vn 0.252f
C278 therm_raw_0/_04_ Vn 0.339f
C279 therm_raw_0/_03_ Vn 0.36f
C280 therm_raw_0/net10 Vn 0.458f
C281 therm_raw_0/_30_/a_109_53# Vn 0.159f
C282 therm_raw_0/_30_/a_215_297# Vn 0.142f
C283 therm_raw_0/_05_ Vn 0.152f
C284 therm_raw_0/net8 Vn 0.386f
C285 therm_raw_0/_31_/a_285_297# Vn 0.00137f
C286 therm_raw_0/_31_/a_35_297# Vn 0.255f
C287 therm_raw_0/_32_/a_27_47# Vn 0.175f
C288 therm_raw_0/_50_/a_343_93# Vn 0.172f
C289 therm_raw_0/_50_/a_223_47# Vn 0.141f
C290 therm_raw_0/_50_/a_27_47# Vn 0.259f
C291 therm_raw_0/_07_ Vn 0.288f
C292 therm_raw_0/_06_ Vn 0.819f
C293 therm_raw_0/net13 Vn 0.379f
C294 therm_raw_0/_33_/a_209_311# Vn 0.143f
C295 therm_raw_0/_33_/a_109_93# Vn 0.158f
C296 therm_raw_0/_08_ Vn 0.131f
C297 therm_raw_0/net12 Vn 0.529f
C298 therm_raw_0/_34_/a_285_47# Vn 0.0174f
C299 therm_raw_0/_34_/a_47_47# Vn 0.199f
C300 therm_raw_0/_23_ Vn 0.106f
C301 therm_raw_0/input15/a_27_47# Vn 0.208f
C302 therm_raw_0/_09_ Vn 0.149f
C303 therm_raw_0/_35_/a_489_413# Vn 0.0254f
C304 therm_raw_0/_35_/a_226_47# Vn 0.162f
C305 therm_raw_0/_35_/a_76_199# Vn 0.141f
C306 therm_raw_0/_24_ Vn 0.135f
C307 therm_raw_0/_12_ Vn 0.387f
C308 therm_raw_0/_52_/a_250_297# Vn 0.0278f
C309 therm_raw_0/_52_/a_93_21# Vn 0.151f
C310 therm_raw_0/_10_ Vn 0.643f
C311 therm_raw_0/_36_/a_27_47# Vn 0.175f
C312 therm_raw_0/input14/a_27_47# Vn 0.208f
C313 therm_raw_0/_53_/a_29_53# Vn 0.18f
C314 therm_raw_0/_11_ Vn 0.267f
C315 therm_raw_0/_37_/a_27_47# Vn 0.175f
C316 therm_raw_0/input13/a_27_47# Vn 0.208f
C317 therm_raw_0/net18 Vn 0.207f
C318 therm_raw_0/_25_ Vn 0.191f
C319 therm_raw_0/_54_/a_75_212# Vn 0.21f
C320 therm_raw_0/_38_/a_27_47# Vn 0.175f
C321 therm_raw_0/net19 Vn 0.177f
C322 therm_raw_0/_22_ Vn 0.216f
C323 therm_raw_0/_14_ Vn 0.228f
C324 therm_raw_0/_15_ Vn 0.338f
C325 therm_raw_0/_55_/a_217_297# Vn 0.00117f
C326 therm_raw_0/_55_/a_80_21# Vn 0.21f
C327 therm_raw_0/input12/a_27_47# Vn 0.208f
C328 therm_raw_0/net9 Vn 0.306f
C329 therm_raw_0/input9/a_75_212# Vn 0.21f
C330 therm_raw_0/_39_/a_285_47# Vn 0.0174f
C331 therm_raw_0/_39_/a_47_47# Vn 0.199f
C332 therm_raw_0/net11 Vn 0.771f
C333 therm_raw_0/input11/a_27_47# Vn 0.208f
C334 therm_raw_0/input8/a_27_47# Vn 0.208f
C335 therm_raw_0/input10/a_27_47# Vn 0.208f
C336 therm_raw_0/net7 Vn 0.462f
C337 therm_raw_0/input7/a_27_47# Vn 0.208f
C338 therm_raw_0/input6/a_27_47# Vn 0.208f
C339 therm_raw_0/net5 Vn 0.842f
C340 therm_raw_0/input5/a_841_47# Vn 0.0929f
C341 therm_raw_0/input5/a_664_47# Vn 0.13f
C342 therm_raw_0/input5/a_558_47# Vn 0.164f
C343 therm_raw_0/input5/a_381_47# Vn 0.11f
C344 therm_raw_0/input5/a_62_47# Vn 0.169f
C345 therm_raw_0/input4/a_75_212# Vn 0.21f
C346 therm_raw_0/input3/a_27_47# Vn 0.208f
C347 therm_raw_0/net2 Vn 0.668f
C348 therm_raw_0/input2/a_27_47# Vn 0.208f
C349 therm_raw_0/net1 Vn 0.342f
C350 Vp Vn 84.8f
C351 therm_raw_0/input1/a_75_212# Vn 0.21f
C352 therm_raw_0/b[3] Vn 0.423f
C353 therm_raw_0/output19/a_27_47# Vn 0.543f
C354 therm_raw_0/b[2] Vn 0.515f
C355 therm_raw_0/output18/a_27_47# Vn 0.543f
C356 therm_raw_0/b[1] Vn 0.483f
C357 therm_raw_0/net17 Vn 0.173f
C358 therm_raw_0/output17/a_27_47# Vn 0.543f
C359 therm_raw_0/_41_/a_59_75# Vn 0.177f
C360 therm_raw_0/b[0] Vn 0.528f
C361 therm_raw_0/output16/a_27_47# Vn 0.543f
C362 therm_raw_0/_16_ Vn 0.125f
C363 therm_raw_0/_42_/a_209_311# Vn 0.143f
C364 therm_raw_0/_42_/a_109_93# Vn 0.158f
C365 therm_raw_0/_17_ Vn 0.251f
C366 therm_raw_0/_00_ Vn 0.377f
C367 therm_raw_0/_43_/a_193_413# Vn 0.136f
C368 therm_raw_0/_43_/a_27_47# Vn 0.224f
C369 therm_raw_0/net6 Vn 0.532f
C370 therm_raw_0/net4 Vn 0.324f
C371 therm_raw_0/_26_/a_29_53# Vn 0.18f
C372 therm_raw_0/_01_ Vn 0.15f
C373 therm_raw_0/net14 Vn 0.516f
C374 therm_raw_0/net3 Vn 0.464f
C375 therm_raw_0/net15 Vn 0.452f
C376 therm_raw_0/_27_/a_27_297# Vn 0.163f
C377 therm_raw_0/_18_ Vn 0.143f
C378 therm_raw_0/_44_/a_250_297# Vn 0.0278f
C379 therm_raw_0/_44_/a_93_21# Vn 0.151f
C380 therm_raw_0/net16 Vn 0.231f
C381 therm_raw_0/_13_ Vn 0.133f
C382 therm_raw_0/_45_/a_193_297# Vn 0.0011f
C383 therm_raw_0/_45_/a_109_297# Vn 7.11e-19
C384 therm_raw_0/_45_/a_27_47# Vn 0.216f
C385 therm_raw_0/_29_/a_29_53# Vn 0.18f
C386 therm_raw_0/_19_ Vn 0.118f
C387 therm_raw_0/_47_/a_299_297# Vn 0.0348f
C388 therm_raw_0/_47_/a_81_21# Vn 0.147f
C389 therm_raw_0/_48_/a_27_47# Vn 0.177f
C390 therm_raw_0/_21_ Vn 0.29f
C391 therm_raw_0/_20_ Vn 0.238f
C392 therm_raw_0/_02_ Vn 0.453f
C393 therm_raw_0/_49_/a_201_297# Vn 0.00345f
C394 therm_raw_0/_49_/a_75_199# Vn 0.205f
.ends

