magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 2572 29 2578
rect -29 2538 -17 2572
rect -29 2532 29 2538
rect -29 -2538 29 -2532
rect -29 -2572 -17 -2538
rect -29 -2578 29 -2572
<< pwell >>
rect -211 -2710 211 2710
<< nmos >>
rect -15 -2500 15 2500
<< ndiff >>
rect -73 2488 -15 2500
rect -73 -2488 -61 2488
rect -27 -2488 -15 2488
rect -73 -2500 -15 -2488
rect 15 2488 73 2500
rect 15 -2488 27 2488
rect 61 -2488 73 2488
rect 15 -2500 73 -2488
<< ndiffc >>
rect -61 -2488 -27 2488
rect 27 -2488 61 2488
<< psubdiff >>
rect -175 2640 -79 2674
rect 79 2640 175 2674
rect -175 2578 -141 2640
rect 141 2578 175 2640
rect -175 -2640 -141 -2578
rect 141 -2640 175 -2578
rect -175 -2674 -79 -2640
rect 79 -2674 175 -2640
<< psubdiffcont >>
rect -79 2640 79 2674
rect -175 -2578 -141 2578
rect 141 -2578 175 2578
rect -79 -2674 79 -2640
<< poly >>
rect -33 2572 33 2588
rect -33 2538 -17 2572
rect 17 2538 33 2572
rect -33 2522 33 2538
rect -15 2500 15 2522
rect -15 -2522 15 -2500
rect -33 -2538 33 -2522
rect -33 -2572 -17 -2538
rect 17 -2572 33 -2538
rect -33 -2588 33 -2572
<< polycont >>
rect -17 2538 17 2572
rect -17 -2572 17 -2538
<< locali >>
rect -175 2640 -79 2674
rect 79 2640 175 2674
rect -175 2578 -141 2640
rect 141 2578 175 2640
rect -33 2538 -17 2572
rect 17 2538 33 2572
rect -61 2488 -27 2504
rect -61 -2504 -27 -2488
rect 27 2488 61 2504
rect 27 -2504 61 -2488
rect -33 -2572 -17 -2538
rect 17 -2572 33 -2538
rect -175 -2640 -141 -2578
rect 141 -2640 175 -2578
rect -175 -2674 -79 -2640
rect 79 -2674 175 -2640
<< viali >>
rect -17 2538 17 2572
rect -61 -2488 -27 2488
rect 27 -2488 61 2488
rect -17 -2572 17 -2538
<< metal1 >>
rect -29 2572 29 2578
rect -29 2538 -17 2572
rect 17 2538 29 2572
rect -29 2532 29 2538
rect -67 2488 -21 2500
rect -67 -2488 -61 2488
rect -27 -2488 -21 2488
rect -67 -2500 -21 -2488
rect 21 2488 67 2500
rect 21 -2488 27 2488
rect 61 -2488 67 2488
rect 21 -2500 67 -2488
rect -29 -2538 29 -2532
rect -29 -2572 -17 -2538
rect 17 -2572 29 -2538
rect -29 -2578 29 -2572
<< properties >>
string FIXED_BBOX -158 -2657 158 2657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 25.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
