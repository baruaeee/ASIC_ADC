magic
tech sky130A
magscale 1 2
timestamp 1704313364
use th13  x1
timestamp 1704313364
transform 1 0 53 0 1 1800
box 240 -1200 2062 556
<< end >>
