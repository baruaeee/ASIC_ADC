magic
tech sky130A
magscale 1 2
timestamp 1706270854
<< psubdiff >>
rect 1839 -1412 1925 -1378
<< locali >>
rect 1493 -66 1522 -32
rect 484 -444 518 -413
rect 1837 -1412 1891 -1378
<< viali >>
rect 1459 -66 1493 -32
rect 484 -479 519 -444
rect 1891 -1412 1925 -1378
<< metal1 >>
rect 1418 -32 1518 6
rect 1418 -66 1459 -32
rect 1493 -35 1518 -32
rect 1493 -66 1519 -35
rect 1418 -94 1519 -66
rect 571 -287 631 -227
rect 1355 -253 1420 -225
rect 1355 -287 1421 -253
rect 472 -444 531 -438
rect 472 -479 484 -444
rect 519 -479 531 -444
rect 472 -485 531 -479
rect 571 -457 605 -287
rect 1046 -370 1096 -346
rect 1040 -422 1046 -370
rect 1098 -422 1104 -370
rect 482 -525 517 -485
rect 571 -501 607 -457
rect 433 -560 517 -525
rect 573 -527 607 -501
rect 433 -787 468 -560
rect 573 -561 1289 -527
rect 1255 -739 1289 -561
rect 1387 -571 1421 -287
rect 1485 -333 1519 -94
rect 1596 -184 1662 -122
rect 1567 -333 1601 -285
rect 1485 -336 1601 -333
rect 1485 -370 1604 -336
rect 1657 -349 1691 -285
rect 1567 -467 1601 -370
rect 1657 -383 1925 -349
rect 1657 -451 1691 -383
rect 1505 -571 1661 -563
rect 1387 -597 1661 -571
rect 1387 -605 1539 -597
rect 1254 -787 1289 -739
rect 433 -851 501 -787
rect 1223 -821 1289 -787
rect 1223 -851 1288 -821
rect 433 -900 468 -851
rect 433 -935 895 -900
rect 402 -1066 454 -1060
rect 340 -1118 402 -1082
rect 1505 -1074 1539 -605
rect 1891 -640 1925 -383
rect 1868 -740 1968 -640
rect 1933 -872 1967 -740
rect 1685 -906 1967 -872
rect 1686 -938 1748 -906
rect 340 -1124 454 -1118
rect 1113 -1108 1640 -1074
rect 340 -1182 440 -1124
rect 1113 -1185 1147 -1108
rect 545 -1268 551 -1216
rect 603 -1268 628 -1216
rect 991 -1219 1251 -1185
rect 548 -1270 628 -1268
rect 1059 -1273 1094 -1271
rect 875 -1308 1257 -1273
rect 1402 -1278 1458 -1214
rect 1700 -1265 1734 -1264
rect 1683 -1299 1753 -1265
rect 1059 -1376 1094 -1308
rect 1700 -1376 1735 -1299
rect 1059 -1379 1735 -1376
rect 1860 -1378 1960 -1344
rect 1860 -1379 1891 -1378
rect 1059 -1411 1891 -1379
rect 1700 -1412 1891 -1411
rect 1925 -1412 1960 -1378
rect 1700 -1413 1960 -1412
rect 1860 -1444 1960 -1413
<< via1 >>
rect 1046 -422 1098 -370
rect 402 -1118 454 -1066
rect 551 -1268 603 -1216
<< metal2 >>
rect 1046 -370 1098 -364
rect 1098 -422 1353 -419
rect 1046 -428 1353 -422
rect 1055 -453 1353 -428
rect 1319 -995 1353 -453
rect 411 -1029 1353 -995
rect 411 -1066 445 -1029
rect 396 -1118 402 -1066
rect 454 -1118 460 -1066
rect 560 -1210 594 -1029
rect 551 -1216 603 -1210
rect 551 -1274 603 -1268
use sky130_fd_pr__nfet_01v8_SHU4BF  XM0
timestamp 1706204487
transform 0 -1 1019 1 0 -1245
box -211 -563 211 563
use sky130_fd_pr__pfet_01v8_HE9GT9  XM1
timestamp 1706204487
transform 1 0 994 0 1 -257
box -546 -261 546 261
use sky130_fd_pr__nfet_01v8_LHD8GA  XM2
timestamp 1706204487
transform 1 0 862 0 1 -820
box -546 -252 546 252
use sky130_fd_pr__pfet_01v8_XJP3BL  XM3
timestamp 1706204487
transform -1 0 1629 0 -1 -365
box -211 -369 211 369
use sky130_fd_pr__nfet_01v8_LH5FDA  XM4
timestamp 1706211875
transform 0 -1 1716 -1 0 -1102
box -260 -252 346 252
<< labels >>
flabel metal1 1860 -1444 1960 -1344 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 1868 -740 1968 -640 0 FreeSans 256 0 0 0 V01
port 2 nsew
flabel metal1 1418 -94 1518 6 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 340 -1182 440 -1082 0 FreeSans 256 0 0 0 Vin
port 1 nsew
<< end >>
