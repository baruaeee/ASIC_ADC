** sch_path: /home/exotic/Desktop/ASIC_ADC/xschem/Transient_Analysis_Inverter_sym_test_banch.sch
.subckt Transient_Analysis_Inverter_sym_test_banch Vin Vout
*.PININFO Vin:I Vout:O
VDD VDD GND 1.8
.save i(vdd)
Vin Vin GND pulse(0 1.8 0ns 1ns 1ns 5ns 10ns)
.save i(vin)
x1 VDD Vin Vout GND make_symbol_Inverter
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.save all





.tran 1n 30n
.control
run
set color0=white
set color1=black
plot Vin Vout
set xbrushwidth=3
.save all
.endc
.end


**** end user architecture code
.ends

* expanding   symbol:  make_symbol_Inverter.sym # of pins=4
** sym_path: /home/exotic/Desktop/ASIC_ADC/xschem/make_symbol_Inverter.sym
** sch_path: /home/exotic/Desktop/ASIC_ADC/xschem/make_symbol_Inverter.sch
.subckt make_symbol_Inverter Vdd Vin Vout GND
*.PININFO Vin:I Vout:O Vdd:B GND:B
XM1 Vout Vin Vdd net1 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 Vout Vin GND net2 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
