* NGSPICE file created from th01_1.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_9DPZTU w_n291_n261# a_n153_n42# a_n95_n139# a_95_n42#
+ VSUBS
X0 a_95_n42# a_n95_n139# a_n153_n42# w_n291_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.95
C0 a_n95_n139# w_n291_n261# 0.419f
C1 a_n95_n139# a_n153_n42# 0.014f
C2 w_n291_n261# a_n153_n42# 0.0499f
C3 a_n95_n139# a_95_n42# 0.014f
C4 w_n291_n261# a_95_n42# 0.0499f
C5 a_95_n42# a_n153_n42# 0.0249f
C6 a_95_n42# VSUBS 0.0313f
C7 a_n153_n42# VSUBS 0.0313f
C8 a_n95_n139# VSUBS 0.289f
C9 w_n291_n261# VSUBS 1.36f
.ends

.subckt sky130_fd_pr__nfet_01v8_586EUA a_n97_n95# a_n199_n269# a_n39_n183# a_39_n95#
X0 a_39_n95# a_n39_n183# a_n97_n95# a_n199_n269# sky130_fd_pr__nfet_01v8 ad=0.275 pd=2.48 as=0.275 ps=2.48 w=0.95 l=0.39
C0 a_n97_n95# a_n39_n183# 0.0127f
C1 a_n97_n95# a_39_n95# 0.1f
C2 a_n39_n183# a_39_n95# 0.0127f
C3 a_39_n95# a_n199_n269# 0.135f
C4 a_n97_n95# a_n199_n269# 0.135f
C5 a_n39_n183# a_n199_n269# 0.381f
.ends

.subckt sky130_fd_pr__nfet_01v8_PJBF84 a_n248_n222# a_n146_n48# a_88_n48# a_n88_n136#
X0 a_88_n48# a_n88_n136# a_n146_n48# a_n248_n222# sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.54 as=0.139 ps=1.54 w=0.48 l=0.88
C0 a_n146_n48# a_n88_n136# 0.0146f
C1 a_n146_n48# a_88_n48# 0.03f
C2 a_n88_n136# a_88_n48# 0.0146f
C3 a_88_n48# a_n248_n222# 0.088f
C4 a_n146_n48# a_n248_n222# 0.088f
C5 a_n88_n136# a_n248_n222# 0.649f
.ends

.subckt sky130_fd_pr__pfet_01v8_RVEGTV a_n69_n175# a_n127_n78# w_n265_n297# a_69_n78#
+ VSUBS
X0 a_69_n78# a_n69_n175# a_n127_n78# w_n265_n297# sky130_fd_pr__pfet_01v8 ad=0.226 pd=2.14 as=0.226 ps=2.14 w=0.78 l=0.69
C0 a_n69_n175# w_n265_n297# 0.338f
C1 a_n69_n175# a_n127_n78# 0.0173f
C2 w_n265_n297# a_n127_n78# 0.0718f
C3 a_n69_n175# a_69_n78# 0.0173f
C4 w_n265_n297# a_69_n78# 0.0718f
C5 a_69_n78# a_n127_n78# 0.0574f
C6 a_69_n78# VSUBS 0.0474f
C7 a_n127_n78# VSUBS 0.0474f
C8 a_n69_n175# VSUBS 0.227f
C9 w_n265_n297# VSUBS 1.41f
.ends

.subckt th01 Vp Vin Vout m1_732_n84# Vn
XXM2 Vp Vp Vin m1_732_n84# Vn sky130_fd_pr__pfet_01v8_9DPZTU
XXM3 Vn Vn Vin m1_732_n84# sky130_fd_pr__nfet_01v8_586EUA
XXM4 Vn Vn Vout m1_732_n84# sky130_fd_pr__nfet_01v8_PJBF84
XXM5 m1_732_n84# Vp Vp Vout Vn sky130_fd_pr__pfet_01v8_RVEGTV
C0 Vn Vin 0.0827f
C1 Vn Vp 0.167f
C2 m1_732_n84# Vout 0.174f
C3 Vin Vout 1.54e-19
C4 Vin m1_732_n84# 0.174f
C5 Vp Vout 0.0895f
C6 Vp m1_732_n84# 0.305f
C7 Vin Vp 0.228f
C8 Vn Vout 0.0643f
C9 Vn m1_732_n84# 0.18f
C10 Vin 0 0.683f
C11 Vp 0 2.57f
C12 Vout 0 0.247f
C13 m1_732_n84# 0 0.96f
C14 Vn 0 0.0948f
.ends

.subckt sky130_fd_pr__pfet_01v8_4N47A3 w_n231_n369# a_n93_n150# a_35_n150# a_n35_n247#
+ VSUBS
X0 a_35_n150# a_n35_n247# a_n93_n150# w_n231_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.35
C0 a_n93_n150# a_35_n150# 0.166f
C1 w_n231_n369# a_n35_n247# 0.233f
C2 a_n93_n150# a_n35_n247# 0.0165f
C3 a_n35_n247# a_35_n150# 0.0165f
C4 w_n231_n369# a_n93_n150# 0.116f
C5 w_n231_n369# a_35_n150# 0.116f
C6 a_35_n150# VSUBS 0.0757f
C7 a_n93_n150# VSUBS 0.0757f
C8 a_n35_n247# VSUBS 0.141f
C9 w_n231_n369# VSUBS 1.52f
.ends

.subckt sky130_fd_pr__nfet_01v8_48YMBA a_n518_n42# a_460_n42# a_n620_n216# a_n460_n130#
X0 a_460_n42# a_n460_n130# a_n518_n42# a_n620_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=4.6
C0 a_n460_n130# a_n518_n42# 0.0236f
C1 a_460_n42# a_n518_n42# 0.00624f
C2 a_n460_n130# a_460_n42# 0.0236f
C3 a_460_n42# a_n620_n216# 0.0868f
C4 a_n518_n42# a_n620_n216# 0.0868f
C5 a_n460_n130# a_n620_n216# 2.69f
.ends

.subckt preamp Vp Vin Vn Vpamp
XXM0 Vpamp Vn Vpamp Vin Vpamp sky130_fd_pr__pfet_01v8_4N47A3
XXM1 Vp Vpamp Vpamp Vin sky130_fd_pr__nfet_01v8_48YMBA
C0 Vin Vn 0.0147f
C1 Vpamp Vp 0.0775f
C2 Vp Vn 0.0228f
C3 Vpamp Vn 0.213f
C4 Vp Vin 0.233f
C5 Vpamp Vin 0.488f
C6 Vpamp 0 1.57f
C7 Vp 0 0.377f
C8 Vin 0 2.67f
C9 Vn 0 0.247f
.ends

.subckt th01_1
Xx1 x2/Vp VSUBS x1/Vout x1/m1_732_n84# VSUBS th01
Xx2 x2/Vp x2/Vin VSUBS VSUBS preamp
C0 x2/Vp x2/Vin 0.173f
C1 x1/m1_732_n84# x2/Vin 0.0029f
C2 x1/Vout x2/Vin 8.58e-20
C3 VSUBS x2/Vp 0.156f
C4 x1/m1_732_n84# VSUBS 0.00347f
C5 VSUBS x1/Vout 1.44e-19
C6 VSUBS x2/Vin 0.00888f
C7 VSUBS 0 2.24f
C8 x2/Vin 0 2.67f
C9 x2/Vp 0 3.38f
C10 x1/Vout 0 0.247f
C11 x1/m1_732_n84# 0 0.96f
.ends

