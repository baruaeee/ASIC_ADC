** sch_path: /home/exotic/Desktop/ASIC_ADC/xschem/Vth_sch/Pre_layout/th04.sch
**.subckt th04 Vin Vout
*.ipin Vin
*.opin Vout
VDD VDD GND 1.8
Vin Vin GND pulse(0 0.2 0ns 1ns 1ns 5ns 10ns)
V_logic_high V_LH GND 1.25
V_logic_low V_LL GND 0.5
x1 VDD Vout Vin GND th04
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.save all





.dc Vin 0 1.8 0.01
*.tran 1n 30n
.control
run
set color0=white
set color1=black
plot Vin Vout V_LH V_LL
set xbrushwidth=3
.save all
.endc
.end


**** end user architecture code
**.ends

* NGSPICE file created from th04.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_42G4RD a_n80_n42# a_n33_n130# a_n182_n216# a_22_n42#
X0 a_22_n42# a_n33_n130# a_n80_n42# a_n182_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_n80_n42# a_22_n42# 0.0604f
C1 a_22_n42# a_n33_n130# 0.00866f
C2 a_n80_n42# a_n33_n130# 0.00866f
C3 a_22_n42# a_n182_n216# 0.0785f
C4 a_n80_n42# a_n182_n216# 0.0785f
C5 a_n33_n130# a_n182_n216# 0.341f
.ends

.subckt sky130_fd_pr__pfet_01v8_DDPLQ8 a_n77_n42# w_n215_n261# a_n33_n139# a_19_n42#
+ VSUBS
X0 a_19_n42# a_n33_n139# a_n77_n42# w_n215_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_19_n42# a_n77_n42# 0.0641f
C1 a_n33_n139# a_19_n42# 0.0127f
C2 a_n33_n139# a_n77_n42# 0.0127f
C3 a_19_n42# w_n215_n261# 0.0484f
C4 a_n77_n42# w_n215_n261# 0.0484f
C5 a_n33_n139# w_n215_n261# 0.234f
C6 a_19_n42# VSUBS 0.0275f
C7 a_n77_n42# VSUBS 0.0275f
C8 a_n33_n139# VSUBS 0.119f
C9 w_n215_n261# VSUBS 1.04f
.ends

.subckt sky130_fd_pr__nfet_01v8_VWP3K3 a_n33_n130# a_15_n42# a_n175_n216# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n42# a_15_n42# 0.0699f
C1 a_15_n42# a_n33_n130# 0.0209f
C2 a_n73_n42# a_n33_n130# 0.0209f
C3 a_15_n42# a_n175_n216# 0.0729f
C4 a_n73_n42# a_n175_n216# 0.0729f
C5 a_n33_n130# a_n175_n216# 0.338f
.ends

.subckt sky130_fd_pr__pfet_01v8_LZD9A4 a_n80_n42# a_22_n42# a_n33_n139# w_n218_n261#
+ VSUBS
X0 a_22_n42# a_n33_n139# a_n80_n42# w_n218_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_22_n42# a_n80_n42# 0.0604f
C1 a_n33_n139# a_22_n42# 0.0084f
C2 a_n33_n139# a_n80_n42# 0.0084f
C3 a_22_n42# w_n218_n261# 0.0496f
C4 a_n80_n42# w_n218_n261# 0.0496f
C5 a_n33_n139# w_n218_n261# 0.233f
C6 a_22_n42# VSUBS 0.0285f
C7 a_n80_n42# VSUBS 0.0285f
C8 a_n33_n139# VSUBS 0.122f
C9 w_n218_n261# VSUBS 1.06f
.ends

.subckt sky130_fd_pr__nfet_01v8_VRD6K3 a_n77_n42# a_n33_n130# a_19_n42# a_n179_n216#
X0 a_19_n42# a_n33_n130# a_n77_n42# a_n179_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_n77_n42# a_19_n42# 0.0641f
C1 a_19_n42# a_n33_n130# 0.0136f
C2 a_n77_n42# a_n33_n130# 0.0136f
C3 a_19_n42# a_n179_n216# 0.0763f
C4 a_n77_n42# a_n179_n216# 0.0763f
C5 a_n33_n130# a_n179_n216# 0.339f
.ends

.subckt th04 Vp V04 Vin Vn
XXM0 m1_960_n972# Vin Vn Vn sky130_fd_pr__nfet_01v8_42G4RD
XXM1 m1_397_n357# Vp Vin m1_960_n972# Vn sky130_fd_pr__pfet_01v8_DDPLQ8
XXM2 Vp m1_397_n357# Vn Vp sky130_fd_pr__nfet_01v8_VWP3K3
XXM3 Vp V04 m1_960_n972# Vp Vn sky130_fd_pr__pfet_01v8_LZD9A4
XXM4 V04 m1_960_n972# Vn Vn sky130_fd_pr__nfet_01v8_VRD6K3
C0 Vp Vin 0.103f
C1 Vin V04 5.12e-19
C2 Vin m1_397_n357# 0.109f
C3 Vp m1_960_n972# 0.257f
C4 Vin Vn 0.0911f
C5 V04 m1_960_n972# 0.39f
C6 m1_397_n357# m1_960_n972# 0.027f
C7 Vn m1_960_n972# 0.346f
C8 Vp V04 0.173f
C9 Vp m1_397_n357# 0.401f
C10 Vp Vn 0.228f
C11 V04 m1_397_n357# 0.0695f
C12 Vn V04 0.181f
C13 Vn m1_397_n357# 0.0588f
C14 Vin m1_960_n972# 0.395f
C15 Vin 0 0.599f
C16 m1_960_n972# 0 0.53f
C17 Vn 0 0.213f
C18 V04 0 0.324f
C19 m1_397_n357# 0 0.189f
C20 Vp 0 2.61f
.ends


.GLOBAL VDD
.GLOBAL GND
.GLOBAL V_LH
.GLOBAL V_LL
.end
