magic
tech sky130A
magscale 1 2
timestamp 1696359958
<< metal1 >>
rect 6246 3586 6446 3672
rect 6246 3468 6958 3586
rect 1142 3154 1492 3220
rect 6246 3218 6524 3468
rect 6834 3266 6958 3468
rect 6682 3236 6958 3266
rect 1142 2544 1240 3154
rect 6246 2914 6524 3156
rect 6682 3146 6854 3236
rect 6940 3146 6958 3236
rect 6682 3108 6958 3146
rect 6246 2804 7192 2914
rect 1142 2478 1492 2544
rect 6246 2540 6524 2804
rect 6682 2554 6958 2590
rect 1142 1868 1238 2478
rect 6246 2252 6524 2480
rect 6682 2464 6854 2554
rect 6940 2464 6958 2554
rect 6682 2432 6958 2464
rect 6834 2252 6958 2432
rect 6246 2112 6960 2252
rect 1142 1802 1488 1868
rect 6246 1864 6524 2112
rect 6836 1914 6960 2112
rect 768 1232 968 1428
rect 1142 1232 1236 1802
rect 6002 1542 6198 1806
rect 6682 1756 6960 1914
rect 7072 1542 7192 2804
rect 6002 1424 7194 1542
rect 768 1198 2090 1232
rect 768 294 850 1198
rect 1116 1076 1508 1160
rect 6992 1158 7192 1424
rect 6516 1076 7192 1158
rect 1116 776 1198 1076
rect 3028 776 3228 934
rect 1116 576 6972 776
rect 3028 574 3228 576
rect 768 260 2092 294
rect 768 -634 850 260
rect 1116 138 1508 222
rect 6898 220 6972 576
rect 6516 138 6972 220
rect 1116 -162 1198 138
rect 3028 -162 3228 -4
rect 6898 -162 6972 -160
rect 1116 -362 6972 -162
rect 3028 -364 3228 -362
rect 768 -668 2094 -634
rect 1114 -790 1500 -706
rect 6898 -708 6972 -362
rect 6518 -790 6972 -708
rect 1114 -1090 1196 -790
rect 3028 -1090 3230 -930
rect 1114 -1102 3230 -1090
rect 1114 -1290 3228 -1102
<< via1 >>
rect 6854 3146 6940 3236
rect 6854 2464 6940 2554
<< metal2 >>
rect 6846 3236 6950 3242
rect 6846 3146 6854 3236
rect 6940 3146 6950 3236
rect 6846 2554 6950 3146
rect 6846 2464 6854 2554
rect 6940 2464 6950 2554
rect 6846 2446 6950 2464
use sky130_fd_pr__pfet_01v8_KGSDF3  XM7
timestamp 1696298453
transform 0 1 4033 -1 0 1835
box -211 -2719 211 2719
use sky130_fd_pr__nfet_01v8_YYPCPJ  XM8
timestamp 1696298453
transform 1 0 4012 0 1 -748
box -2696 -252 2696 252
use sky130_fd_pr__nfet_01v8_YYPCPJ  XM9
timestamp 1696298453
transform 1 0 4008 0 1 180
box -2696 -252 2696 252
use sky130_fd_pr__nfet_01v8_YYPCPJ  XM10
timestamp 1696298453
transform 1 0 4008 0 1 1116
box -2696 -252 2696 252
use sky130_fd_pr__pfet_01v8_KGSDF3  XM11
timestamp 1696298453
transform 0 1 4033 -1 0 2511
box -211 -2719 211 2719
use sky130_fd_pr__pfet_01v8_KGSDF3  XM12
timestamp 1696298453
transform 0 1 4033 -1 0 3187
box -211 -2719 211 2719
<< labels >>
flabel metal1 3028 -1290 3228 -1090 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 768 1228 968 1428 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 6992 1342 7192 1542 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 6246 3472 6446 3672 0 FreeSans 256 0 0 0 Vp
port 0 nsew
<< end >>
