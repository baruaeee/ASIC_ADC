** sch_path: /home/exotic/Desktop/ASIC_ADC/xschem/Vth_sch/test_ngspice/test_script.sch
**.subckt test_script Vin Vin Vout
*.ipin Vin
*.ipin Vin
*.opin Vout
VDD VDD GND 1.8
Vin Vin GND 0.621200000V

XM1 Vout Vin VDD net1 sky130_fd_pr__pfet_01v8 L=0.7100000000000004 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout Vin GND net2 sky130_fd_pr__nfet_01v8 L=0.153 W=2.315 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1

V_logic_high V_LH GND 1.25
V_logic_low V_LL GND 0.5
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.save all





.control
op
*run
.endc
.end


**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.GLOBAL V_LH
.GLOBAL V_LL
.end
