magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_s >>
rect 546 1069 581 1087
rect 510 1068 581 1069
rect 1800 1070 1858 1076
rect 510 583 580 1068
rect 1800 1036 1812 1070
rect 1800 1030 1858 1036
rect 692 1000 750 1006
rect 692 966 704 1000
rect 692 960 750 966
rect 862 963 896 981
rect 1654 963 1688 981
rect 862 927 932 963
rect 879 893 950 927
rect 692 666 750 672
rect 692 632 704 666
rect 692 626 750 632
rect 510 547 563 583
rect 879 530 949 893
rect 879 494 932 530
rect 1618 477 1688 963
rect 1800 560 1858 566
rect 1800 526 1812 560
rect 1800 520 1858 526
rect 1618 441 1671 477
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_VZ9GC6  XM1
timestamp 1703732895
transform 1 0 1275 0 1 702
box -396 -261 396 261
use sky130_fd_pr__nfet_01v8_ATLS57  XM3
timestamp 1703732895
transform 1 0 1829 0 1 798
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_PZD9SE  XM7
timestamp 1703732895
transform 1 0 255 0 1 808
box -308 -261 308 261
use sky130_fd_pr__nfet_01v8_UNLS3X  XM10
timestamp 1703732895
transform 1 0 721 0 1 816
box -211 -322 211 322
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
