magic
tech sky130A
magscale 1 2
timestamp 1704501257
<< error_p >>
rect -29 1181 29 1187
rect -29 1147 -17 1181
rect -29 1141 29 1147
rect -29 -1147 29 -1141
rect -29 -1181 -17 -1147
rect -29 -1187 29 -1181
<< nwell >>
rect -214 -1319 214 1319
<< pmos >>
rect -18 -1100 18 1100
<< pdiff >>
rect -76 1088 -18 1100
rect -76 -1088 -64 1088
rect -30 -1088 -18 1088
rect -76 -1100 -18 -1088
rect 18 1088 76 1100
rect 18 -1088 30 1088
rect 64 -1088 76 1088
rect 18 -1100 76 -1088
<< pdiffc >>
rect -64 -1088 -30 1088
rect 30 -1088 64 1088
<< nsubdiff >>
rect -178 1249 -82 1283
rect 82 1249 178 1283
rect -178 1187 -144 1249
rect 144 1187 178 1249
rect -178 -1249 -144 -1187
rect 144 -1249 178 -1187
rect -178 -1283 -82 -1249
rect 82 -1283 178 -1249
<< nsubdiffcont >>
rect -82 1249 82 1283
rect -178 -1187 -144 1187
rect 144 -1187 178 1187
rect -82 -1283 82 -1249
<< poly >>
rect -33 1181 33 1197
rect -33 1147 -17 1181
rect 17 1147 33 1181
rect -33 1131 33 1147
rect -18 1100 18 1131
rect -18 -1131 18 -1100
rect -33 -1147 33 -1131
rect -33 -1181 -17 -1147
rect 17 -1181 33 -1147
rect -33 -1197 33 -1181
<< polycont >>
rect -17 1147 17 1181
rect -17 -1181 17 -1147
<< locali >>
rect -178 1249 -82 1283
rect 82 1249 178 1283
rect -178 1187 -144 1249
rect 144 1187 178 1249
rect -33 1147 -17 1181
rect 17 1147 33 1181
rect -64 1088 -30 1104
rect -64 -1104 -30 -1088
rect 30 1088 64 1104
rect 30 -1104 64 -1088
rect -33 -1181 -17 -1147
rect 17 -1181 33 -1147
rect -178 -1249 -144 -1187
rect 144 -1249 178 -1187
rect -178 -1283 -82 -1249
rect 82 -1283 178 -1249
<< viali >>
rect -17 1147 17 1181
rect -64 -1088 -30 1088
rect 30 -1088 64 1088
rect -17 -1181 17 -1147
<< metal1 >>
rect -29 1181 29 1187
rect -29 1147 -17 1181
rect 17 1147 29 1181
rect -29 1141 29 1147
rect -70 1088 -24 1100
rect -70 -1088 -64 1088
rect -30 -1088 -24 1088
rect -70 -1100 -24 -1088
rect 24 1088 70 1100
rect 24 -1088 30 1088
rect 64 -1088 70 1088
rect 24 -1100 70 -1088
rect -29 -1147 29 -1141
rect -29 -1181 -17 -1147
rect 17 -1181 29 -1147
rect -29 -1187 29 -1181
<< properties >>
string FIXED_BBOX -161 -1266 161 1266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 11.0 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
