magic
tech sky130A
magscale 1 2
timestamp 1704389634
<< nwell >>
rect -308 -261 308 261
<< pmos >>
rect -112 -42 112 42
<< pdiff >>
rect -170 30 -112 42
rect -170 -30 -158 30
rect -124 -30 -112 30
rect -170 -42 -112 -30
rect 112 30 170 42
rect 112 -30 124 30
rect 158 -30 170 30
rect 112 -42 170 -30
<< pdiffc >>
rect -158 -30 -124 30
rect 124 -30 158 30
<< nsubdiff >>
rect -272 191 -176 225
rect 176 191 272 225
rect -272 129 -238 191
rect 238 129 272 191
rect -272 -191 -238 -129
rect 238 -191 272 -129
rect -272 -225 -176 -191
rect 176 -225 272 -191
<< nsubdiffcont >>
rect -176 191 176 225
rect -272 -129 -238 129
rect 238 -129 272 129
rect -176 -225 176 -191
<< poly >>
rect -112 123 112 139
rect -112 89 -96 123
rect 96 89 112 123
rect -112 42 112 89
rect -112 -89 112 -42
rect -112 -123 -96 -89
rect 96 -123 112 -89
rect -112 -139 112 -123
<< polycont >>
rect -96 89 96 123
rect -96 -123 96 -89
<< locali >>
rect -272 191 -176 225
rect 176 191 272 225
rect -272 129 -238 191
rect 238 129 272 191
rect -112 89 -96 123
rect 96 89 112 123
rect -158 30 -124 46
rect -158 -46 -124 -30
rect 124 30 158 46
rect 124 -46 158 -30
rect -112 -123 -96 -89
rect 96 -123 112 -89
rect -272 -191 -238 -129
rect 238 -191 272 -129
rect -272 -225 -176 -191
rect 176 -225 272 -191
<< viali >>
rect -96 89 96 123
rect -158 -30 -124 30
rect 124 -30 158 30
rect -96 -123 96 -89
<< metal1 >>
rect -108 123 108 129
rect -108 89 -96 123
rect 96 89 108 123
rect -108 83 108 89
rect -164 30 -118 42
rect -164 -30 -158 30
rect -124 -30 -118 30
rect -164 -42 -118 -30
rect 118 30 164 42
rect 118 -30 124 30
rect 158 -30 164 30
rect 118 -42 164 -30
rect -108 -89 108 -83
rect -108 -123 -96 -89
rect 96 -123 108 -89
rect -108 -129 108 -123
<< properties >>
string FIXED_BBOX -255 -208 255 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 1.12 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
