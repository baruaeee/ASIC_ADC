magic
tech sky130A
magscale 1 2
timestamp 1706270854
<< nsubdiff >>
rect 1275 94 1327 128
<< locali >>
rect 642 168 667 202
rect 1300 94 1326 128
rect 1610 -1034 1644 -959
<< viali >>
rect 607 168 642 203
rect 1265 94 1300 129
rect 1610 -1069 1645 -1034
<< metal1 >>
rect 601 203 648 215
rect 601 168 607 203
rect 642 168 648 203
rect 601 162 648 168
rect 576 110 582 162
rect 634 156 648 162
rect 634 110 640 156
rect 1196 141 1296 204
rect 1196 129 1306 141
rect 1196 104 1265 129
rect 1259 94 1265 104
rect 1300 94 1306 129
rect 1259 82 1306 94
rect 638 -57 743 7
rect 1041 -32 1182 3
rect 1041 -57 1076 -32
rect 638 -527 672 -57
rect 864 -146 916 -118
rect 858 -198 864 -146
rect 916 -198 922 -146
rect 1147 -301 1182 -32
rect 1259 -129 1293 82
rect 1374 -20 1436 42
rect 1343 -129 1377 -93
rect 1259 -130 1377 -129
rect 1259 -163 1379 -130
rect 1280 -164 1379 -163
rect 1435 -133 1469 -103
rect 1343 -205 1377 -164
rect 1435 -167 1562 -133
rect 1435 -211 1469 -167
rect 1145 -335 1435 -301
rect 1145 -336 1434 -335
rect 1316 -342 1434 -336
rect 765 -442 771 -390
rect 823 -442 829 -390
rect 971 -481 1058 -447
rect 977 -489 1058 -481
rect 638 -591 701 -527
rect 1009 -553 1058 -489
rect 1024 -587 1058 -553
rect 1316 -713 1351 -342
rect 1055 -715 1351 -713
rect 1528 -476 1562 -167
rect 1528 -576 1630 -476
rect 1055 -745 1417 -715
rect 890 -747 1417 -745
rect 890 -779 1089 -747
rect 1259 -749 1417 -747
rect 1316 -750 1350 -749
rect 556 -840 656 -824
rect 556 -902 688 -840
rect 890 -844 950 -779
rect 1528 -799 1562 -576
rect 1016 -852 1022 -850
rect 984 -888 1022 -852
rect 556 -924 656 -902
rect 771 -935 911 -901
rect 1016 -902 1022 -888
rect 1074 -902 1080 -850
rect 1116 -860 1172 -800
rect 1495 -859 1562 -799
rect 825 -1049 859 -935
rect 1116 -1049 1150 -860
rect 1580 -1034 1680 -982
rect 1580 -1049 1610 -1034
rect 825 -1069 1610 -1049
rect 1645 -1069 1680 -1034
rect 825 -1082 1680 -1069
rect 825 -1083 1597 -1082
<< via1 >>
rect 582 110 634 162
rect 864 -198 916 -146
rect 771 -442 823 -390
rect 1022 -902 1074 -850
<< metal2 >>
rect 582 162 634 168
rect 561 110 582 133
rect 561 104 634 110
rect 561 99 625 104
rect 561 -225 595 99
rect 864 -146 916 -140
rect 864 -204 916 -198
rect 561 -259 814 -225
rect 780 -384 814 -259
rect 873 -243 907 -204
rect 873 -277 1087 -243
rect 771 -390 823 -384
rect 1053 -389 1087 -277
rect 1053 -423 1174 -389
rect 771 -448 823 -442
rect 1140 -643 1174 -423
rect 1069 -677 1174 -643
rect 1069 -753 1103 -677
rect 1031 -787 1103 -753
rect 1031 -844 1065 -787
rect 1022 -850 1074 -844
rect 1022 -908 1074 -902
use sky130_fd_pr__nfet_01v8_X33H33  XM0
timestamp 1706216322
transform 0 -1 836 1 0 -871
box -211 -320 211 320
use sky130_fd_pr__pfet_01v8_AMA9E4  XM1
timestamp 1706216322
transform 1 0 892 0 1 -25
box -332 -263 332 263
use sky130_fd_pr__nfet_01v8_LH5FDA  XM2
timestamp 1706211875
transform -1 0 862 0 1 -558
box -260 -252 346 252
use sky130_fd_pr__pfet_01v8_8DZSNJ  XM3
timestamp 1706216322
transform 1 0 1406 0 1 -155
box -212 -319 212 319
use sky130_fd_pr__nfet_01v8_LH5FDA  XM4
timestamp 1706211875
transform 1 0 1334 0 1 -830
box -260 -252 346 252
<< labels >>
flabel metal1 1580 -1082 1680 -982 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 1530 -576 1630 -476 0 FreeSans 256 0 0 0 V03
port 1 nsew
flabel metal1 1196 104 1296 204 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 556 -924 656 -824 0 FreeSans 256 0 0 0 Vin
port 2 nsew
<< end >>
