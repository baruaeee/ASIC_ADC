magic
tech sky130A
magscale 1 2
timestamp 1706224144
<< error_p >>
rect -325 159 -308 265
rect -289 195 -272 229
<< nwell >>
rect -308 -269 308 269
<< pmos >>
rect -112 -50 112 50
<< pdiff >>
rect -170 38 -112 50
rect -170 -38 -158 38
rect -124 -38 -112 38
rect -170 -50 -112 -38
rect 112 38 170 50
rect 112 -38 124 38
rect 158 -38 170 38
rect 112 -50 170 -38
<< pdiffc >>
rect -158 -38 -124 38
rect 124 -38 158 38
<< nsubdiff >>
rect -289 195 -176 229
rect 176 195 238 229
<< nsubdiffcont >>
rect -176 195 176 229
<< poly >>
rect -112 131 112 147
rect -112 97 -96 131
rect 96 97 112 131
rect -112 50 112 97
rect -112 -97 112 -50
rect -112 -131 -96 -97
rect 96 -131 112 -97
rect -112 -147 112 -131
<< polycont >>
rect -96 97 96 131
rect -96 -131 96 -97
<< locali >>
rect -283 195 -176 229
rect 176 195 238 229
rect -112 97 -96 131
rect 96 97 112 131
rect -158 38 -124 54
rect -158 -54 -124 -38
rect 124 38 158 54
rect 124 -54 158 -38
rect -112 -131 -96 -97
rect 96 -131 112 -97
<< viali >>
rect -96 97 96 131
rect -158 -38 -124 38
rect 124 -38 158 38
rect -96 -131 96 -97
<< metal1 >>
rect -108 131 108 137
rect -108 97 -96 131
rect 96 97 108 131
rect -108 91 108 97
rect -164 38 -118 50
rect -164 -38 -158 38
rect -124 -38 -118 38
rect -164 -50 -118 -38
rect 118 38 164 50
rect 118 -38 124 38
rect 158 -38 164 38
rect 118 -50 164 -38
rect -108 -97 108 -91
rect -108 -131 -96 -97
rect 96 -131 108 -97
rect -108 -137 108 -131
<< properties >>
string FIXED_BBOX -255 -216 255 216
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 1.12 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
