magic
tech sky130A
magscale 1 2
timestamp 1704371799
<< locali >>
rect 826 -144 970 -38
rect 880 -1464 964 -1316
<< metal1 >>
rect 894 255 1094 398
rect 753 221 1321 255
rect 753 -65 787 221
rect 894 198 1094 221
rect 1287 179 1321 221
rect 1287 145 1387 179
rect 1287 129 1351 145
rect 1353 129 1387 145
rect 1287 95 1387 129
rect 1729 119 1820 159
rect 1287 91 1347 95
rect 1725 85 1820 119
rect 968 8 1026 68
rect 1115 11 1467 45
rect 1785 20 1820 85
rect 753 -175 788 -65
rect 753 -209 971 -175
rect 1115 -245 1149 11
rect 1025 -247 1149 -245
rect 1025 -281 1487 -247
rect 1025 -343 1114 -281
rect 1785 -319 1819 20
rect 754 -425 1033 -391
rect 754 -580 788 -425
rect 670 -780 870 -580
rect 754 -985 788 -780
rect 1080 -849 1114 -343
rect 1286 -377 1389 -331
rect 1731 -357 1819 -319
rect 1283 -391 1389 -377
rect 1283 -411 1381 -391
rect 1283 -741 1320 -411
rect 1727 -415 1819 -357
rect 1718 -741 1918 -648
rect 1283 -775 1918 -741
rect 1283 -829 1323 -775
rect 925 -883 1205 -849
rect 1283 -863 1449 -829
rect 1718 -848 1918 -775
rect 925 -943 959 -883
rect 891 -977 959 -943
rect 754 -1039 837 -985
rect 1171 -1071 1205 -883
rect 1415 -1049 1449 -863
rect 1313 -1071 1347 -1051
rect 1171 -1105 1347 -1071
rect 886 -1317 958 -1310
rect 886 -1360 973 -1317
rect 1196 -1360 1396 -1292
rect 1455 -1360 1509 -1103
rect 1730 -1112 1782 -1046
rect 886 -1412 1509 -1360
rect 889 -1414 1509 -1412
rect 1196 -1492 1396 -1414
use sky130_fd_pr__nfet_01v8_JLSX9N  XM0
timestamp 1704371799
transform 0 -1 922 1 0 -1145
box -353 -252 353 252
use sky130_fd_pr__pfet_01v8_XYZSMQ  XM1
timestamp 1704371799
transform -1 0 999 0 -1 -185
box -211 -377 211 377
use sky130_fd_pr__pfet_01v8_AZD9DW  XM2
timestamp 1704371799
transform 1 0 1557 0 1 137
box -353 -261 353 261
use sky130_fd_pr__pfet_01v8_AZD9DW  XM3
timestamp 1704371799
transform 1 0 1561 0 1 -373
box -353 -261 353 261
use sky130_fd_pr__nfet_01v8_T8HSQ7  XM4
timestamp 1704371799
transform 0 -1 1541 1 0 -1077
box -211 -367 211 367
<< labels >>
flabel metal1 1718 -848 1918 -648 0 FreeSans 256 0 0 0 V09
port 1 nsew
flabel metal1 1196 -1492 1396 -1292 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 670 -780 870 -580 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 894 198 1094 398 0 FreeSans 256 0 0 0 Vp
port 0 nsew
<< end >>
