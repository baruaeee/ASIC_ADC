magic
tech sky130A
magscale 1 2
timestamp 1705015045
<< error_s >>
rect 590 765 631 797
rect 996 717 1037 749
rect 1494 669 1535 701
rect 1808 621 1849 653
rect 2306 573 2347 605
rect 2620 525 2657 557
rect 2934 477 2975 509
rect 3248 429 3289 461
rect 3746 381 3787 413
rect 4558 285 4599 317
rect 4964 237 5005 269
rect 5278 189 5315 221
rect 5684 141 5713 173
rect 6274 93 6315 125
rect 6588 45 6625 77
rect 7086 -3 7127 29
rect 8082 -99 8123 -67
rect 9668 -243 9697 -211
rect 10166 -291 10207 -259
rect 11254 -387 11295 -355
rect 11844 -435 11885 -403
rect 13798 -579 13837 -547
rect 14702 -675 14743 -643
rect 15108 -723 15137 -691
rect 15422 -771 15463 -739
rect 15920 -819 15961 -787
rect 16640 -915 16677 -883
rect 17636 -1011 17649 -979
rect 238 -7387 279 -7355
rect 644 -7435 685 -7403
rect 1142 -7483 1183 -7451
rect 1456 -7531 1497 -7499
rect 1954 -7579 1995 -7547
rect 2268 -7627 2305 -7595
rect 2582 -7675 2623 -7643
rect 2896 -7723 2937 -7691
rect 3394 -7771 3435 -7739
rect 4206 -7867 4247 -7835
rect 4612 -7915 4653 -7883
rect 4926 -7963 4963 -7931
rect 5332 -8011 5361 -7979
rect 5922 -8059 5963 -8027
rect 6236 -8107 6273 -8075
rect 6734 -8155 6775 -8123
rect 7730 -8251 7771 -8219
rect 9316 -8395 9345 -8363
rect 9814 -8443 9855 -8411
rect 10902 -8539 10943 -8507
rect 11492 -8587 11533 -8555
rect 13446 -8731 13485 -8699
rect 14350 -8827 14391 -8795
rect 14756 -8875 14785 -8843
rect 15070 -8923 15111 -8891
rect 15568 -8971 15609 -8939
rect 16288 -9067 16325 -9035
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
use sky130_fd_sc_hd__a22oi_1  sky130_fd_sc_hd__a22oi_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 5370 0 1 -8272
box -38 -48 590 592
use sky130_fd_sc_hd__a32oi_1  sky130_fd_sc_hd__a32oi_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 12120 0 1 -8896
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  sky130_fd_sc_hd__a211oi_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 11530 0 1 -8848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3432 0 1 -8032
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  sky130_fd_sc_hd__lpflow_inputiso1p_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 6772 0 1 -8416
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 -38 0 1 -7600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1696625445
transform 1 0 1180 0 1 -7744
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_2
timestamp 1696625445
transform 1 0 2306 0 1 -7888
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_3
timestamp 1696625445
transform 1 0 2620 0 1 -7936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_4
timestamp 1696625445
transform 1 0 3930 0 1 -8080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_5
timestamp 1696625445
transform 1 0 14074 0 1 -9040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_6
timestamp 1696625445
transform 1 0 14794 0 1 -9136
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_7
timestamp 1696625445
transform 1 0 15284 0 1 -6676
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  sky130_fd_sc_hd__nand2b_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 7768 0 1 -8512
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 276 0 1 -7648
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_1
timestamp 1696625445
transform 1 0 4244 0 1 -8128
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  sky130_fd_sc_hd__nand3b_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 13484 0 1 -8992
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  sky130_fd_sc_hd__nand4_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 682 0 1 -7696
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  sky130_fd_sc_hd__nand4_1_1
timestamp 1696625445
transform 1 0 1494 0 1 -7792
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  sky130_fd_sc_hd__nand4_1_2
timestamp 1696625445
transform 1 0 15108 0 1 -9184
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 1992 0 1 -7840
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1696625445
transform 1 0 4650 0 1 -8176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_2
timestamp 1696625445
transform 1 0 5960 0 1 -8320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_3
timestamp 1696625445
transform 1 0 16012 0 1 -9280
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  sky130_fd_sc_hd__nor3_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 4964 0 1 -8224
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  sky130_fd_sc_hd__nor3_1_1
timestamp 1696625445
transform 1 0 8948 0 1 -8608
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  sky130_fd_sc_hd__nor3_1_2
timestamp 1696625445
transform 1 0 14388 0 1 -9088
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  sky130_fd_sc_hd__nor4_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 2934 0 1 -7984
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  sky130_fd_sc_hd__nor4_1_1
timestamp 1696625445
transform 1 0 7270 0 1 -8464
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  sky130_fd_sc_hd__nor4_1_2
timestamp 1696625445
transform 1 0 9354 0 1 -8656
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  sky130_fd_sc_hd__nor4b_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 8266 0 1 -8560
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_0  sky130_fd_sc_hd__o21ai_0_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 9852 0 1 -8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_0  sky130_fd_sc_hd__o21ai_0_1
timestamp 1696625445
transform 1 0 15606 0 1 -9232
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_0  sky130_fd_sc_hd__o21ai_0_2
timestamp 1696625445
transform 1 0 16326 0 1 -9328
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  sky130_fd_sc_hd__o31ai_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 16732 0 1 -9376
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  sky130_fd_sc_hd__o2111ai_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 12802 0 1 -8944
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  sky130_fd_sc_hd__or3_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 6274 0 1 -8368
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  sky130_fd_sc_hd__or3b_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 10258 0 1 -8752
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  sky130_fd_sc_hd__or4_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 10940 0 1 -8800
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_1  x0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 0 0 1 600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x1
timestamp 1696625445
transform 1 0 314 0 1 552
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  x2
timestamp 1696625445
transform 1 0 628 0 1 504
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  x3
timestamp 1696625445
transform 1 0 1034 0 1 456
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  x4
timestamp 1696625445
transform 1 0 1532 0 1 408
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  x5
timestamp 1696625445
transform 1 0 1846 0 1 360
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  x6
timestamp 1696625445
transform 1 0 2344 0 1 312
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x7
timestamp 1696625445
transform 1 0 2658 0 1 264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x8
timestamp 1696625445
transform 1 0 2972 0 1 216
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  x9
timestamp 1696625445
transform 1 0 3286 0 1 168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x10
timestamp 1696625445
transform 1 0 3784 0 1 120
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  x11
timestamp 1696625445
transform 1 0 4282 0 1 72
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  x12
timestamp 1696625445
transform 1 0 4596 0 1 24
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  x13
timestamp 1696625445
transform 1 0 5002 0 1 -24
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  x14
timestamp 1696625445
transform 1 0 5316 0 1 -72
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  x15
timestamp 1696625445
transform 1 0 5722 0 1 -120
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  x16
timestamp 1696625445
transform 1 0 6312 0 1 -168
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  x17
timestamp 1696625445
transform 1 0 6626 0 1 -216
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  x18
timestamp 1696625445
transform 1 0 7124 0 1 -264
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  x19
timestamp 1696625445
transform 1 0 7622 0 1 -312
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  x20
timestamp 1696625445
transform 1 0 8120 0 1 -360
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  x21
timestamp 1696625445
transform 1 0 8618 0 1 -408
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  x22
timestamp 1696625445
transform 1 0 9300 0 1 -456
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  x23
timestamp 1696625445
transform 1 0 9706 0 1 -504
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_0  x24
timestamp 1696625445
transform 1 0 10204 0 1 -552
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  x25
timestamp 1696625445
transform 1 0 10610 0 1 -600
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  x26
timestamp 1696625445
transform 1 0 11292 0 1 -648
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  x27
timestamp 1696625445
transform 1 0 11882 0 1 -696
box -38 -48 590 592
use sky130_fd_sc_hd__a32oi_1  x28
timestamp 1696625445
transform 1 0 12472 0 1 -744
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  x29
timestamp 1696625445
transform 1 0 13154 0 1 -792
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  x30
timestamp 1696625445
transform 1 0 13836 0 1 -840
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  x31
timestamp 1696625445
transform 1 0 14426 0 1 -888
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  x32
timestamp 1696625445
transform 1 0 14740 0 1 -936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  x33
timestamp 1696625445
transform 1 0 15146 0 1 -984
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  x34
timestamp 1696625445
transform 1 0 15460 0 1 -1032
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_0  x35
timestamp 1696625445
transform 1 0 15958 0 1 -1080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  x36
timestamp 1696625445
transform 1 0 16364 0 1 -1128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_0  x37
timestamp 1696625445
transform 1 0 16678 0 1 -1176
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  x38
timestamp 1696625445
transform 1 0 17084 0 1 -1224
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  x39
timestamp 1696625445
transform 1 0 17674 0 1 -1272
box -38 -48 314 592
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {p\[0\]}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 {p\[1\]}
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 {p\[2\]}
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 {b\[0\]}
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 {p\[3\]}
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 {p\[4\]}
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 {b\[1\]}
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 {p\[5\]}
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 {p\[6\]}
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 {p\[7\]}
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 {b\[2\]}
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 {p\[8\]}
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 {p\[9\]}
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 {b\[3\]}
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 {p\[10\]}
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 {p\[11\]}
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 {}
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 {p\[12\]}
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 {p\[13\]}
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 {p\[14\]}
port 19 nsew
<< end >>
