** sch_path: /home/exotic/Desktop/ASIC_ADC/xschem/Vth_sch/Pre_layout/th01_1.sch
**.subckt th01_1 Vin Vout Vin
*.ipin Vin
*.opin Vout
*.ipin Vin
VDD VDD GND 1.8
Vin Vin GND pulse(0 0.2 0ns 1ns 1ns 5ns 10ns)
V_logic_high V_LH GND 1.25
V_logic_low V_LL GND 0.5
x1 VDD net1 Vout GND th01
x2 VDD Vin net1 GND preamp
C0 Vp net1 0.173f
C1 net1 Vin 0.0029f
C2 Vout Vin 8.58e-20
C3 net1 Vp 0.156f
C4 net1 Vn 0.00347f
C5 Vp Vout 1.44e-19
C6 net1 Vin 0.00888f
C7 net1 0 2.24f
C8 Vin 0 2.67f
C9 Vp 0 3.38f
C10 Vout 0 0.247f
C11 net1 0 0.96f
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.save all





.dc Vin 0 1.8 0.01
*.tran 1n 30n
.control
run
set color0=white
set color1=black
plot Vin Vout V_LH V_LL
set xbrushwidth=3
.save all
.endc
.end


**** end user architecture code
**.ends

* NGSPICE file created from th01.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_9DPZTU w_n291_n261# a_n153_n42# a_n95_n139# a_95_n42#
+ VSUBS
X0 a_95_n42# a_n95_n139# a_n153_n42# w_n291_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.95
C0 w_n291_n261# a_n153_n42# 0.0499f
C1 a_n95_n139# a_n153_n42# 0.014f
C2 a_n95_n139# w_n291_n261# 0.419f
C3 a_n153_n42# a_95_n42# 0.0249f
C4 w_n291_n261# a_95_n42# 0.0499f
C5 a_n95_n139# a_95_n42# 0.014f
C6 a_95_n42# VSUBS 0.0313f
C7 a_n153_n42# VSUBS 0.0313f
C8 a_n95_n139# VSUBS 0.289f
C9 w_n291_n261# VSUBS 1.36f
.ends

.subckt sky130_fd_pr__nfet_01v8_586EUA a_n97_n95# a_n199_n269# a_n39_n183# a_39_n95#
X0 a_39_n95# a_n39_n183# a_n97_n95# a_n199_n269# sky130_fd_pr__nfet_01v8 ad=0.275 pd=2.48 as=0.275 ps=2.48 w=0.95 l=0.39
C0 a_n39_n183# a_39_n95# 0.0127f
C1 a_n97_n95# a_39_n95# 0.1f
C2 a_n97_n95# a_n39_n183# 0.0127f
C3 a_39_n95# a_n199_n269# 0.135f
C4 a_n97_n95# a_n199_n269# 0.135f
C5 a_n39_n183# a_n199_n269# 0.381f
.ends

.subckt sky130_fd_pr__nfet_01v8_PJBF84 a_n248_n222# a_n146_n48# a_88_n48# a_n88_n136#
X0 a_88_n48# a_n88_n136# a_n146_n48# a_n248_n222# sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.54 as=0.139 ps=1.54 w=0.48 l=0.88
C0 a_n88_n136# a_88_n48# 0.0146f
C1 a_n146_n48# a_88_n48# 0.03f
C2 a_n146_n48# a_n88_n136# 0.0146f
C3 a_88_n48# a_n248_n222# 0.088f
C4 a_n146_n48# a_n248_n222# 0.088f
C5 a_n88_n136# a_n248_n222# 0.649f
.ends

.subckt sky130_fd_pr__pfet_01v8_RVEGTV a_n69_n175# a_n127_n78# w_n265_n297# a_69_n78#
+ VSUBS
X0 a_69_n78# a_n69_n175# a_n127_n78# w_n265_n297# sky130_fd_pr__pfet_01v8 ad=0.226 pd=2.14 as=0.226 ps=2.14 w=0.78 l=0.69
C0 w_n265_n297# a_n127_n78# 0.0718f
C1 a_n69_n175# a_n127_n78# 0.0173f
C2 a_n69_n175# w_n265_n297# 0.338f
C3 a_n127_n78# a_69_n78# 0.0574f
C4 w_n265_n297# a_69_n78# 0.0718f
C5 a_n69_n175# a_69_n78# 0.0173f
C6 a_69_n78# VSUBS 0.0474f
C7 a_n127_n78# VSUBS 0.0474f
C8 a_n69_n175# VSUBS 0.227f
C9 w_n265_n297# VSUBS 1.41f
.ends

.subckt th01 Vp Vin Vout Vn
XXM2 Vp Vp Vin m1_732_n84# Vn sky130_fd_pr__pfet_01v8_9DPZTU
XXM3 Vn Vn Vin m1_732_n84# sky130_fd_pr__nfet_01v8_586EUA
XXM4 Vn Vn Vout m1_732_n84# sky130_fd_pr__nfet_01v8_PJBF84
XXM5 m1_732_n84# Vp Vp Vout Vn sky130_fd_pr__pfet_01v8_RVEGTV
C0 Vn Vp 0.167f
C1 Vn Vin 0.0827f
C2 Vn m1_732_n84# 0.18f
C3 Vout Vp 0.0895f
C4 Vout Vin 1.54e-19
C5 Vout m1_732_n84# 0.174f
C6 Vin Vp 0.228f
C7 Vn Vout 0.0643f
C8 m1_732_n84# Vp 0.305f
C9 m1_732_n84# Vin 0.174f
C10 Vin 0 0.683f
C11 Vp 0 2.57f
C12 Vout 0 0.247f
C13 m1_732_n84# 0 0.96f
C14 Vn 0 0.0948f
.ends



* NGSPICE file created from preamp.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_4N47A3 w_n231_n369# a_n93_n150# a_35_n150# a_n35_n247#
+ VSUBS
X0 a_35_n150# a_n35_n247# a_n93_n150# w_n231_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.35
C0 a_35_n150# a_n35_n247# 0.0165f
C1 a_n93_n150# a_n35_n247# 0.0165f
C2 a_n93_n150# a_35_n150# 0.166f
C3 a_n35_n247# w_n231_n369# 0.233f
C4 a_35_n150# w_n231_n369# 0.116f
C5 a_n93_n150# w_n231_n369# 0.116f
C6 a_35_n150# VSUBS 0.0757f
C7 a_n93_n150# VSUBS 0.0757f
C8 a_n35_n247# VSUBS 0.141f
C9 w_n231_n369# VSUBS 1.52f
.ends

.subckt sky130_fd_pr__nfet_01v8_48YMBA a_n518_n42# a_460_n42# a_n620_n216# a_n460_n130#
X0 a_460_n42# a_n460_n130# a_n518_n42# a_n620_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=4.6
C0 a_460_n42# a_n518_n42# 0.00624f
C1 a_n518_n42# a_n460_n130# 0.0236f
C2 a_460_n42# a_n460_n130# 0.0236f
C3 a_460_n42# a_n620_n216# 0.0868f
C4 a_n518_n42# a_n620_n216# 0.0868f
C5 a_n460_n130# a_n620_n216# 2.69f
.ends

.subckt preamp Vp Vin Vpamp Vn
XXM0 Vpamp Vn Vpamp Vin Vpamp sky130_fd_pr__pfet_01v8_4N47A3
XXM1 Vp Vpamp Vpamp Vin sky130_fd_pr__nfet_01v8_48YMBA
C0 Vn Vpamp 0.213f
C1 Vpamp Vp 0.0775f
C2 Vin Vpamp 0.488f
C3 Vn Vp 0.0228f
C4 Vin Vn 0.0147f
C5 Vin Vp 0.233f
C6 Vpamp 0 1.57f
C7 Vp 0 0.377f
C8 Vin 0 2.67f
C9 Vn 0 0.247f
.ends


.GLOBAL VDD
.GLOBAL GND
.GLOBAL V_LH
.GLOBAL V_LL
.end
