/home/cae3/Desktop/ADC/ASIC_ADC/PNR/lef/pre_therm_MACRO.lef