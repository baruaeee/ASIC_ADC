magic
tech sky130A
magscale 1 2
timestamp 1704730646
<< pwell >>
rect -201 -1798 201 1798
<< psubdiff >>
rect -165 1728 -69 1762
rect 69 1728 165 1762
rect -165 1666 -131 1728
rect 131 1666 165 1728
rect -165 -1728 -131 -1666
rect 131 -1728 165 -1666
rect -165 -1762 -69 -1728
rect 69 -1762 165 -1728
<< psubdiffcont >>
rect -69 1728 69 1762
rect -165 -1666 -131 1666
rect 131 -1666 165 1666
rect -69 -1762 69 -1728
<< xpolycontact >>
rect -35 1200 35 1632
rect -35 -1632 35 -1200
<< xpolyres >>
rect -35 -1200 35 1200
<< locali >>
rect -165 1728 -69 1762
rect 69 1728 165 1762
rect -165 1666 -131 1728
rect 131 1666 165 1728
rect -165 -1728 -131 -1666
rect 131 -1728 165 -1666
rect -165 -1762 -69 -1728
rect 69 -1762 165 -1728
<< viali >>
rect -19 1217 19 1614
rect -19 -1614 19 -1217
<< metal1 >>
rect -25 1614 25 1626
rect -25 1217 -19 1614
rect 19 1217 25 1614
rect -25 1205 25 1217
rect -25 -1217 25 -1205
rect -25 -1614 -19 -1217
rect 19 -1614 25 -1217
rect -25 -1626 25 -1614
<< properties >>
string FIXED_BBOX -148 -1745 148 1745
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 12.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 69.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
