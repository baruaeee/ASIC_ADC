magic
tech sky130A
timestamp 1706134018
<< pwell >>
rect -273 -155 273 155
<< nmos >>
rect -175 -50 175 50
<< ndiff >>
rect -204 44 -175 50
rect -204 -44 -198 44
rect -181 -44 -175 44
rect -204 -50 -175 -44
rect 175 44 204 50
rect 175 -44 181 44
rect 198 -44 204 44
rect 175 -50 204 -44
<< ndiffc >>
rect -198 -44 -181 44
rect 181 -44 198 44
<< psubdiff >>
rect -255 120 -207 137
rect 207 120 255 137
rect -255 89 -238 120
rect 238 89 255 120
rect -255 -120 -238 -89
rect 238 -120 255 -89
rect -255 -137 -207 -120
rect 207 -137 255 -120
<< psubdiffcont >>
rect -207 120 207 137
rect -255 -89 -238 89
rect 238 -89 255 89
rect -207 -137 207 -120
<< poly >>
rect -175 86 175 94
rect -175 69 -167 86
rect 167 69 175 86
rect -175 50 175 69
rect -175 -69 175 -50
rect -175 -86 -167 -69
rect 167 -86 175 -69
rect -175 -94 175 -86
<< polycont >>
rect -167 69 167 86
rect -167 -86 167 -69
<< locali >>
rect -255 120 -207 137
rect 207 120 255 137
rect -255 89 -238 120
rect 238 89 255 120
rect -175 69 -167 86
rect 167 69 175 86
rect -198 44 -181 52
rect -198 -52 -181 -44
rect 181 44 198 52
rect 181 -52 198 -44
rect -175 -86 -167 -69
rect 167 -86 175 -69
rect -255 -120 -238 -89
rect 238 -120 255 -89
rect -255 -137 -207 -120
rect 207 -137 255 -120
<< viali >>
rect -167 69 167 86
rect -198 -44 -181 44
rect 181 -44 198 44
rect -167 -86 167 -69
<< metal1 >>
rect -173 86 173 89
rect -173 69 -167 86
rect 167 69 173 86
rect -173 66 173 69
rect -201 44 -178 50
rect -201 -44 -198 44
rect -181 -44 -178 44
rect -201 -50 -178 -44
rect 178 44 201 50
rect 178 -44 181 44
rect 198 -44 201 44
rect 178 -50 201 -44
rect -173 -69 173 -66
rect -173 -86 -167 -69
rect 167 -86 173 -69
rect -173 -89 173 -86
<< properties >>
string FIXED_BBOX -246 -128 246 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 3.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
