* NGSPICE file created from th13.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n73_n100# w_n211_n319# 0.0813f
C1 a_n33_n197# w_n211_n319# 0.246f
C2 a_n33_n197# a_n73_n100# 0.0281f
C3 a_15_n100# w_n211_n319# 0.0815f
C4 a_15_n100# a_n73_n100# 0.162f
C5 a_15_n100# a_n33_n197# 0.0262f
C6 a_15_n100# VSUBS 0.0492f
C7 a_n73_n100# VSUBS 0.0487f
C8 a_n33_n197# VSUBS 0.129f
C9 w_n211_n319# VSUBS 1.23f
.ends

.subckt sky130_fd_pr__nfet_01v8_L6G859 a_n288_n42# a_230_n42# a_n390_n216# a_n230_n130#
X0 a_230_n42# a_n230_n130# a_n288_n42# a_n390_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.3
C0 a_230_n42# a_n230_n130# 0.0204f
C1 a_n288_n42# a_n230_n130# 0.0204f
C2 a_n288_n42# a_230_n42# 0.0119f
C3 a_230_n42# a_n390_n216# 0.0846f
C4 a_n288_n42# a_n390_n216# 0.0846f
C5 a_n230_n130# a_n390_n216# 1.43f
.ends

.subckt sky130_fd_pr__pfet_01v8_XW9KDL a_n73_n230# a_n33_n327# a_15_n230# w_n211_n449#
+ VSUBS
X0 a_15_n230# a_n33_n327# a_n73_n230# w_n211_n449# sky130_fd_pr__pfet_01v8 ad=0.667 pd=5.18 as=0.667 ps=5.18 w=2.3 l=0.15
C0 a_n73_n230# w_n211_n449# 0.161f
C1 a_n33_n327# w_n211_n449# 0.246f
C2 a_n33_n327# a_n73_n230# 0.0338f
C3 a_15_n230# w_n211_n449# 0.161f
C4 a_15_n230# a_n73_n230# 0.369f
C5 a_15_n230# a_n33_n327# 0.0338f
C6 a_15_n230# VSUBS 0.102f
C7 a_n73_n230# VSUBS 0.102f
C8 a_n33_n327# VSUBS 0.129f
C9 w_n211_n449# VSUBS 1.69f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GC6 a_200_n42# w_n396_n261# a_n200_n139# a_n258_n42#
+ VSUBS
X0 a_200_n42# a_n200_n139# a_n258_n42# w_n396_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_n258_n42# w_n396_n261# 0.0498f
C1 a_n200_n139# w_n396_n261# 0.743f
C2 a_n200_n139# a_n258_n42# 0.0196f
C3 a_200_n42# w_n396_n261# 0.0498f
C4 a_200_n42# a_n258_n42# 0.0134f
C5 a_200_n42# a_n200_n139# 0.0196f
C6 a_200_n42# VSUBS 0.0338f
C7 a_n258_n42# VSUBS 0.0338f
C8 a_n200_n139# VSUBS 0.554f
C9 w_n396_n261# VSUBS 1.79f
.ends

.subckt sky130_fd_pr__nfet_01v8_ATLS57 a_15_n200# a_n175_n374# a_n73_n200# a_n33_n288#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n175_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_15_n200# a_n33_n288# 0.0357f
C1 a_n73_n200# a_n33_n288# 0.0336f
C2 a_n73_n200# a_15_n200# 0.321f
C3 a_15_n200# a_n175_n374# 0.232f
C4 a_n73_n200# a_n175_n374# 0.232f
C5 a_n33_n288# a_n175_n374# 0.358f
.ends

.subckt th13 Vp Vout Vin Vn
XXM0 m1_724_n958# Vn Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 m1_546_n454# m1_724_n958# Vn Vin sky130_fd_pr__nfet_01v8_L6G859
XXM2 m1_546_n454# Vin Vp Vp Vn sky130_fd_pr__pfet_01v8_XW9KDL
XXM3 Vout Vp m1_546_n454# Vp Vn sky130_fd_pr__pfet_01v8_VZ9GC6
XXM4 Vout Vn Vn m1_546_n454# sky130_fd_pr__nfet_01v8_ATLS57
C0 Vn Vout 0.147f
C1 Vin Vp 0.151f
C2 Vp m1_724_n958# 0.312f
C3 Vin Vout 0.00172f
C4 m1_546_n454# Vp 0.574f
C5 Vout m1_724_n958# 0.00247f
C6 m1_546_n454# Vout 0.546f
C7 Vin Vn 0.126f
C8 Vp Vout 0.346f
C9 Vn m1_724_n958# 0.0967f
C10 m1_546_n454# Vn 0.331f
C11 Vin m1_724_n958# 0.14f
C12 Vin m1_546_n454# 0.349f
C13 m1_546_n454# m1_724_n958# 0.0214f
C14 Vp Vn 0.589f
C15 Vn 0 0.573f
C16 Vout 0 0.513f
C17 Vp 0 4.74f
C18 m1_546_n454# 0 1.54f
C19 Vin 0 1.66f
C20 m1_724_n958# 0 0.188f
.ends

