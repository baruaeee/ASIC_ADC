magic
tech sky130A
magscale 1 2
timestamp 1704387829
<< pwell >>
rect 528 -874 598 -705
<< locali >>
rect 342 -244 492 -156
rect 724 -422 1097 -357
rect 742 -812 1097 -726
rect 524 -1089 594 -920
<< metal1 >>
rect 342 -26 1146 62
rect 342 -156 430 -26
rect 800 -138 1000 -26
rect 342 -244 492 -156
rect 605 -225 715 -155
rect 608 -244 715 -225
rect 504 -287 594 -286
rect 504 -365 595 -287
rect 324 -431 595 -365
rect 645 -288 715 -244
rect 1058 -160 1146 -26
rect 1058 -248 1234 -160
rect 1342 -232 1528 -168
rect 645 -342 1332 -288
rect 324 -476 390 -431
rect 310 -676 510 -476
rect 324 -864 390 -676
rect 645 -705 715 -342
rect 528 -775 715 -705
rect 951 -659 1005 -342
rect 1464 -468 1528 -232
rect 1342 -604 1542 -468
rect 951 -713 1127 -659
rect 324 -930 484 -864
rect 528 -874 598 -775
rect 524 -1019 594 -926
rect 630 -932 700 -862
rect 1073 -875 1127 -713
rect 1252 -668 1542 -604
rect 1167 -875 1207 -859
rect 1252 -868 1316 -668
rect 822 -1019 1022 -906
rect 1073 -929 1207 -875
rect 1255 -1019 1325 -923
rect 1362 -928 1422 -864
rect 524 -1089 1325 -1019
rect 822 -1106 1022 -1089
use sky130_fd_pr__nfet_01v8_L7T3GD  XM0
timestamp 1704387395
transform 0 -1 560 1 0 -899
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_NZD9V2  XM1
timestamp 1704387395
transform 1 0 551 0 1 -199
box -243 -261 243 261
use sky130_fd_pr__pfet_01v8_3PDS9J  XM2
timestamp 1704387395
transform 1 0 1288 0 1 -201
box -240 -261 240 261
use sky130_fd_pr__nfet_01v8_97T34Z  XM3
timestamp 1704387395
transform 0 -1 1286 1 0 -895
box -211 -256 211 256
<< labels >>
flabel metal1 310 -676 510 -476 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 800 -138 1000 62 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 822 -1106 1022 -906 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 1342 -668 1542 -468 0 FreeSans 256 0 0 0 V06
port 2 nsew
<< end >>
