magic
tech sky130A
magscale 1 2
timestamp 1706233216
<< nwell >>
rect -244 -262 244 262
<< pmos >>
rect -48 -43 48 43
<< pdiff >>
rect -106 31 -48 43
rect -106 -31 -94 31
rect -60 -31 -48 31
rect -106 -43 -48 -31
rect 48 31 106 43
rect 48 -31 60 31
rect 94 -31 106 31
rect 48 -43 106 -31
<< pdiffc >>
rect -94 -31 -60 31
rect 60 -31 94 31
<< nsubdiff >>
rect -174 192 -112 226
rect 112 192 174 226
<< nsubdiffcont >>
rect -112 192 112 226
<< poly >>
rect -48 124 48 140
rect -48 90 -32 124
rect 32 90 48 124
rect -48 43 48 90
rect -48 -90 48 -43
rect -48 -124 -32 -90
rect 32 -124 48 -90
rect -48 -140 48 -124
<< polycont >>
rect -32 90 32 124
rect -32 -124 32 -90
<< locali >>
rect -174 192 -112 226
rect 112 192 174 226
rect -48 90 -32 124
rect 32 90 48 124
rect -94 31 -60 47
rect -94 -47 -60 -31
rect 60 31 94 47
rect 60 -47 94 -31
rect -48 -124 -32 -90
rect 32 -124 48 -90
<< viali >>
rect -32 90 32 124
rect -94 -31 -60 31
rect 60 -31 94 31
rect -32 -124 32 -90
<< metal1 >>
rect -44 124 44 130
rect -44 90 -32 124
rect 32 90 44 124
rect -44 84 44 90
rect -100 31 -54 43
rect -100 -31 -94 31
rect -60 -31 -54 31
rect -100 -43 -54 -31
rect 54 31 100 43
rect 54 -31 60 31
rect 94 -31 100 31
rect 54 -43 100 -31
rect -44 -90 44 -84
rect -44 -124 -32 -90
rect 32 -124 44 -90
rect -44 -130 44 -124
<< properties >>
string FIXED_BBOX -191 -209 191 209
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.43 l 0.48 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
