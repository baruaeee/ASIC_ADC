magic
tech sky130A
magscale 1 2
timestamp 1706458547
<< nwell >>
rect 532 -558 570 -68
<< pwell >>
rect 1472 -222 1506 -162
<< nsubdiff >>
rect 609 386 663 420
<< locali >>
rect 641 386 666 420
rect 1742 -711 1776 -693
<< viali >>
rect 607 386 641 420
rect 1040 -373 1074 -339
rect 1742 -745 1776 -711
<< metal1 >>
rect 536 432 636 454
rect 536 420 647 432
rect 536 386 607 420
rect 641 417 647 420
rect 641 386 1079 417
rect 536 383 1079 386
rect 536 374 647 383
rect 536 354 636 374
rect 1037 254 1079 383
rect 901 199 935 223
rect 1037 211 1098 254
rect 901 165 1005 199
rect 1064 194 1098 211
rect 1799 193 1867 255
rect 901 139 935 165
rect 971 135 1005 165
rect 971 101 1417 135
rect 778 20 784 72
rect 836 20 842 72
rect 800 -16 840 20
rect 753 -163 843 -161
rect 745 -167 843 -163
rect 737 -201 843 -167
rect 669 -325 727 -251
rect 807 -296 843 -201
rect 1132 -268 1166 101
rect 1833 -51 1867 193
rect 1472 -55 1947 -51
rect 1471 -89 1947 -55
rect 1471 -191 1507 -89
rect 1869 -94 1947 -89
rect 1869 -117 1980 -94
rect 1311 -225 1649 -191
rect 1880 -194 1980 -117
rect 1366 -281 1400 -276
rect 669 -534 703 -325
rect 807 -379 844 -296
rect 1225 -305 1673 -281
rect 1209 -315 1673 -305
rect 1037 -333 1087 -325
rect 1209 -333 1400 -315
rect 1034 -339 1400 -333
rect 1034 -373 1040 -339
rect 1074 -373 1400 -339
rect 1034 -379 1400 -373
rect 739 -413 1087 -379
rect 751 -417 1087 -413
rect 1037 -423 1087 -417
rect 1755 -449 1789 -229
rect 1660 -483 1789 -449
rect 1660 -531 1695 -483
rect 669 -568 1205 -534
rect 1171 -597 1205 -568
rect 1627 -595 1695 -531
rect 830 -667 930 -626
rect 830 -719 870 -667
rect 922 -719 930 -667
rect 1232 -667 1600 -646
rect 1232 -680 1360 -667
rect 830 -726 930 -719
rect 1412 -680 1600 -667
rect 1360 -725 1412 -719
rect 1706 -711 1806 -668
rect 1706 -745 1742 -711
rect 1776 -745 1806 -711
rect 1706 -768 1806 -745
<< via1 >>
rect 784 20 836 72
rect 870 -719 922 -667
rect 1360 -719 1412 -667
<< metal2 >>
rect 784 72 836 78
rect 836 20 840 46
rect 784 14 840 20
rect 793 -7 840 14
rect 793 -41 919 -7
rect 885 -667 919 -41
rect 864 -719 870 -667
rect 922 -676 928 -667
rect 1354 -676 1360 -667
rect 922 -710 1360 -676
rect 922 -719 928 -710
rect 1354 -719 1360 -710
rect 1412 -719 1418 -667
use sky130_fd_pr__pfet_01v8_LDQF7K  XM0
timestamp 1706457568
transform 1 0 769 0 1 -289
box -225 -269 225 269
use sky130_fd_pr__nfet_01v8_HZA4VB  XM1
timestamp 1706458450
transform 1 0 1416 0 1 -566
box -396 -206 396 252
use sky130_fd_pr__pfet_01v8_TM5S5A  XM2
timestamp 1706457568
transform 1 0 810 0 1 187
box -276 -269 276 269
use sky130_fd_pr__pfet_01v8_KQKFM4  XM3
timestamp 1706457568
transform 1 0 1458 0 1 223
box -526 -261 526 261
use sky130_fd_pr__nfet_01v8_KQFF5S  XM4
timestamp 1706458547
transform 0 -1 1464 1 0 -251
box -211 -460 155 444
<< labels >>
flabel metal1 536 354 636 454 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 1880 -194 1980 -94 0 FreeSans 256 0 0 0 V15
port 1 nsew
flabel metal1 830 -726 930 -626 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 1706 -768 1806 -668 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
