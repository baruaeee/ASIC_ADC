magic
tech sky130A
magscale 1 2
timestamp 1705440580
<< psubdiff >>
rect 1136 -1531 1170 -1292
<< locali >>
rect 1136 -923 1170 152
rect 3798 -208 3898 129
rect 2410 -1086 2562 -1082
rect 2410 -1096 2570 -1086
rect 2398 -1112 2570 -1096
rect 2410 -1116 2562 -1112
<< viali >>
rect 3798 129 3898 200
<< metal1 >>
rect 3870 606 4395 677
rect 3870 502 3941 606
rect 4146 502 4208 556
rect 3467 426 3542 446
rect 3744 426 3944 502
rect 3467 412 3944 426
rect 3469 401 3944 412
rect 1199 285 1283 377
rect 3495 375 3944 401
rect 3508 362 3944 375
rect 3519 355 3944 362
rect 1199 51 1241 285
rect 3744 200 3944 355
rect 4324 338 4395 606
rect 4203 267 4395 338
rect 3744 129 3798 200
rect 3898 129 3944 200
rect 3744 124 3944 129
rect 3786 123 3910 124
rect 1199 9 1534 51
rect 1114 -491 1314 -426
rect 1492 -444 1534 9
rect 3780 -434 3884 -366
rect 1114 -533 1671 -491
rect 1114 -626 1314 -533
rect 1232 -1082 1274 -626
rect 3816 -740 3884 -434
rect 1510 -774 3884 -740
rect 1510 -808 1514 -774
rect 1566 -808 3884 -774
rect 1514 -832 1566 -826
rect 1522 -1018 1558 -832
rect 2840 -1082 3040 -1076
rect 2301 -1116 3040 -1082
rect 1524 -1373 1560 -1176
rect 2840 -1265 3040 -1116
rect 2835 -1276 3040 -1265
rect 1514 -1379 1566 -1373
rect 2835 -1377 2883 -1276
rect 1514 -1437 1566 -1431
rect 1775 -1431 2883 -1377
rect 1775 -1475 1829 -1431
rect 1181 -1529 1829 -1475
rect 1181 -1661 1235 -1529
rect 3214 -1630 3282 -808
rect 3650 -1138 4148 -986
rect 3544 -1186 4148 -1138
rect 1181 -1753 1283 -1661
rect 3544 -1672 3592 -1186
rect 3508 -1750 3592 -1672
rect 3355 -1817 3513 -1789
rect 3355 -1844 3517 -1817
rect 4147 -1844 4201 -1779
rect 3355 -1898 4201 -1844
<< via1 >>
rect 1514 -826 1566 -774
rect 1514 -1431 1566 -1379
<< metal2 >>
rect 1508 -826 1514 -774
rect 1566 -783 1572 -774
rect 1566 -817 1649 -783
rect 1566 -826 1572 -817
rect 1508 -1431 1514 -1379
rect 1566 -1388 1572 -1379
rect 1615 -1388 1649 -817
rect 1566 -1422 1650 -1388
rect 1566 -1431 1572 -1422
use sky130_fd_pr__nfet_01v8_9GNSAK  XM0
timestamp 1704501535
transform 0 -1 1860 1 0 -1099
box -263 -760 263 760
use sky130_fd_pr__pfet_01v8_UTD9YE  XM1
timestamp 1704501257
transform 1 0 2682 0 1 -399
box -1296 -261 1296 261
use sky130_fd_pr__nfet_01v8_VZ7MP4  XM2
timestamp 1704501257
transform 1 0 2396 0 1 334
box -1296 -252 1296 252
use sky130_fd_pr__pfet_01v8_UGSTRG  XM3
timestamp 1704501257
transform 1 0 4178 0 1 -639
box -214 -1319 214 1319
use sky130_fd_pr__nfet_01v8_VZ7MP4  XM4
timestamp 1704501257
transform 1 0 2396 0 1 -1708
box -1296 -252 1296 252
<< labels >>
flabel metal1 1114 -626 1314 -426 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 3650 -1186 3850 -986 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 2840 -1276 3040 -1076 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 3744 302 3944 502 0 FreeSans 256 0 0 0 Vp
port 0 nsew
<< end >>
