magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< nwell >>
rect -488 -261 488 261
<< pmos >>
rect -292 -42 292 42
<< pdiff >>
rect -350 30 -292 42
rect -350 -30 -338 30
rect -304 -30 -292 30
rect -350 -42 -292 -30
rect 292 30 350 42
rect 292 -30 304 30
rect 338 -30 350 30
rect 292 -42 350 -30
<< pdiffc >>
rect -338 -30 -304 30
rect 304 -30 338 30
<< nsubdiff >>
rect -452 191 -356 225
rect 356 191 452 225
rect -452 129 -418 191
rect 418 129 452 191
rect -452 -191 -418 -129
rect 418 -191 452 -129
rect -452 -225 -356 -191
rect 356 -225 452 -191
<< nsubdiffcont >>
rect -356 191 356 225
rect -452 -129 -418 129
rect 418 -129 452 129
rect -356 -225 356 -191
<< poly >>
rect -292 123 292 139
rect -292 89 -276 123
rect 276 89 292 123
rect -292 42 292 89
rect -292 -89 292 -42
rect -292 -123 -276 -89
rect 276 -123 292 -89
rect -292 -139 292 -123
<< polycont >>
rect -276 89 276 123
rect -276 -123 276 -89
<< locali >>
rect -452 191 -356 225
rect 356 191 452 225
rect -452 129 -418 191
rect 418 129 452 191
rect -292 89 -276 123
rect 276 89 292 123
rect -338 30 -304 46
rect -338 -46 -304 -30
rect 304 30 338 46
rect 304 -46 338 -30
rect -292 -123 -276 -89
rect 276 -123 292 -89
rect -452 -191 -418 -129
rect 418 -191 452 -129
rect -452 -225 -356 -191
rect 356 -225 452 -191
<< viali >>
rect -276 89 276 123
rect -338 -30 -304 30
rect 304 -30 338 30
rect -276 -123 276 -89
<< metal1 >>
rect -288 123 288 129
rect -288 89 -276 123
rect 276 89 288 123
rect -288 83 288 89
rect -344 30 -298 42
rect -344 -30 -338 30
rect -304 -30 -298 30
rect -344 -42 -298 -30
rect 298 30 344 42
rect 298 -30 304 30
rect 338 -30 344 30
rect 298 -42 344 -30
rect -288 -89 288 -83
rect -288 -123 -276 -89
rect 276 -123 288 -89
rect -288 -129 288 -123
<< properties >>
string FIXED_BBOX -435 -208 435 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 2.92 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
