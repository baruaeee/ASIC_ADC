magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 114 29 120
rect -29 80 -17 114
rect -29 74 29 80
rect -29 -80 29 -74
rect -29 -114 -17 -80
rect -29 -120 29 -114
<< pwell >>
rect -212 -252 212 252
<< nmos >>
rect -16 -42 16 42
<< ndiff >>
rect -74 30 -16 42
rect -74 -30 -62 30
rect -28 -30 -16 30
rect -74 -42 -16 -30
rect 16 30 74 42
rect 16 -30 28 30
rect 62 -30 74 30
rect 16 -42 74 -30
<< ndiffc >>
rect -62 -30 -28 30
rect 28 -30 62 30
<< psubdiff >>
rect -176 182 -80 216
rect 80 182 176 216
rect -176 120 -142 182
rect 142 120 176 182
rect -176 -182 -142 -120
rect 142 -182 176 -120
rect -176 -216 -80 -182
rect 80 -216 176 -182
<< psubdiffcont >>
rect -80 182 80 216
rect -176 -120 -142 120
rect 142 -120 176 120
rect -80 -216 80 -182
<< poly >>
rect -33 114 33 130
rect -33 80 -17 114
rect 17 80 33 114
rect -33 64 33 80
rect -16 42 16 64
rect -16 -64 16 -42
rect -33 -80 33 -64
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -33 -130 33 -114
<< polycont >>
rect -17 80 17 114
rect -17 -114 17 -80
<< locali >>
rect -176 182 -80 216
rect 80 182 176 216
rect -176 120 -142 182
rect 142 120 176 182
rect -33 80 -17 114
rect 17 80 33 114
rect -62 30 -28 46
rect -62 -46 -28 -30
rect 28 30 62 46
rect 28 -46 62 -30
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -176 -182 -142 -120
rect 142 -182 176 -120
rect -176 -216 -80 -182
rect 80 -216 176 -182
<< viali >>
rect -17 80 17 114
rect -62 -30 -28 30
rect 28 -30 62 30
rect -17 -114 17 -80
<< metal1 >>
rect -29 114 29 120
rect -29 80 -17 114
rect 17 80 29 114
rect -29 74 29 80
rect -68 30 -22 42
rect -68 -30 -62 30
rect -28 -30 -22 30
rect -68 -42 -22 -30
rect 22 30 68 42
rect 22 -30 28 30
rect 62 -30 68 30
rect 22 -42 68 -30
rect -29 -80 29 -74
rect -29 -114 -17 -80
rect 17 -114 29 -80
rect -29 -120 29 -114
<< properties >>
string FIXED_BBOX -159 -199 159 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.155 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
