magic
tech sky130A
timestamp 1704310896
<< pwell >>
rect -213 -126 213 126
<< nmos >>
rect -115 -21 115 21
<< ndiff >>
rect -144 15 -115 21
rect -144 -15 -138 15
rect -121 -15 -115 15
rect -144 -21 -115 -15
rect 115 15 144 21
rect 115 -15 121 15
rect 138 -15 144 15
rect 115 -21 144 -15
<< ndiffc >>
rect -138 -15 -121 15
rect 121 -15 138 15
<< psubdiff >>
rect -195 91 -147 108
rect 147 91 195 108
rect -195 60 -178 91
rect 178 60 195 91
rect -195 -91 -178 -60
rect 178 -91 195 -60
rect -195 -108 -147 -91
rect 147 -108 195 -91
<< psubdiffcont >>
rect -147 91 147 108
rect -195 -60 -178 60
rect 178 -60 195 60
rect -147 -108 147 -91
<< poly >>
rect -115 57 115 65
rect -115 40 -107 57
rect 107 40 115 57
rect -115 21 115 40
rect -115 -40 115 -21
rect -115 -57 -107 -40
rect 107 -57 115 -40
rect -115 -65 115 -57
<< polycont >>
rect -107 40 107 57
rect -107 -57 107 -40
<< locali >>
rect -195 91 -147 108
rect 147 91 195 108
rect -195 60 -178 91
rect 178 60 195 91
rect -115 40 -107 57
rect 107 40 115 57
rect -138 15 -121 23
rect -138 -23 -121 -15
rect 121 15 138 23
rect 121 -23 138 -15
rect -115 -57 -107 -40
rect 107 -57 115 -40
rect -195 -91 -178 -60
rect 178 -91 195 -60
rect -195 -108 -147 -91
rect 147 -108 195 -91
<< viali >>
rect -107 40 107 57
rect -138 -15 -121 15
rect 121 -15 138 15
rect -107 -57 107 -40
<< metal1 >>
rect -113 57 113 60
rect -113 40 -107 57
rect 107 40 113 57
rect -113 37 113 40
rect -141 15 -118 21
rect -141 -15 -138 15
rect -121 -15 -118 15
rect -141 -21 -118 -15
rect 118 15 141 21
rect 118 -15 121 15
rect 138 -15 141 15
rect 118 -21 141 -15
rect -113 -40 113 -37
rect -113 -57 -107 -40
rect 107 -57 113 -40
rect -113 -60 113 -57
<< properties >>
string FIXED_BBOX -186 -99 186 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 2.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
