magic
tech sky130A
timestamp 1706204487
<< pwell >>
rect -273 -126 273 126
<< nmos >>
rect -175 -21 175 21
<< ndiff >>
rect -204 15 -175 21
rect -204 -15 -198 15
rect -181 -15 -175 15
rect -204 -21 -175 -15
rect 175 15 204 21
rect 175 -15 181 15
rect 198 -15 204 15
rect 175 -21 204 -15
<< ndiffc >>
rect -198 -15 -181 15
rect 181 -15 198 15
<< psubdiff >>
rect -255 60 -238 91
rect -255 -91 -238 -60
<< psubdiffcont >>
rect -255 -60 -238 60
<< poly >>
rect -175 57 175 65
rect -175 40 -167 57
rect 167 40 175 57
rect -175 21 175 40
rect -175 -40 175 -21
rect -175 -57 -167 -40
rect 167 -57 175 -40
rect -175 -65 175 -57
<< polycont >>
rect -167 40 167 57
rect -167 -57 167 -40
<< locali >>
rect -255 60 -238 91
rect -175 40 -167 57
rect 167 40 175 57
rect -198 15 -181 23
rect -198 -23 -181 -15
rect 181 15 198 23
rect 181 -23 198 -15
rect -175 -57 -167 -40
rect 167 -57 175 -40
rect -255 -91 -238 -60
<< viali >>
rect -167 40 167 57
rect -198 -15 -181 15
rect 181 -15 198 15
rect -167 -57 167 -40
<< metal1 >>
rect -173 57 173 60
rect -173 40 -167 57
rect 167 40 173 57
rect -173 37 173 40
rect -201 15 -178 21
rect -201 -15 -198 15
rect -181 -15 -178 15
rect -201 -21 -178 -15
rect 178 15 201 21
rect 178 -15 181 15
rect 198 -15 201 15
rect 178 -21 201 -15
rect -173 -40 173 -37
rect -173 -57 -167 -40
rect 167 -57 173 -40
rect -173 -60 173 -57
<< properties >>
string FIXED_BBOX -246 -99 246 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 3.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
