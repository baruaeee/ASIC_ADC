magic
tech sky130A
magscale 1 2
timestamp 1704301096
<< error_p >>
rect -29 129 29 135
rect -29 95 -17 129
rect -29 89 29 95
rect -29 -95 29 -89
rect -29 -129 -17 -95
rect -29 -135 29 -129
<< nwell >>
rect -211 -267 211 267
<< pmos >>
rect -15 -48 15 48
<< pdiff >>
rect -73 36 -15 48
rect -73 -36 -61 36
rect -27 -36 -15 36
rect -73 -48 -15 -36
rect 15 36 73 48
rect 15 -36 27 36
rect 61 -36 73 36
rect 15 -48 73 -36
<< pdiffc >>
rect -61 -36 -27 36
rect 27 -36 61 36
<< nsubdiff >>
rect -175 197 -79 231
rect 79 197 175 231
rect -175 135 -141 197
rect 141 135 175 197
rect -175 -197 -141 -135
rect 141 -197 175 -135
rect -175 -231 -79 -197
rect 79 -231 175 -197
<< nsubdiffcont >>
rect -79 197 79 231
rect -175 -135 -141 135
rect 141 -135 175 135
rect -79 -231 79 -197
<< poly >>
rect -33 129 33 145
rect -33 95 -17 129
rect 17 95 33 129
rect -33 79 33 95
rect -15 48 15 79
rect -15 -79 15 -48
rect -33 -95 33 -79
rect -33 -129 -17 -95
rect 17 -129 33 -95
rect -33 -145 33 -129
<< polycont >>
rect -17 95 17 129
rect -17 -129 17 -95
<< locali >>
rect -175 197 -79 231
rect 79 197 175 231
rect -175 135 -141 197
rect 141 135 175 197
rect -33 95 -17 129
rect 17 95 33 129
rect -61 36 -27 52
rect -61 -52 -27 -36
rect 27 36 61 52
rect 27 -52 61 -36
rect -33 -129 -17 -95
rect 17 -129 33 -95
rect -175 -197 -141 -135
rect 141 -197 175 -135
rect -175 -231 -79 -197
rect 79 -231 175 -197
<< viali >>
rect -17 95 17 129
rect -61 -36 -27 36
rect 27 -36 61 36
rect -17 -129 17 -95
<< metal1 >>
rect -29 129 29 135
rect -29 95 -17 129
rect 17 95 29 129
rect -29 89 29 95
rect -67 36 -21 48
rect -67 -36 -61 36
rect -27 -36 -21 36
rect -67 -48 -21 -36
rect 21 36 67 48
rect 21 -36 27 36
rect 61 -36 67 36
rect 21 -48 67 -36
rect -29 -95 29 -89
rect -29 -129 -17 -95
rect 17 -129 29 -95
rect -29 -135 29 -129
<< properties >>
string FIXED_BBOX -158 -214 158 214
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.48 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
