magic
tech sky130A
magscale 1 2
timestamp 1706479318
<< pwell >>
rect 620 -642 654 -582
<< psubdiff >>
rect 983 -718 1083 -684
<< locali >>
rect 735 454 827 488
rect 989 -718 1025 -684
rect 1059 -718 1075 -684
<< viali >>
rect 827 454 861 488
rect 1025 -718 1059 -684
<< metal1 >>
rect 726 500 826 502
rect 726 489 867 500
rect 401 488 867 489
rect 401 455 827 488
rect 401 374 435 455
rect 726 454 827 455
rect 861 454 867 488
rect 726 442 867 454
rect 726 436 826 442
rect 726 426 768 436
rect 392 274 492 374
rect 574 342 636 400
rect 762 384 768 426
rect 820 384 826 436
rect 963 406 1377 407
rect 962 372 1405 406
rect 963 341 1027 372
rect 1343 341 1405 372
rect 1076 279 1111 328
rect 401 142 435 274
rect 401 108 581 142
rect 631 117 665 209
rect 871 117 905 243
rect 1076 188 1115 279
rect 1249 188 1283 263
rect 1076 178 1111 188
rect 1283 178 1286 188
rect 1076 158 1286 178
rect 1080 146 1286 158
rect 631 83 905 117
rect 631 25 665 83
rect 397 -91 635 -57
rect 397 -126 431 -91
rect 396 -226 496 -126
rect 715 -223 749 83
rect 871 31 905 83
rect 1081 57 1115 146
rect 1249 67 1283 146
rect 1358 1 1392 2
rect 968 -27 1020 -21
rect 1339 -33 1403 1
rect 968 -85 1020 -79
rect 1358 -217 1393 -33
rect 1500 -217 1600 -200
rect 397 -609 431 -226
rect 715 -257 1125 -223
rect 715 -273 749 -257
rect 485 -307 749 -273
rect 485 -349 519 -307
rect 485 -471 520 -349
rect 485 -505 551 -471
rect 486 -531 551 -505
rect 892 -524 995 -490
rect 486 -532 520 -531
rect 620 -609 775 -581
rect 397 -615 775 -609
rect 397 -643 655 -615
rect 961 -652 995 -524
rect 1091 -567 1125 -257
rect 1358 -251 1600 -217
rect 1358 -482 1393 -251
rect 1500 -300 1600 -251
rect 1241 -517 1451 -482
rect 1518 -514 1570 -512
rect 924 -672 1024 -652
rect 924 -684 1065 -672
rect 924 -718 1025 -684
rect 1059 -718 1065 -684
rect 924 -719 1065 -718
rect 1304 -719 1338 -569
rect 1514 -574 1570 -514
rect 1514 -576 1566 -574
rect 924 -752 1338 -719
rect 977 -753 1338 -752
<< via1 >>
rect 768 384 820 436
rect 968 -79 1020 -27
<< metal2 >>
rect 768 436 820 442
rect 768 378 820 384
rect 776 -36 811 378
rect 962 -36 968 -27
rect 776 -71 968 -36
rect 962 -79 968 -71
rect 1020 -79 1026 -27
use sky130_fd_pr__nfet_01v8_2V6S9N  XM0
timestamp 1706236419
transform 1 0 722 0 1 -502
box -354 -252 354 252
use sky130_fd_pr__pfet_01v8_XYZSMQ  XM1
timestamp 1706236419
transform 1 0 605 0 1 147
box -211 -377 211 377
use sky130_fd_pr__pfet_01v8_AZD9DW  XM2
timestamp 1706479318
transform 0 -1 993 1 0 171
box -353 -261 353 261
use sky130_fd_pr__pfet_01v8_AZD9DW  XM3
timestamp 1706479318
transform 0 -1 1373 1 0 171
box -353 -261 353 261
use sky130_fd_pr__nfet_01v8_T8HSQ7  XM4
timestamp 1706236419
transform 0 -1 1325 1 0 -543
box -211 -367 211 367
<< labels >>
flabel metal1 924 -752 1024 -652 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 396 -226 496 -126 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 1500 -300 1600 -200 0 FreeSans 256 0 0 0 V09
port 1 nsew
flabel metal1 392 274 492 374 0 FreeSans 256 0 0 0 Vp
port 0 nsew
<< end >>
