magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< nwell >>
rect -2696 -261 2696 261
<< pmos >>
rect -2500 -42 2500 42
<< pdiff >>
rect -2558 30 -2500 42
rect -2558 -30 -2546 30
rect -2512 -30 -2500 30
rect -2558 -42 -2500 -30
rect 2500 30 2558 42
rect 2500 -30 2512 30
rect 2546 -30 2558 30
rect 2500 -42 2558 -30
<< pdiffc >>
rect -2546 -30 -2512 30
rect 2512 -30 2546 30
<< nsubdiff >>
rect -2660 191 -2564 225
rect 2564 191 2660 225
rect -2660 129 -2626 191
rect 2626 129 2660 191
rect -2660 -191 -2626 -129
rect 2626 -191 2660 -129
rect -2660 -225 -2564 -191
rect 2564 -225 2660 -191
<< nsubdiffcont >>
rect -2564 191 2564 225
rect -2660 -129 -2626 129
rect 2626 -129 2660 129
rect -2564 -225 2564 -191
<< poly >>
rect -2500 123 2500 139
rect -2500 89 -2484 123
rect 2484 89 2500 123
rect -2500 42 2500 89
rect -2500 -89 2500 -42
rect -2500 -123 -2484 -89
rect 2484 -123 2500 -89
rect -2500 -139 2500 -123
<< polycont >>
rect -2484 89 2484 123
rect -2484 -123 2484 -89
<< locali >>
rect -2660 191 -2564 225
rect 2564 191 2660 225
rect -2660 129 -2626 191
rect 2626 129 2660 191
rect -2500 89 -2484 123
rect 2484 89 2500 123
rect -2546 30 -2512 46
rect -2546 -46 -2512 -30
rect 2512 30 2546 46
rect 2512 -46 2546 -30
rect -2500 -123 -2484 -89
rect 2484 -123 2500 -89
rect -2660 -191 -2626 -129
rect 2626 -191 2660 -129
rect -2660 -225 -2564 -191
rect 2564 -225 2660 -191
<< viali >>
rect -2484 89 2484 123
rect -2546 -30 -2512 30
rect 2512 -30 2546 30
rect -2484 -123 2484 -89
<< metal1 >>
rect -2496 123 2496 129
rect -2496 89 -2484 123
rect 2484 89 2496 123
rect -2496 83 2496 89
rect -2552 30 -2506 42
rect -2552 -30 -2546 30
rect -2512 -30 -2506 30
rect -2552 -42 -2506 -30
rect 2506 30 2552 42
rect 2506 -30 2512 30
rect 2546 -30 2552 30
rect 2506 -42 2552 -30
rect -2496 -89 2496 -83
rect -2496 -123 -2484 -89
rect 2484 -123 2496 -89
rect -2496 -129 2496 -123
<< properties >>
string FIXED_BBOX -2643 -208 2643 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 25.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
