magic
tech sky130A
magscale 1 2
timestamp 1706204487
<< error_p >>
rect -29 231 29 237
rect -29 197 -17 231
rect -29 191 29 197
rect -29 -197 29 -191
rect -29 -231 -17 -197
rect -29 -237 29 -231
<< nwell >>
rect -211 -369 211 369
<< pmos >>
rect -15 -150 15 150
<< pdiff >>
rect -73 138 -15 150
rect -73 -138 -61 138
rect -27 -138 -15 138
rect -73 -150 -15 -138
rect 15 138 73 150
rect 15 -138 27 138
rect 61 -138 73 138
rect 15 -150 73 -138
<< pdiffc >>
rect -61 -138 -27 138
rect 27 -138 61 138
<< nsubdiff >>
rect -141 -333 -79 -299
rect 79 -333 141 -299
<< nsubdiffcont >>
rect -79 -333 79 -299
<< poly >>
rect -33 231 33 247
rect -33 197 -17 231
rect 17 197 33 231
rect -33 181 33 197
rect -15 150 15 181
rect -15 -181 15 -150
rect -33 -197 33 -181
rect -33 -231 -17 -197
rect 17 -231 33 -197
rect -33 -247 33 -231
<< polycont >>
rect -17 197 17 231
rect -17 -231 17 -197
<< locali >>
rect -33 197 -17 231
rect 17 197 33 231
rect -61 138 -27 154
rect -61 -154 -27 -138
rect 27 138 61 154
rect 27 -154 61 -138
rect -33 -231 -17 -197
rect 17 -231 33 -197
rect -141 -333 -79 -299
rect 79 -333 141 -299
<< viali >>
rect -17 197 17 231
rect -61 -138 -27 138
rect 27 -138 61 138
rect -17 -231 17 -197
<< metal1 >>
rect -29 231 29 237
rect -29 197 -17 231
rect 17 197 29 231
rect -29 191 29 197
rect -67 138 -21 150
rect -67 -138 -61 138
rect -27 -138 -21 138
rect -67 -150 -21 -138
rect 21 138 67 150
rect 21 -138 27 138
rect 61 -138 67 138
rect 21 -150 67 -138
rect -29 -197 29 -191
rect -29 -231 -17 -197
rect 17 -231 29 -197
rect -29 -237 29 -231
<< properties >>
string FIXED_BBOX -158 -316 158 316
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
