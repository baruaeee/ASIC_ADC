magic
tech sky130A
magscale 1 2
timestamp 1704418840
<< nwell >>
rect -335 -261 335 261
<< pmos >>
rect -139 -42 139 42
<< pdiff >>
rect -197 30 -139 42
rect -197 -30 -185 30
rect -151 -30 -139 30
rect -197 -42 -139 -30
rect 139 30 197 42
rect 139 -30 151 30
rect 185 -30 197 30
rect 139 -42 197 -30
<< pdiffc >>
rect -185 -30 -151 30
rect 151 -30 185 30
<< nsubdiff >>
rect -299 191 -203 225
rect 203 191 299 225
rect -299 129 -265 191
rect 265 129 299 191
rect -299 -191 -265 -129
rect 265 -191 299 -129
rect -299 -225 -203 -191
rect 203 -225 299 -191
<< nsubdiffcont >>
rect -203 191 203 225
rect -299 -129 -265 129
rect 265 -129 299 129
rect -203 -225 203 -191
<< poly >>
rect -139 123 139 139
rect -139 89 -123 123
rect 123 89 139 123
rect -139 42 139 89
rect -139 -89 139 -42
rect -139 -123 -123 -89
rect 123 -123 139 -89
rect -139 -139 139 -123
<< polycont >>
rect -123 89 123 123
rect -123 -123 123 -89
<< locali >>
rect -299 191 -203 225
rect 203 191 299 225
rect -299 129 -265 191
rect 265 129 299 191
rect -139 89 -123 123
rect 123 89 139 123
rect -185 30 -151 46
rect -185 -46 -151 -30
rect 151 30 185 46
rect 151 -46 185 -30
rect -139 -123 -123 -89
rect 123 -123 139 -89
rect -299 -191 -265 -129
rect 265 -191 299 -129
rect -299 -225 -203 -191
rect 203 -225 299 -191
<< viali >>
rect -123 89 123 123
rect -185 -30 -151 30
rect 151 -30 185 30
rect -123 -123 123 -89
<< metal1 >>
rect -135 123 135 129
rect -135 89 -123 123
rect 123 89 135 123
rect -135 83 135 89
rect -191 30 -145 42
rect -191 -30 -185 30
rect -151 -30 -145 30
rect -191 -42 -145 -30
rect 145 30 191 42
rect 145 -30 151 30
rect 185 -30 191 30
rect 145 -42 191 -30
rect -135 -89 135 -83
rect -135 -123 -123 -89
rect 123 -123 135 -89
rect -135 -129 135 -123
<< properties >>
string FIXED_BBOX -282 -208 282 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 1.39 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
