// This is the unpowered netlist.
module ADC (b,
    p);
 output [3:0] b;
 input [14:0] p;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__decap_4 FILLER_0_0_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__or3_1 _26_ (.A(net5),
    .B(net4),
    .C(net6),
    .X(_00_));
 sky130_fd_sc_hd__or4_1 _27_ (.A(net14),
    .B(net15),
    .C(net3),
    .D(net2),
    .X(_01_));
 sky130_fd_sc_hd__nor2_1 _28_ (.A(_00_),
    .B(_01_),
    .Y(_02_));
 sky130_fd_sc_hd__or3_1 _29_ (.A(net11),
    .B(net13),
    .C(net12),
    .X(_03_));
 sky130_fd_sc_hd__or4b_1 _30_ (.A(net9),
    .B(net10),
    .C(_03_),
    .D_N(net1),
    .X(_04_));
 sky130_fd_sc_hd__xor2_1 _31_ (.A(net7),
    .B(net8),
    .X(_05_));
 sky130_fd_sc_hd__and4_1 _32_ (.A(net7),
    .B(net1),
    .C(net9),
    .D(net8),
    .X(_06_));
 sky130_fd_sc_hd__and3b_1 _33_ (.A_N(net13),
    .B(_06_),
    .C(net10),
    .X(_07_));
 sky130_fd_sc_hd__xnor2_1 _34_ (.A(net11),
    .B(net12),
    .Y(_08_));
 sky130_fd_sc_hd__a2bb2o_1 _35_ (.A1_N(_04_),
    .A2_N(_05_),
    .B1(_07_),
    .B2(_08_),
    .X(_09_));
 sky130_fd_sc_hd__and4_1 _36_ (.A(net11),
    .B(net10),
    .C(net13),
    .D(net12),
    .X(_10_));
 sky130_fd_sc_hd__and4_1 _37_ (.A(net14),
    .B(net15),
    .C(net3),
    .D(net2),
    .X(_11_));
 sky130_fd_sc_hd__and4_1 _38_ (.A(net4),
    .B(_06_),
    .C(_10_),
    .D(_11_),
    .X(_12_));
 sky130_fd_sc_hd__xnor2_1 _39_ (.A(net5),
    .B(net6),
    .Y(_13_));
 sky130_fd_sc_hd__nor4_1 _40_ (.A(net15),
    .B(net3),
    .C(net2),
    .D(_00_),
    .Y(_14_));
 sky130_fd_sc_hd__and2_1 _41_ (.A(_06_),
    .B(_10_),
    .X(_15_));
 sky130_fd_sc_hd__and3b_1 _42_ (.A_N(net3),
    .B(net15),
    .C(net14),
    .X(_16_));
 sky130_fd_sc_hd__and4b_1 _43_ (.A_N(_00_),
    .B(_06_),
    .C(_10_),
    .D(_16_),
    .X(_17_));
 sky130_fd_sc_hd__a32o_1 _44_ (.A1(net14),
    .A2(_14_),
    .A3(_15_),
    .B1(_17_),
    .B2(net2),
    .X(_18_));
 sky130_fd_sc_hd__a221o_1 _45_ (.A1(_02_),
    .A2(_09_),
    .B1(_12_),
    .B2(_13_),
    .C1(_18_),
    .X(net16));
 sky130_fd_sc_hd__inv_2 _46_ (.A(_04_),
    .Y(_19_));
 sky130_fd_sc_hd__a21o_1 _47_ (.A1(net5),
    .A2(_12_),
    .B1(_17_),
    .X(_20_));
 sky130_fd_sc_hd__and3_1 _48_ (.A(net11),
    .B(_02_),
    .C(_07_),
    .X(_21_));
 sky130_fd_sc_hd__a311o_1 _49_ (.A1(net7),
    .A2(_02_),
    .A3(_19_),
    .B1(_20_),
    .C1(_21_),
    .X(net17));
 sky130_fd_sc_hd__and4bb_1 _50_ (.A_N(net5),
    .B_N(net6),
    .C(_15_),
    .D(_11_),
    .X(_22_));
 sky130_fd_sc_hd__inv_2 _51_ (.A(_03_),
    .Y(_23_));
 sky130_fd_sc_hd__a32o_1 _52_ (.A1(_02_),
    .A2(_06_),
    .A3(_23_),
    .B1(_12_),
    .B2(net5),
    .X(_24_));
 sky130_fd_sc_hd__or3_1 _53_ (.A(_21_),
    .B(_22_),
    .C(_24_),
    .X(_25_));
 sky130_fd_sc_hd__clkbuf_1 _54_ (.A(_25_),
    .X(net18));
 sky130_fd_sc_hd__a211o_1 _55_ (.A1(_14_),
    .A2(_15_),
    .B1(_20_),
    .C1(_22_),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(p[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(p[4]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(p[5]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(p[6]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(p[7]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(p[8]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(p[9]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input2 (.A(p[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(p[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(p[12]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(p[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(p[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(p[1]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(p[2]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(p[3]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output16 (.A(net16),
    .X(b[0]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(b[1]));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(b[2]));
 sky130_fd_sc_hd__clkbuf_4 output19 (.A(net19),
    .X(b[3]));
endmodule

