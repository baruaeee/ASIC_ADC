magic
tech sky130A
magscale 1 2
timestamp 1706211875
<< nwell >>
rect 0 0 516 1512
<< pmos >>
rect 200 420 230 714
rect 286 420 316 714
<< pdiff >>
rect 147 606 200 714
rect 147 572 155 606
rect 189 572 200 606
rect 147 538 200 572
rect 147 504 155 538
rect 189 504 200 538
rect 147 470 200 504
rect 147 436 155 470
rect 189 436 200 470
rect 147 420 200 436
rect 230 606 286 714
rect 230 572 241 606
rect 275 572 286 606
rect 230 538 286 572
rect 230 504 241 538
rect 275 504 286 538
rect 230 470 286 504
rect 230 436 241 470
rect 275 436 286 470
rect 230 420 286 436
rect 316 606 369 714
rect 316 572 327 606
rect 361 572 369 606
rect 316 538 369 572
rect 316 504 327 538
rect 361 504 369 538
rect 316 470 369 504
rect 316 436 327 470
rect 361 436 369 470
rect 316 420 369 436
<< pdiffc >>
rect 155 572 189 606
rect 155 504 189 538
rect 155 436 189 470
rect 241 572 275 606
rect 241 504 275 538
rect 241 436 275 470
rect 327 572 361 606
rect 327 504 361 538
rect 327 436 361 470
<< nsubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
<< nsubdiffcont >>
rect 241 1327 275 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 714 230 897
rect 286 714 316 897
rect 200 252 230 420
rect 286 252 316 420
<< polycont >>
rect 241 907 275 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 147 606 197 773
rect 147 572 155 606
rect 189 572 197 606
rect 147 538 197 572
rect 147 504 155 538
rect 189 504 197 538
rect 147 470 197 504
rect 147 436 155 470
rect 189 436 197 470
rect 147 185 197 436
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 606 283 773
rect 233 572 241 606
rect 275 572 283 606
rect 233 538 283 572
rect 233 504 241 538
rect 275 504 283 538
rect 233 470 283 504
rect 233 436 241 470
rect 275 436 283 470
rect 233 101 283 436
rect 233 67 241 101
rect 275 67 283 101
rect 319 606 369 773
rect 319 572 327 606
rect 361 572 369 606
rect 319 538 369 572
rect 319 504 327 538
rect 361 504 369 538
rect 319 470 369 504
rect 319 436 327 470
rect 361 436 369 470
rect 319 185 369 436
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
<< viali >>
rect 241 1327 275 1361
rect 241 907 275 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
<< metal1 >>
rect 138 1370 378 1372
rect 138 1361 318 1370
rect 138 1327 241 1361
rect 275 1327 318 1361
rect 138 1318 318 1327
rect 370 1318 378 1370
rect 138 1316 378 1318
rect 52 941 292 952
rect 52 907 241 941
rect 275 907 292 941
rect 52 896 292 907
rect 138 194 378 196
rect 138 185 318 194
rect 138 151 155 185
rect 189 151 318 185
rect 138 142 318 151
rect 370 142 378 194
rect 138 140 378 142
rect 52 101 292 112
rect 52 67 241 101
rect 275 67 292 101
rect 52 56 292 67
<< via1 >>
rect 318 1318 370 1370
rect 318 185 370 194
rect 318 151 327 185
rect 327 151 361 185
rect 361 151 370 185
rect 318 142 370 151
<< metal2 >>
rect 316 1370 372 1376
rect 316 1318 318 1370
rect 370 1318 372 1370
rect 316 194 372 1318
rect 316 142 318 194
rect 370 142 372 194
rect 316 136 372 142
<< end >>
