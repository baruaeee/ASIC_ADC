magic
tech sky130A
magscale 1 2
timestamp 1706216322
<< error_p >>
rect -29 181 29 187
rect -29 147 -17 181
rect -29 141 29 147
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect -29 -187 29 -181
<< nwell >>
rect -212 -319 212 319
<< pmos >>
rect -16 -100 16 100
<< pdiff >>
rect -74 88 -16 100
rect -74 -88 -62 88
rect -28 -88 -16 88
rect -74 -100 -16 -88
rect 16 88 74 100
rect 16 -88 28 88
rect 62 -88 74 88
rect 16 -100 74 -88
<< pdiffc >>
rect -62 -88 -28 88
rect 28 -88 62 88
<< nsubdiff >>
rect -142 249 -80 283
rect 80 249 142 283
<< nsubdiffcont >>
rect -80 249 80 283
<< poly >>
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect -16 100 16 131
rect -16 -131 16 -100
rect -33 -147 33 -131
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -197 33 -181
<< polycont >>
rect -17 147 17 181
rect -17 -181 17 -147
<< locali >>
rect -142 249 -80 283
rect 80 249 142 283
rect -33 147 -17 181
rect 17 147 33 181
rect -62 88 -28 104
rect -62 -104 -28 -88
rect 28 88 62 104
rect 28 -104 62 -88
rect -33 -181 -17 -147
rect 17 -181 33 -147
<< viali >>
rect -17 147 17 181
rect -62 -88 -28 88
rect 28 -88 62 88
rect -17 -181 17 -147
<< metal1 >>
rect -29 181 29 187
rect -29 147 -17 181
rect 17 147 29 181
rect -29 141 29 147
rect -68 88 -22 100
rect -68 -88 -62 88
rect -28 -88 -22 88
rect -68 -100 -22 -88
rect 22 88 68 100
rect 22 -88 28 88
rect 62 -88 68 88
rect 22 -100 68 -88
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect 17 -181 29 -147
rect -29 -187 29 -181
<< properties >>
string FIXED_BBOX -159 -266 159 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.156 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
