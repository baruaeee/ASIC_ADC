* NGSPICE file created from th05.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_ATLS57 a_15_n200# a_n175_n374# a_n73_n200# a_n33_n288#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n175_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n73_n200# a_n33_n288# 0.0312f
C1 a_n73_n200# a_15_n200# 0.321f
C2 a_15_n200# a_n33_n288# 0.0312f
C3 a_15_n200# a_n175_n374# 0.233f
C4 a_n73_n200# a_n175_n374# 0.233f
C5 a_n33_n288# a_n175_n374# 0.347f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GC6 a_200_n42# w_n396_n261# a_n200_n139# a_n258_n42#
+ VSUBS
X0 a_200_n42# a_n200_n139# a_n258_n42# w_n396_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 w_n396_n261# a_n200_n139# 0.743f
C1 a_200_n42# a_n258_n42# 0.0134f
C2 a_200_n42# a_n200_n139# 0.0196f
C3 a_n200_n139# a_n258_n42# 0.0196f
C4 a_200_n42# w_n396_n261# 0.0498f
C5 w_n396_n261# a_n258_n42# 0.0498f
C6 a_200_n42# VSUBS 0.0338f
C7 a_n258_n42# VSUBS 0.0338f
C8 a_n200_n139# VSUBS 0.554f
C9 w_n396_n261# VSUBS 1.79f
.ends

.subckt sky130_fd_pr__pfet_01v8_PZD9SE a_n112_n139# w_n308_n261# a_112_n42# a_n170_n42#
+ VSUBS
X0 a_112_n42# a_n112_n139# a_n170_n42# w_n308_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.12
C0 a_n170_n42# a_n112_n139# 0.0153f
C1 a_112_n42# w_n308_n261# 0.0499f
C2 a_n112_n139# a_112_n42# 0.0153f
C3 a_n112_n139# w_n308_n261# 0.472f
C4 a_n170_n42# a_112_n42# 0.0219f
C5 a_n170_n42# w_n308_n261# 0.0499f
C6 a_112_n42# VSUBS 0.0318f
C7 a_n170_n42# VSUBS 0.0318f
C8 a_n112_n139# VSUBS 0.332f
C9 w_n308_n261# VSUBS 1.43f
.ends

.subckt sky130_fd_pr__nfet_01v8_UNLS3X a_n33_n200# a_n175_n286# a_n73_n112# a_15_n112#
X0 a_15_n112# a_n33_n200# a_n73_n112# a_n175_n286# sky130_fd_pr__nfet_01v8 ad=0.325 pd=2.82 as=0.325 ps=2.82 w=1.12 l=0.15
C0 a_n33_n200# a_n73_n112# 0.0262f
C1 a_n73_n112# a_15_n112# 0.181f
C2 a_n33_n200# a_15_n112# 0.0262f
C3 a_15_n112# a_n175_n286# 0.144f
C4 a_n73_n112# a_n175_n286# 0.144f
C5 a_n33_n200# a_n175_n286# 0.344f
.ends

.subckt th05 Vp V05 Vin Vn
XXM0 m1_836_n724# Vn Vn Vin sky130_fd_pr__nfet_01v8_ATLS57
XXM1 m1_836_n724# Vp Vin Vp Vn sky130_fd_pr__pfet_01v8_VZ9GC6
XXM2 m1_836_n724# Vp V05 Vp Vn sky130_fd_pr__pfet_01v8_PZD9SE
XXM3 m1_836_n724# Vn Vn V05 sky130_fd_pr__nfet_01v8_UNLS3X
C0 m1_836_n724# V05 0.122f
C1 Vin V05 5.09e-20
C2 m1_836_n724# Vin 0.187f
C3 Vp V05 0.103f
C4 m1_836_n724# Vp 0.372f
C5 Vin Vp 0.324f
C6 Vin Vn 1.06f
C7 V05 Vn 0.48f
C8 m1_836_n724# Vn 1.23f
C9 Vp Vn 3.53f
.ends

