* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : pre_therm                                    *
* Netlisted  : Mon Dec  9 01:54:35 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733705663440                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733705663440 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6.5e-07 W=4.45e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733705663440

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733705663441                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733705663441 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=6.3e-07 W=7.9e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733705663441

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv01f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv01f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_733705663440 $T=295 475 0 0 $X=-110 $Y=325
X5 VDD Y A pfet_01v8_CDNS_733705663441 $T=295 2820 0 0 $X=-150 $Y=2640
.ends inv01f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733705663442                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733705663442 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 pfet_01v8 L=1.05e-06 W=5.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733705663442

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733705663443                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733705663443 1 2 3 4
** N=10 EP=4 FDC=1
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=1.02e-06 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733705663443

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: preampF                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt preampF VDD VSS A Y
** N=9 EP=4 FDC=2
X5 Y VSS A VDD pfet_01v8_CDNS_733705663442 $T=825 3430 0 270 $X=645 $Y=1935
X6 Y VDD A VSS nfet_01v8_CDNS_733705663443 $T=430 485 1 180 $X=-125 $Y=335
.ends preampF

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733705663444                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733705663444 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.5e-07 W=8e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733705663444

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733705663445                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733705663445 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=2.85e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733705663445

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv02f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv02f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VDD Y A pfet_01v8_CDNS_733705663444 $T=335 2855 0 0 $X=-110 $Y=2675
X5 VSS Y A nfet_01v8_CDNS_733705663445 $T=315 640 0 0 $X=-90 $Y=490
.ends inv02f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733705663446                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733705663446 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 pfet_01v8 L=2.5e-07 W=5.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733705663446

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733705663447                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733705663447 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 nfet_01v8 L=5.5e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733705663447

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: preamp1F                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt preamp1F VDD VSS A Y
** N=9 EP=4 FDC=2
X3 Y VSS A VDD pfet_01v8_CDNS_733705663446 $T=840 2840 0 90 $X=110 $Y=2395
X4 Y VDD A VSS nfet_01v8_CDNS_733705663447 $T=610 1275 0 270 $X=460 $Y=320
.ends preamp1F

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733705663448                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733705663448 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=3.5e-07 W=6.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733705663448

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733705663449                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733705663449 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=4.5e-07 W=6.4e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733705663449

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv03f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv03f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VDD Y A pfet_01v8_CDNS_733705663448 $T=335 3045 0 0 $X=-110 $Y=2865
X5 VSS Y A nfet_01v8_CDNS_733705663449 $T=290 640 0 0 $X=-115 $Y=490
.ends inv03f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634410                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634410 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.9e-07 W=6.2e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634410

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634411                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634411 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6e-07 W=7.05e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634411

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv04f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv04f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VDD Y A pfet_01v8_CDNS_7337056634410 $T=380 2650 0 0 $X=-65 $Y=2470
X5 VSS Y A nfet_01v8_CDNS_7337056634411 $T=280 715 0 0 $X=-125 $Y=565
.ends inv04f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634412                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634412 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=6.95e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634412

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634413                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634413 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=4e-07 W=6.5e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634413

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv05f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv05f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VDD Y A pfet_01v8_CDNS_7337056634412 $T=360 2825 0 0 $X=-85 $Y=2645
X5 VSS Y A nfet_01v8_CDNS_7337056634413 $T=315 630 0 0 $X=-90 $Y=480
.ends inv05f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634414                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634414 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3.2e-07 W=7.25e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634414

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634415                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634415 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=4.35e-07 W=5.6e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634415

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv06f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv06f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7337056634414 $T=395 685 0 0 $X=-10 $Y=535
X5 VDD Y A pfet_01v8_CDNS_7337056634415 $T=335 3005 0 0 $X=-110 $Y=2825
.ends inv06f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634416                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634416 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3e-07 W=9.8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634416

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634417                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634417 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.55e-07 W=5.7e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634417

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv07f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv07f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7337056634416 $T=315 460 0 0 $X=-90 $Y=310
X5 VDD Y A pfet_01v8_CDNS_7337056634417 $T=360 2950 0 0 $X=-85 $Y=2770
.ends inv07f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634418                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634418 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=9.9e-07 W=4.9e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634418

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634419                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634419 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.65e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634419

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv08f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv08f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7337056634418 $T=1280 740 0 90 $X=640 $Y=335
X5 VDD Y A pfet_01v8_CDNS_7337056634419 $T=360 2755 0 0 $X=-85 $Y=2575
.ends inv08f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634420                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634420 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.1e-06 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634420

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634421                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634421 1 2 3
** N=9 EP=3 FDC=2
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.7e-07 $X=0 $Y=0 $dt=8
M1 1 3 2 1 pfet_01v8 L=1.5e-07 W=7.7e-07 $X=430 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634421

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv09f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv09f VDD VSS A Y
** N=9 EP=4 FDC=3
X4 VSS Y A nfet_01v8_CDNS_7337056634420 $T=905 695 0 90 $X=335 $Y=290
X5 VDD Y A pfet_01v8_CDNS_7337056634421 $T=400 2840 0 0 $X=-45 $Y=2660
.ends inv09f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634422                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634422 1 2 3
** N=7 EP=3 FDC=1
M0 2 2 1 3 pfet_01v8 L=1.5e-07 W=1e-06 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634422

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: div_fixed                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt div_fixed A VSS Y
** N=8 EP=3 FDC=2
X4 A Y VSS A pfet_01v8_CDNS_733705663442 $T=1625 3880 1 270 $X=895 $Y=2385
X5 Y VSS A pfet_01v8_CDNS_7337056634422 $T=470 1900 0 180 $X=-125 $Y=720
.ends div_fixed

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634423                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634423 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.55e-07 W=9.45e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634423

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634424                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634424 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.45e-07 W=8.65e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634424

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv10f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv10f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7337056634423 $T=425 555 0 0 $X=20 $Y=405
X5 VDD Y A pfet_01v8_CDNS_7337056634424 $T=385 2670 0 0 $X=-60 $Y=2490
.ends inv10f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634425                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634425 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=9.5e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634425

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634426                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634426 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.6e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634426

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv11f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv11f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7337056634425 $T=215 700 0 0 $X=-190 $Y=550
X5 VDD Y A pfet_01v8_CDNS_7337056634426 $T=350 2610 0 0 $X=-95 $Y=2430
.ends inv11f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634427                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634427 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3.3e-07 W=8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634427

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634428                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634428 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634428

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv12f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv12f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7337056634427 $T=340 555 0 0 $X=-65 $Y=405
X5 VDD Y A pfet_01v8_CDNS_7337056634428 $T=385 2785 0 0 $X=-60 $Y=2605
.ends inv12f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634429                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634429 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=5.5e-07 W=5.4e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634429

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634430                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634430 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.6e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634430

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv13f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv13f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7337056634429 $T=360 720 0 0 $X=-45 $Y=570
X5 VDD Y A pfet_01v8_CDNS_7337056634430 $T=385 2685 0 0 $X=-60 $Y=2505
.ends inv13f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7337056634431                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7337056634431 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6.75e-07 W=4.8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7337056634431

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634432                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634432 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.65e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634432

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv14f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv14f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7337056634431 $T=350 675 0 0 $X=-55 $Y=525
X5 VDD Y A pfet_01v8_CDNS_7337056634432 $T=445 2705 0 0 $X=0 $Y=2525
.ends inv14f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7337056634433                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7337056634433 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7337056634433

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv15f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv15f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7337056634425 $T=215 700 0 0 $X=-190 $Y=550
X5 VDD Y A pfet_01v8_CDNS_7337056634433 $T=620 2635 0 0 $X=175 $Y=2455
.ends inv15f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pre_therm                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pre_therm IN VDD VSS Y01 Y02 Y03 Y04 Y05 Y06 Y07
+ Y08 Y09 Y10 Y11 Y12 Y13 Y14 Y15
** N=21 EP=18 FDC=37
X54 VDD VSS 2 Y01 inv01f $T=1740 9060 1 0 $X=1560 $Y=4615
X55 VDD VSS IN 2 preampF $T=0 9060 1 0 $X=-180 $Y=4615
X56 VDD VSS 2 Y02 inv02f $T=3480 9060 1 0 $X=3300 $Y=4615
X57 VDD VSS IN 3 preamp1F $T=0 255 0 0 $X=-180 $Y=-10
X58 VDD VSS 3 Y03 inv03f $T=1740 260 0 0 $X=1560 $Y=-5
X59 VDD VSS 3 Y04 inv04f $T=3480 260 0 0 $X=3300 $Y=-5
X60 VDD VSS 3 Y05 inv05f $T=5220 260 0 0 $X=5040 $Y=-5
X61 VDD VSS IN Y06 inv06f $T=6960 260 0 0 $X=6780 $Y=-5
X62 VDD VSS IN Y07 inv07f $T=8700 260 0 0 $X=8520 $Y=-5
X63 VDD VSS IN Y08 inv08f $T=5220 9060 1 0 $X=5040 $Y=4615
X64 VDD VSS IN Y09 inv09f $T=6970 9060 1 0 $X=6780 $Y=4615
X65 IN VSS 8 div_fixed $T=0 9580 0 0 $X=-180 $Y=9315
X66 VDD VSS 8 Y10 inv10f $T=4040 9585 0 0 $X=3860 $Y=9320
X67 VDD VSS 8 Y11 inv11f $T=5735 9585 0 0 $X=5545 $Y=9320
X68 VDD VSS 8 Y12 inv12f $T=7430 9580 0 0 $X=7250 $Y=9315
X69 VDD VSS 8 Y13 inv13f $T=9060 9580 0 0 $X=8880 $Y=9315
X70 VDD VSS 8 Y14 inv14f $T=8665 9060 1 0 $X=8485 $Y=4615
X71 VDD VSS 8 Y15 inv15f $T=10360 9060 1 0 $X=10170 $Y=4615
.ends pre_therm
