module therm ( VNB, VPWR, clk, rst, p, b);

input VNB, VPWR;
input clk;
input rst;
input [14:0] p;
output [3:0] b;

sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_1 ( .VNB(VNB), .VPWR(VPWR), .A(_47__2_), .X(b[2]) );
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_2 ( .VNB(VNB), .VPWR(VPWR), .A(_47__3_), .X(b[3]) );
sky130_fd_sc_hd__dfrtp_1 sky130_fd_sc_hd__dfrtp_1_1 ( .VNB(VNB), .VPWR(VPWR), .CLK(clk), .D(_0__0_), .Q(_47__0_), .RESET_B(_1_) );
sky130_fd_sc_hd__dfrtp_1 sky130_fd_sc_hd__dfrtp_1_2 ( .VNB(VNB), .VPWR(VPWR), .CLK(clk), .D(_0__1_), .Q(_47__1_), .RESET_B(_1_) );
sky130_fd_sc_hd__dfrtp_1 sky130_fd_sc_hd__dfrtp_1_3 ( .VNB(VNB), .VPWR(VPWR), .CLK(clk), .D(_0__2_), .Q(_47__2_), .RESET_B(_1_) );
sky130_fd_sc_hd__dfrtp_1 sky130_fd_sc_hd__dfrtp_1_4 ( .VNB(VNB), .VPWR(VPWR), .CLK(clk), .D(_0__3_), .Q(_47__3_), .RESET_B(_1_) );
sky130_fd_sc_hd__nor3_4 sky130_fd_sc_hd__nor3_4_1 ( .VNB(VNB), .VPWR(VPWR), .A(p[12]), .B(p[13]), .C(p[14]), .Y(_2_) );
sky130_fd_sc_hd__nor2_1 sky130_fd_sc_hd__nor2_1_1 ( .VNB(VNB), .VPWR(VPWR), .A(p[10]), .B(p[11]), .Y(_3_) );
sky130_fd_sc_hd__nor2_1 sky130_fd_sc_hd__nor2_1_2 ( .VNB(VNB), .VPWR(VPWR), .A(p[8]), .B(p[9]), .Y(_4_) );
sky130_fd_sc_hd__nand3_1 sky130_fd_sc_hd__nand3_1_1 ( .VNB(VNB), .VPWR(VPWR), .A(_2_), .B(_3_), .C(_4_), .Y(_5_) );
sky130_fd_sc_hd__nand4_1 sky130_fd_sc_hd__nand4_1_1 ( .VNB(VNB), .VPWR(VPWR), .A(p[0]), .B(p[1]), .C(p[2]), .D(p[3]), .Y(_6_) );
sky130_fd_sc_hd__clkinv_1 sky130_fd_sc_hd__clkinv_1_1 ( .VNB(VNB), .VPWR(VPWR), .A(_6_), .Y(_7_) );
sky130_fd_sc_hd__clkinv_1 sky130_fd_sc_hd__clkinv_1_2 ( .VNB(VNB), .VPWR(VPWR), .A(p[5]), .Y(_8_) );
sky130_fd_sc_hd__clkinv_1 sky130_fd_sc_hd__clkinv_1_3 ( .VNB(VNB), .VPWR(VPWR), .A(p[6]), .Y(_9_) );
sky130_fd_sc_hd__clkinv_1 sky130_fd_sc_hd__clkinv_1_4 ( .VNB(VNB), .VPWR(VPWR), .A(p[7]), .Y(_10_) );
sky130_fd_sc_hd__nand4_1 sky130_fd_sc_hd__nand4_1_2 ( .VNB(VNB), .VPWR(VPWR), .A(_8_), .B(_9_), .C(_10_), .D(p[4]), .Y(_11_) );
sky130_fd_sc_hd__nand2_1 sky130_fd_sc_hd__nand2_1_1 ( .VNB(VNB), .VPWR(VPWR), .A(p[4]), .B(p[5]), .Y(_12_) );
sky130_fd_sc_hd__nand2_1 sky130_fd_sc_hd__nand2_1_2 ( .VNB(VNB), .VPWR(VPWR), .A(_10_), .B(p[6]), .Y(_13_) );
sky130_fd_sc_hd__o21ai_0 sky130_fd_sc_hd__o21ai_0_1 ( .VNB(VNB), .VPWR(VPWR), .A1(_12_), .A2(_13_), .B1(_11_), .Y(_14_) );
sky130_fd_sc_hd__nand2_1 sky130_fd_sc_hd__nand2_1_3 ( .VNB(VNB), .VPWR(VPWR), .A(p[1]), .B(p[2]), .Y(_15_) );
sky130_fd_sc_hd__or2_2 sky130_fd_sc_hd__or2_2_1 ( .VNB(VNB), .VPWR(VPWR), .A(p[1]), .B(p[2]), .X(_16_) );
sky130_fd_sc_hd__nand2_1 sky130_fd_sc_hd__nand2_1_4 ( .VNB(VNB), .VPWR(VPWR), .A(_16_), .B(_15_), .Y(_17_) );
sky130_fd_sc_hd__nor3_1 sky130_fd_sc_hd__nor3_1_1 ( .VNB(VNB), .VPWR(VPWR), .A(p[5]), .B(p[6]), .C(p[7]), .Y(_18_) );
sky130_fd_sc_hd__nor3b_1 sky130_fd_sc_hd__nor3b_1_1 ( .VNB(VNB), .VPWR(VPWR), .A(p[3]), .B(p[4]), .C_N(p[0]), .Y(_19_) );
sky130_fd_sc_hd__a32oi_1 sky130_fd_sc_hd__a32oi_1_1 ( .VNB(VNB), .VPWR(VPWR), .A1(_17_), .A2(_18_), .A3(_19_), .B1(_14_), .B2(_7_), .Y(_20_) );
sky130_fd_sc_hd__nor4_1 sky130_fd_sc_hd__nor4_1_1 ( .VNB(VNB), .VPWR(VPWR), .A(_9_), .B(_10_), .C(_12_), .D(_6_), .Y(_21_) );
sky130_fd_sc_hd__nor2_1 sky130_fd_sc_hd__nor2_1_3 ( .VNB(VNB), .VPWR(VPWR), .A(p[13]), .B(p[14]), .Y(_22_) );
sky130_fd_sc_hd__nand2_1 sky130_fd_sc_hd__nand2_1_5 ( .VNB(VNB), .VPWR(VPWR), .A(p[8]), .B(p[9]), .Y(_23_) );
sky130_fd_sc_hd__nand2_1 sky130_fd_sc_hd__nand2_1_6 ( .VNB(VNB), .VPWR(VPWR), .A(p[10]), .B(p[11]), .Y(_24_) );
sky130_fd_sc_hd__nor2_1 sky130_fd_sc_hd__nor2_1_4 ( .VNB(VNB), .VPWR(VPWR), .A(_23_), .B(_24_), .Y(_25_) );
sky130_fd_sc_hd__and2_2 sky130_fd_sc_hd__and2_2_1 ( .VNB(VNB), .VPWR(VPWR), .A(p[13]), .B(p[14]), .X(_26_) );
sky130_fd_sc_hd__o211ai_1 sky130_fd_sc_hd__o211ai_1_1 ( .VNB(VNB), .VPWR(VPWR), .A1(_22_), .A2(_26_), .B1(p[12]), .C1(_25_), .Y(_27_) );
sky130_fd_sc_hd__clkinv_1 sky130_fd_sc_hd__clkinv_1_5 ( .VNB(VNB), .VPWR(VPWR), .A(p[9]), .Y(_28_) );
sky130_fd_sc_hd__nand4_1 sky130_fd_sc_hd__nand4_1_3 ( .VNB(VNB), .VPWR(VPWR), .A(_2_), .B(p[8]), .C(_28_), .D(_3_), .Y(_29_) );
sky130_fd_sc_hd__clkinv_1 sky130_fd_sc_hd__clkinv_1_6 ( .VNB(VNB), .VPWR(VPWR), .A(p[11]), .Y(_30_) );
sky130_fd_sc_hd__and2_2 sky130_fd_sc_hd__and2_2_2 ( .VNB(VNB), .VPWR(VPWR), .A(p[8]), .B(p[9]), .X(_31_) );
sky130_fd_sc_hd__nand4_1 sky130_fd_sc_hd__nand4_1_4 ( .VNB(VNB), .VPWR(VPWR), .A(_2_), .B(p[10]), .C(_31_), .D(_30_), .Y(_32_) );
sky130_fd_sc_hd__nand3_1 sky130_fd_sc_hd__nand3_1_2 ( .VNB(VNB), .VPWR(VPWR), .A(_27_), .B(_29_), .C(_32_), .Y(_33_) );
sky130_fd_sc_hd__o2bb2ai_1 sky130_fd_sc_hd__o2bb2ai_1_1 ( .VNB(VNB), .VPWR(VPWR), .A1_N(_21_), .A2_N(_33_), .B1(_5_), .B2(_20_), .Y(_0__0_) );
sky130_fd_sc_hd__nand2_1 sky130_fd_sc_hd__nand2_1_7 ( .VNB(VNB), .VPWR(VPWR), .A(_19_), .B(_18_), .Y(_34_) );
sky130_fd_sc_hd__nand4_1 sky130_fd_sc_hd__nand4_1_5 ( .VNB(VNB), .VPWR(VPWR), .A(_2_), .B(p[1]), .C(_3_), .D(_4_), .Y(_35_) );
sky130_fd_sc_hd__nor3_1 sky130_fd_sc_hd__nor3_1_2 ( .VNB(VNB), .VPWR(VPWR), .A(_9_), .B(_10_), .C(_12_), .Y(_36_) );
sky130_fd_sc_hd__and2_2 sky130_fd_sc_hd__and2_2_3 ( .VNB(VNB), .VPWR(VPWR), .A(p[12]), .B(p[13]), .X(_37_) );
sky130_fd_sc_hd__nand4_1 sky130_fd_sc_hd__nand4_1_6 ( .VNB(VNB), .VPWR(VPWR), .A(_36_), .B(_7_), .C(_25_), .D(_37_), .Y(_38_) );
sky130_fd_sc_hd__nor2_1 sky130_fd_sc_hd__nor2_1_5 ( .VNB(VNB), .VPWR(VPWR), .A(p[11]), .B(_23_), .Y(_39_) );
sky130_fd_sc_hd__nand3_1 sky130_fd_sc_hd__nand3_1_3 ( .VNB(VNB), .VPWR(VPWR), .A(_21_), .B(_2_), .C(_39_), .Y(_40_) );
sky130_fd_sc_hd__nor3_1 sky130_fd_sc_hd__nor3_1_3 ( .VNB(VNB), .VPWR(VPWR), .A(p[7]), .B(_12_), .C(_6_), .Y(_41_) );
sky130_fd_sc_hd__nand4_1 sky130_fd_sc_hd__nand4_1_7 ( .VNB(VNB), .VPWR(VPWR), .A(_41_), .B(_2_), .C(_3_), .D(_4_), .Y(_42_) );
sky130_fd_sc_hd__o2111ai_1 sky130_fd_sc_hd__o2111ai_1_1 ( .VNB(VNB), .VPWR(VPWR), .A1(_35_), .A2(_34_), .B1(_42_), .C1(_38_), .D1(_40_), .Y(_0__1_) );
sky130_fd_sc_hd__nand2_1 sky130_fd_sc_hd__nand2_1_8 ( .VNB(VNB), .VPWR(VPWR), .A(_36_), .B(_7_), .Y(_43_) );
sky130_fd_sc_hd__nand2_1 sky130_fd_sc_hd__nand2_1_9 ( .VNB(VNB), .VPWR(VPWR), .A(_7_), .B(_18_), .Y(_44_) );
sky130_fd_sc_hd__o21ai_0 sky130_fd_sc_hd__o21ai_0_2 ( .VNB(VNB), .VPWR(VPWR), .A1(_22_), .A2(_37_), .B1(_25_), .Y(_45_) );
sky130_fd_sc_hd__o221ai_1 sky130_fd_sc_hd__o221ai_1_1 ( .VNB(VNB), .VPWR(VPWR), .A1(_5_), .A2(_44_), .B1(_45_), .B2(_43_), .C1(_42_), .Y(_0__2_) );
sky130_fd_sc_hd__nand2_1 sky130_fd_sc_hd__nand2_1_10 ( .VNB(VNB), .VPWR(VPWR), .A(_39_), .B(_2_), .Y(_46_) );
sky130_fd_sc_hd__a41oi_1 sky130_fd_sc_hd__a41oi_1_1 ( .VNB(VNB), .VPWR(VPWR), .A1(_29_), .A2(_45_), .A3(_46_), .A4(_5_), .B1(_43_), .Y(_0__3_) );
sky130_fd_sc_hd__clkinv_1 sky130_fd_sc_hd__clkinv_1_7 ( .VNB(VNB), .VPWR(VPWR), .A(rst), .Y(_1_) );
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_3 ( .VNB(VNB), .VPWR(VPWR), .A(_47__0_), .X(b[0]) );
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_4 ( .VNB(VNB), .VPWR(VPWR), .A(_47__1_), .X(b[1]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_1 ( .VNB(VNB), .VPWR(VPWR), .DIODE(clk) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_2 ( .VNB(VNB), .VPWR(VPWR), .DIODE(rst) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_3 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[0]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_4 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[1]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_5 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[2]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_6 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[3]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_7 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[4]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_8 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[5]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_9 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[6]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_10 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[7]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_11 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[8]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_12 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[9]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_13 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[10]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_14 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[11]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_15 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[12]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_16 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[13]) );
sky130_fd_sc_hd__diode_2 sky130_fd_sc_hd__diode_2_17 ( .VNB(VNB), .VPWR(VPWR), .DIODE(p[14]) );
endmodule
