magic
tech sky130A
magscale 1 2
timestamp 1704877912
<< error_p >>
rect -31 231 31 237
rect -31 197 -19 231
rect -31 191 31 197
rect -31 -197 31 -191
rect -31 -231 -19 -197
rect -31 -237 31 -231
<< nwell >>
rect -231 -369 231 369
<< pmos >>
rect -35 -150 35 150
<< pdiff >>
rect -93 138 -35 150
rect -93 -138 -81 138
rect -47 -138 -35 138
rect -93 -150 -35 -138
rect 35 138 93 150
rect 35 -138 47 138
rect 81 -138 93 138
rect 35 -150 93 -138
<< pdiffc >>
rect -81 -138 -47 138
rect 47 -138 81 138
<< nsubdiff >>
rect -195 299 -99 333
rect 99 299 195 333
rect -195 237 -161 299
rect 161 237 195 299
rect -195 -299 -161 -237
rect 161 -299 195 -237
rect -195 -333 -99 -299
rect 99 -333 195 -299
<< nsubdiffcont >>
rect -99 299 99 333
rect -195 -237 -161 237
rect 161 -237 195 237
rect -99 -333 99 -299
<< poly >>
rect -35 231 35 247
rect -35 197 -19 231
rect 19 197 35 231
rect -35 150 35 197
rect -35 -197 35 -150
rect -35 -231 -19 -197
rect 19 -231 35 -197
rect -35 -247 35 -231
<< polycont >>
rect -19 197 19 231
rect -19 -231 19 -197
<< locali >>
rect -195 299 -99 333
rect 99 299 195 333
rect -195 237 -161 299
rect 161 237 195 299
rect -35 197 -19 231
rect 19 197 35 231
rect -81 138 -47 154
rect -81 -154 -47 -138
rect 47 138 81 154
rect 47 -154 81 -138
rect -35 -231 -19 -197
rect 19 -231 35 -197
rect -195 -299 -161 -237
rect 161 -299 195 -237
rect -195 -333 -99 -299
rect 99 -333 195 -299
<< viali >>
rect -19 197 19 231
rect -81 -138 -47 138
rect 47 -138 81 138
rect -19 -231 19 -197
<< metal1 >>
rect -31 231 31 237
rect -31 197 -19 231
rect 19 197 31 231
rect -31 191 31 197
rect -87 138 -41 150
rect -87 -138 -81 138
rect -47 -138 -41 138
rect -87 -150 -41 -138
rect 41 138 87 150
rect 41 -138 47 138
rect 81 -138 87 138
rect 41 -150 87 -138
rect -31 -197 31 -191
rect -31 -231 -19 -197
rect 19 -231 31 -197
rect -31 -237 31 -231
<< properties >>
string FIXED_BBOX -178 -316 178 316
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
