magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_s >>
rect 298 999 333 1016
rect 299 998 333 999
rect 721 1009 756 1016
rect 721 998 755 1009
rect 299 962 369 998
rect 129 931 187 937
rect 129 897 141 931
rect 316 928 387 962
rect 129 891 187 897
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 928
rect 498 860 556 866
rect 498 826 510 860
rect 498 820 556 826
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 316 547 369 583
rect 685 530 755 998
rect 867 941 925 947
rect 867 907 879 941
rect 867 901 925 907
rect 1037 874 1071 928
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 685 494 738 530
rect 1056 477 1071 874
rect 1090 840 1125 874
rect 1405 840 1440 874
rect 1090 477 1124 840
rect 1406 821 1440 840
rect 1236 772 1294 778
rect 1236 738 1248 772
rect 1236 732 1294 738
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1090 443 1105 477
rect 1425 424 1440 821
rect 1459 787 1494 821
rect 1774 787 1809 804
rect 1459 424 1493 787
rect 1775 786 1809 787
rect 1775 750 1845 786
rect 1605 719 1663 725
rect 1605 685 1617 719
rect 1792 716 1863 750
rect 1605 679 1663 685
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1459 390 1474 424
rect 1792 371 1862 716
rect 1974 648 2032 654
rect 1974 614 1986 648
rect 1974 608 2032 614
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1792 335 1845 371
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_M479BZ  XM1
timestamp 1703732895
transform 1 0 158 0 1 808
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 1703732895
transform 1 0 896 0 1 760
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_L7T3GD  XM3
timestamp 1703732895
transform 1 0 527 0 1 746
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_M479BZ  XM7
timestamp 1703732895
transform 1 0 1265 0 1 649
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_M479BZ  XM9
timestamp 1703732895
transform 1 0 1634 0 1 596
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_L7T3GD  XM10
timestamp 1703732895
transform 1 0 2003 0 1 534
box -211 -252 211 252
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
