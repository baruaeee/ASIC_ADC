magic
tech sky130A
magscale 1 2
timestamp 1704322866
<< error_p >>
rect -29 216 29 222
rect -29 182 -17 216
rect -29 176 29 182
rect -29 -182 29 -176
rect -29 -216 -17 -182
rect -29 -222 29 -216
<< nwell >>
rect -211 -354 211 354
<< pmos >>
rect -15 -135 15 135
<< pdiff >>
rect -73 123 -15 135
rect -73 -123 -61 123
rect -27 -123 -15 123
rect -73 -135 -15 -123
rect 15 123 73 135
rect 15 -123 27 123
rect 61 -123 73 123
rect 15 -135 73 -123
<< pdiffc >>
rect -61 -123 -27 123
rect 27 -123 61 123
<< nsubdiff >>
rect -175 284 -79 318
rect 79 284 175 318
rect -175 222 -141 284
rect 141 222 175 284
rect -175 -284 -141 -222
rect 141 -284 175 -222
rect -175 -318 -79 -284
rect 79 -318 175 -284
<< nsubdiffcont >>
rect -79 284 79 318
rect -175 -222 -141 222
rect 141 -222 175 222
rect -79 -318 79 -284
<< poly >>
rect -33 216 33 232
rect -33 182 -17 216
rect 17 182 33 216
rect -33 166 33 182
rect -15 135 15 166
rect -15 -166 15 -135
rect -33 -182 33 -166
rect -33 -216 -17 -182
rect 17 -216 33 -182
rect -33 -232 33 -216
<< polycont >>
rect -17 182 17 216
rect -17 -216 17 -182
<< locali >>
rect -175 284 -79 318
rect 79 284 175 318
rect -175 222 -141 284
rect 141 222 175 284
rect -33 182 -17 216
rect 17 182 33 216
rect -61 123 -27 139
rect -61 -139 -27 -123
rect 27 123 61 139
rect 27 -139 61 -123
rect -33 -216 -17 -182
rect 17 -216 33 -182
rect -175 -284 -141 -222
rect 141 -284 175 -222
rect -175 -318 -79 -284
rect 79 -318 175 -284
<< viali >>
rect -17 182 17 216
rect -61 -123 -27 123
rect 27 -123 61 123
rect -17 -216 17 -182
<< metal1 >>
rect -29 216 29 222
rect -29 182 -17 216
rect 17 182 29 216
rect -29 176 29 182
rect -67 123 -21 135
rect -67 -123 -61 123
rect -27 -123 -21 123
rect -67 -135 -21 -123
rect 21 123 67 135
rect 21 -123 27 123
rect 61 -123 67 123
rect 21 -135 67 -123
rect -29 -182 29 -176
rect -29 -216 -17 -182
rect 17 -216 29 -182
rect -29 -222 29 -216
<< properties >>
string FIXED_BBOX -158 -301 158 301
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.349 l 0.151 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
