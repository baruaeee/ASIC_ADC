VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO oaTaper STRING ;
  MACRO CatenaDesignType STRING ;
  MACRO lastSavedExtractCounter INTEGER ;
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_WIDTH STRING ;
END PROPERTYDEFINITIONS

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER dnwell
  TYPE MASTERSLICE ;
END dnwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
  PROPERTY LEF58_SPACING "SPACING 1.27 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.84 ;" ;
END nwell

LAYER diff
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
  PROPERTY LEF58_SPACING "SPACING 0.27 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.15 ;" ;
END diff

LAYER tap
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
  PROPERTY LEF58_SPACING "SPACING 0.27 ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.15 ;" ;
END tap

LAYER nsdm
  TYPE IMPLANT ;
  WIDTH 0.38 ;
  SPACING 0.38 ;
  AREA 0.265 ;
END nsdm

LAYER psdm
  TYPE IMPLANT ;
  WIDTH 0.38 ;
  SPACING 0.38 ;
  AREA 0.255 ;
END psdm

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER npc
  TYPE CUT ;
  SPACING 0.27 ;
  WIDTH 0.27 ;
  ANTENNAMODEL OXIDE1 ;
END npc

LAYER licon1
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE MEOL ;" ;
END licon1

LAYER li1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.17 ;
  AREA 0.056 ;
  SPACING 0.17 ;
  SPACING 0.17 SAMENET ;
  RESISTANCE RPERSQ 12.2 ;
  CAPACITANCE CPERSQDIST 3.69e-05 ;
  THICKNESS 0.1 ;
  EDGECAPACITANCE 3.26e-06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 75 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 75 ) ( 0.0125 75 ) ( 0.0225 85.125 ) ( 22.5 10200 ) ) ;
END li1

LAYER mcon
  TYPE CUT ;
  SPACING 0.19 ;
  WIDTH 0.17 ;
  ENCLOSURE BELOW 0 0 ;
  ENCLOSURE ABOVE 0.03 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 3 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 3 ) ( 0.0125 3 ) ( 0.0225 3.405 ) ( 22.5 408 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.36 ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.28 0.28 ;
  WIDTH 0.14 ;
  OFFSET 0.14 0.14 ;
  AREA 0.083 ;
  SPACING 0.14 ;
  SPACING 0.28 RANGE 3.005 10000 ;
  SPACING 0.14 SAMENET ;
  SPACING 0.28 RANGE 3.005 10000 INFLUENCE 0.28 ;
  MAXWIDTH 4 ;
  MINENCLOSEDAREA 0.14 ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 2.58e-05 ;
  THICKNESS 0.35 ;
  EDGECAPACITANCE 1.79e-06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
  ACCURRENTDENSITY RMS 6.1 ;
  DCCURRENTDENSITY AVERAGE 2.8 ;
END met1

LAYER via
  TYPE CUT ;
  SPACING 0.17 ;
  WIDTH 0.15 ;
  ENCLOSURE BELOW 0.055 0.085 ;
  ENCLOSURE ABOVE 0.055 0.085 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 6 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.29 ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.28 0.28 ;
  WIDTH 0.14 ;
  OFFSET 0.14 0.14 ;
  AREA 0.0676 ;
  SPACING 0.14 ;
  SPACING 0.28 RANGE 3.005 10000 ;
  SPACING 0.14 SAMENET ;
  SPACING 0.28 RANGE 3.005 10000 INFLUENCE 0.28 ;
  MAXWIDTH 4 ;
  MINENCLOSEDAREA 0.14 ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 1.75e-05 ;
  THICKNESS 0.35 ;
  EDGECAPACITANCE 1.22e-06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
  ACCURRENTDENSITY RMS 6.1 ;
  DCCURRENTDENSITY AVERAGE 2.8 ;
END met2

LAYER via2
  TYPE CUT ;
  SPACING 0.2 ;
  WIDTH 0.2 ;
  ENCLOSURE BELOW 0.04 0.085 ;
  ENCLOSURE ABOVE 0.065 0.065 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 6 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.6 0.6 ;
  WIDTH 0.3 ;
  OFFSET 0.3 0.3 ;
  AREA 0.24 ;
  SPACING 0.3 ;
  SPACING 0.4 RANGE 3.005 10000 ;
  SPACING 0.3 SAMENET ;
  SPACING 0.4 RANGE 3.005 10000 INFLUENCE 0.4 ;
  MAXWIDTH 4 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.047 ;
  CAPACITANCE CPERSQDIST 1.26e-05 ;
  THICKNESS 0.8 ;
  EDGECAPACITANCE 1.86e-06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
  ACCURRENTDENSITY RMS 14.9 ;
  DCCURRENTDENSITY AVERAGE 6.8 ;
END met3

LAYER via3
  TYPE CUT ;
  SPACING 0.2 ;
  WIDTH 0.2 ;
  ENCLOSURE BELOW 0.06 0.09 ;
  ENCLOSURE ABOVE 0.065 0.065 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 6 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.6 0.6 ;
  WIDTH 0.3 ;
  OFFSET 0.3 0.3 ;
  AREA 0.24 ;
  SPACING 0.3 ;
  SPACING 0.4 RANGE 3.005 10000 ;
  SPACING 0.3 SAMENET ;
  SPACING 0.4 RANGE 3.005 10000 INFLUENCE 0.4 ;
  MAXWIDTH 10 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.047 ;
  CAPACITANCE CPERSQDIST 8.67e-06 ;
  THICKNESS 0.8 ;
  EDGECAPACITANCE 1.29e-06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
  ACCURRENTDENSITY RMS 14.9 ;
  DCCURRENTDENSITY AVERAGE 6.8 ;
END met4

LAYER via4
  TYPE CUT ;
  SPACING 0.8 ;
  WIDTH 0.8 ;
  ENCLOSURE BELOW 0.19 0.19 ;
  ENCLOSURE ABOVE 0.31 0.31 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 6 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 2.49 ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.2 3.2 ;
  WIDTH 1.6 ;
  OFFSET 1.6 1.6 ;
  AREA 4 ;
  SPACING 1.6 ;
  SPACING 1.6 SAMENET ;
  RESISTANCE RPERSQ 0.0285 ;
  CAPACITANCE CPERSQDIST 6.48e-06 ;
  THICKNESS 1.2 ;
  EDGECAPACITANCE 4.96e-06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
  ACCURRENTDENSITY RMS 22.34 ;
  DCCURRENTDENSITY AVERAGE 10.17 ;
END met5

LAYER rdl
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 10 ;
  SPACING 10 ;
  RESISTANCE RPERSQ 0.005 ;
  CAPACITANCE CPERSQDIST 2.66e-06 ;
  THICKNESS 2 ;
  EDGECAPACITANCE 6.2e-06 ;
  ANTENNAMODEL OXIDE1 ;
END rdl

VIARULE M4M5_C GENERATE DEFAULT
  LAYER met5 ;
    ENCLOSURE 0.31 0.31 ;
  LAYER met4 ;
    ENCLOSURE 0.19 0.19 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.6 BY 1.6 ;
    RESISTANCE 0.380000 ;
END M4M5_C

VIARULE M3M4_C GENERATE DEFAULT
  LAYER met4 ;
    ENCLOSURE 0.065 0.065 ;
  LAYER met3 ;
    ENCLOSURE 0.06 0.09 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.4 BY 0.4 ;
    RESISTANCE 3.410000 ;
END M3M4_C

VIARULE M2M3_C GENERATE DEFAULT
  LAYER met3 ;
    ENCLOSURE 0.065 0.065 ;
  LAYER met2 ;
    ENCLOSURE 0.04 0.085 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.4 BY 0.4 ;
    RESISTANCE 3.410000 ;
END M2M3_C

VIARULE M1M2_C GENERATE DEFAULT
  LAYER met2 ;
    ENCLOSURE 0.055 0.085 ;
  LAYER met1 ;
    ENCLOSURE 0.055 0.085 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
    SPACING 0.32 BY 0.32 ;
    RESISTANCE 4.500000 ;
END M1M2_C

VIARULE L1M1_C GENERATE DEFAULT
  LAYER met1 ;
    ENCLOSURE 0.03 0.06 ;
  LAYER li1 ;
    ENCLOSURE 0 0.08 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
    SPACING 0.36 BY 0.36 ;
    RESISTANCE 9.300000 ;
END L1M1_C

VIA PYL1CON_C_0
  VIARULE PYL1CON_C ;
  CUTSIZE 0.37 0.37 ;
  LAYERS poly npc licon1 ;
  CUTSPACING 0.27 0.27 ;
  ENCLOSURE -0.05 -0.02 -0.1 -0.1 ;
  ROWCOL 1 1 ;
END PYL1CON_C_0

VIA PYL1CON_C_1
  VIARULE PYL1CON_C ;
  CUTSIZE 0.37 0.37 ;
  LAYERS poly npc licon1 ;
  CUTSPACING 0.27 0.27 ;
  ENCLOSURE -0.05 -0.02 -0.1 -0.1 ;
  ROWCOL 1 1 ;
END PYL1CON_C_1

VIA L1M1_C_2
  VIARULE L1M1_C ;
  CUTSIZE 0.17 0.17 ;
  LAYERS li1 mcon met1 ;
  CUTSPACING 0.19 0.19 ;
  ENCLOSURE 0 0.08 0.03 0.06 ;
  ROWCOL 1 1 ;
END L1M1_C_2

VIA L1M1_C_3
  VIARULE L1M1_C ;
  CUTSIZE 0.17 0.17 ;
  LAYERS li1 mcon met1 ;
  CUTSPACING 0.19 0.19 ;
  ENCLOSURE 0.08 0 0.03 0.06 ;
  ROWCOL 1 1 ;
END L1M1_C_3

VIA L1M1_C_4
  VIARULE L1M1_C ;
  CUTSIZE 0.17 0.17 ;
  LAYERS li1 mcon met1 ;
  CUTSPACING 0.19 0.19 ;
  ENCLOSURE 0 0.08 0.03 0.06 ;
  ROWCOL 2 1 ;
END L1M1_C_4

VIA L1M1_C_5
  VIARULE L1M1_C ;
  CUTSIZE 0.17 0.17 ;
  LAYERS li1 mcon met1 ;
  CUTSPACING 0.19 0.19 ;
  ENCLOSURE 0 0.08 0.03 0.06 ;
  ROWCOL 1 1 ;
END L1M1_C_5

MACRO inv01f
  ORIGIN 0 0 ;
  FOREIGN inv01f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.43 1.39 0.78 1.64 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 1.03 -0.17 1.38 0.08 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 1.03 3.835 1.38 4.085 ;
    END
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.25 0.96 1.5 1.31 ;
    END
  END Y
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY lastSavedExtractCounter 5684 ;
END inv01f

END LIBRARY
