magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< nwell >>
rect -240 -261 240 261
<< pmos >>
rect -44 -42 44 42
<< pdiff >>
rect -102 30 -44 42
rect -102 -30 -90 30
rect -56 -30 -44 30
rect -102 -42 -44 -30
rect 44 30 102 42
rect 44 -30 56 30
rect 90 -30 102 30
rect 44 -42 102 -30
<< pdiffc >>
rect -90 -30 -56 30
rect 56 -30 90 30
<< nsubdiff >>
rect -204 191 -108 225
rect 108 191 204 225
rect -204 129 -170 191
rect 170 129 204 191
rect -204 -191 -170 -129
rect 170 -191 204 -129
rect -204 -225 -108 -191
rect 108 -225 204 -191
<< nsubdiffcont >>
rect -108 191 108 225
rect -204 -129 -170 129
rect 170 -129 204 129
rect -108 -225 108 -191
<< poly >>
rect -44 123 44 139
rect -44 89 -28 123
rect 28 89 44 123
rect -44 42 44 89
rect -44 -89 44 -42
rect -44 -123 -28 -89
rect 28 -123 44 -89
rect -44 -139 44 -123
<< polycont >>
rect -28 89 28 123
rect -28 -123 28 -89
<< locali >>
rect -204 191 -108 225
rect 108 191 204 225
rect -204 129 -170 191
rect 170 129 204 191
rect -44 89 -28 123
rect 28 89 44 123
rect -90 30 -56 46
rect -90 -46 -56 -30
rect 56 30 90 46
rect 56 -46 90 -30
rect -44 -123 -28 -89
rect 28 -123 44 -89
rect -204 -191 -170 -129
rect 170 -191 204 -129
rect -204 -225 -108 -191
rect 108 -225 204 -191
<< viali >>
rect -28 89 28 123
rect -90 -30 -56 30
rect 56 -30 90 30
rect -28 -123 28 -89
<< metal1 >>
rect -40 123 40 129
rect -40 89 -28 123
rect 28 89 40 123
rect -40 83 40 89
rect -96 30 -50 42
rect -96 -30 -90 30
rect -56 -30 -50 30
rect -96 -42 -50 -30
rect 50 30 96 42
rect 50 -30 56 30
rect 90 -30 96 30
rect 50 -42 96 -30
rect -40 -89 40 -83
rect -40 -123 -28 -89
rect 28 -123 40 -89
rect -40 -129 40 -123
<< properties >>
string FIXED_BBOX -187 -208 187 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.436 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
