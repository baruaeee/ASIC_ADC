magic
tech sky130A
magscale 1 2
timestamp 1708346635
<< checkpaint >>
rect -1313 2318 2299 2427
rect -1313 -713 2668 2318
rect -1260 -766 2668 -713
rect -1260 -2460 1460 -766
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_MWHFPY  XM0
timestamp 0
transform 1 0 1197 0 1 776
box -211 -282 211 282
use sky130_fd_pr__nfet_01v8_DPSGWY  XM1
timestamp 0
transform 1 0 493 0 1 857
box -546 -310 546 310
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vpamp
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
