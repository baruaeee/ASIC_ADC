magic
tech sky130A
magscale 1 2
timestamp 1706402911
<< psubdiff >>
rect 447 686 891 720
rect 1416 254 1422 261
rect 1416 195 1450 254
<< locali >>
rect 706 1268 786 1304
rect 455 686 863 720
rect 1416 254 1422 259
rect 1416 233 1450 254
<< viali >>
rect 672 1268 706 1304
rect 863 686 897 720
rect 1416 199 1450 233
<< metal1 >>
rect 556 1317 656 1330
rect 556 1312 714 1317
rect 556 1304 715 1312
rect 556 1268 672 1304
rect 706 1268 715 1304
rect 556 1260 715 1268
rect 556 1256 714 1260
rect 556 1230 656 1256
rect 571 1166 615 1230
rect 511 1114 517 1166
rect 569 1122 615 1166
rect 896 1162 954 1222
rect 569 1114 575 1122
rect 953 1105 987 1109
rect 647 1032 653 1084
rect 705 1076 711 1084
rect 705 1042 898 1076
rect 953 1071 1365 1105
rect 705 1032 711 1042
rect 953 1009 987 1071
rect 1331 1040 1365 1071
rect 394 948 494 984
rect 394 914 947 948
rect 1300 940 1400 1040
rect 394 884 494 914
rect 510 784 517 836
rect 569 784 575 836
rect 510 535 542 784
rect 607 617 641 914
rect 770 800 822 806
rect 770 742 822 748
rect 779 728 822 742
rect 857 728 903 732
rect 779 720 903 728
rect 779 686 863 720
rect 897 719 903 720
rect 897 686 909 719
rect 779 685 909 686
rect 857 674 903 685
rect 607 583 1029 617
rect 1331 535 1365 940
rect 510 514 579 535
rect 511 501 579 514
rect 512 359 579 501
rect 1303 534 1365 535
rect 512 358 546 359
rect 1303 357 1366 534
rect 1457 239 1494 254
rect 1404 236 1494 239
rect 1390 233 1494 236
rect 1390 199 1416 233
rect 1450 199 1494 233
rect 1390 172 1494 199
rect 1390 136 1490 172
<< via1 >>
rect 517 1114 569 1166
rect 653 1032 705 1084
rect 517 784 569 836
rect 770 748 822 800
<< metal2 >>
rect 517 1166 569 1172
rect 517 1108 569 1114
rect 526 842 560 1108
rect 653 1084 705 1090
rect 653 1026 705 1032
rect 517 836 569 842
rect 517 778 569 784
rect 662 791 696 1026
rect 764 791 770 800
rect 662 757 770 791
rect 764 748 770 757
rect 822 748 828 800
use sky130_fd_pr__pfet_01v8_MWHFPY  XM0
timestamp 1706203507
transform 1 0 925 0 1 1058
box -211 -282 211 282
use sky130_fd_pr__nfet_01v8_DPSGWY  XM1
timestamp 1706134018
transform 1 0 940 0 1 446
box -546 -310 546 310
<< labels >>
flabel metal1 556 1230 656 1330 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 1390 136 1490 236 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 1300 940 1400 1040 0 FreeSans 256 0 0 0 Vpamp
port 2 nsew
flabel metal1 394 884 494 984 0 FreeSans 256 0 0 0 Vin
port 1 nsew
<< end >>
