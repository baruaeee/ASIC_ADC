magic
tech sky130A
magscale 1 2
timestamp 1704305861
<< error_p >>
rect -29 531 29 537
rect -29 497 -17 531
rect -29 491 29 497
rect -29 -497 29 -491
rect -29 -531 -17 -497
rect -29 -537 29 -531
<< nwell >>
rect -211 -669 211 669
<< pmos >>
rect -15 -450 15 450
<< pdiff >>
rect -73 438 -15 450
rect -73 -438 -61 438
rect -27 -438 -15 438
rect -73 -450 -15 -438
rect 15 438 73 450
rect 15 -438 27 438
rect 61 -438 73 438
rect 15 -450 73 -438
<< pdiffc >>
rect -61 -438 -27 438
rect 27 -438 61 438
<< nsubdiff >>
rect -175 599 -79 633
rect 79 599 175 633
rect -175 537 -141 599
rect 141 537 175 599
rect -175 -599 -141 -537
rect 141 -599 175 -537
rect -175 -633 -79 -599
rect 79 -633 175 -599
<< nsubdiffcont >>
rect -79 599 79 633
rect -175 -537 -141 537
rect 141 -537 175 537
rect -79 -633 79 -599
<< poly >>
rect -33 531 33 547
rect -33 497 -17 531
rect 17 497 33 531
rect -33 481 33 497
rect -15 450 15 481
rect -15 -481 15 -450
rect -33 -497 33 -481
rect -33 -531 -17 -497
rect 17 -531 33 -497
rect -33 -547 33 -531
<< polycont >>
rect -17 497 17 531
rect -17 -531 17 -497
<< locali >>
rect -175 599 -79 633
rect 79 599 175 633
rect -175 537 -141 599
rect 141 537 175 599
rect -33 497 -17 531
rect 17 497 33 531
rect -61 438 -27 454
rect -61 -454 -27 -438
rect 27 438 61 454
rect 27 -454 61 -438
rect -33 -531 -17 -497
rect 17 -531 33 -497
rect -175 -599 -141 -537
rect 141 -599 175 -537
rect -175 -633 -79 -599
rect 79 -633 175 -599
<< viali >>
rect -17 497 17 531
rect -61 -438 -27 438
rect 27 -438 61 438
rect -17 -531 17 -497
<< metal1 >>
rect -29 531 29 537
rect -29 497 -17 531
rect 17 497 29 531
rect -29 491 29 497
rect -67 438 -21 450
rect -67 -438 -61 438
rect -27 -438 -21 438
rect -67 -450 -21 -438
rect 21 438 67 450
rect 21 -438 27 438
rect 61 -438 67 438
rect 21 -450 67 -438
rect -29 -497 29 -491
rect -29 -531 -17 -497
rect 17 -531 29 -497
rect -29 -537 29 -531
<< properties >>
string FIXED_BBOX -158 -616 158 616
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
