* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : inv09f                                       *
* Netlisted  : Sun Dec  1 16:07:56 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733065665430                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733065665430 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.1e-06 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733065665430

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733065665431                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733065665431 1 2 3
** N=9 EP=3 FDC=2
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.7e-07 $X=0 $Y=0 $dt=8
M1 1 3 2 1 pfet_01v8 L=1.5e-07 W=7.7e-07 $X=430 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733065665431

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv09f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv09f A VDD VSS Y
** N=9 EP=4 FDC=3
X2 VSS Y A nfet_01v8_CDNS_733065665430 $T=905 695 0 90 $X=335 $Y=290
X3 VDD Y A pfet_01v8_CDNS_733065665431 $T=400 2840 0 0 $X=-45 $Y=2660
.ends inv09f
