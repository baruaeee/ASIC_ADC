* NGSPICE file created from th05.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_Q7AWK3 a_n180_n340# a_20_n200# a_n78_n200# a_n33_n288#
X0 a_20_n200# a_n33_n288# a_n78_n200# a_n180_n340# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
C0 a_n78_n200# a_n33_n288# 0.024f
C1 a_20_n200# a_n78_n200# 0.288f
C2 a_20_n200# a_n33_n288# 0.024f
C3 a_20_n200# a_n180_n340# 0.202f
C4 a_n78_n200# a_n180_n340# 0.237f
C5 a_n33_n288# a_n180_n340# 0.325f
.ends

.subckt sky130_fd_pr__pfet_01v8_EXJYQP w_n359_n261# a_n163_n139# a_n221_n42# a_163_n42#
+ VSUBS
X0 a_163_n42# a_n163_n139# a_n221_n42# w_n359_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.63
C0 a_n163_n139# w_n359_n261# 0.413f
C1 a_n221_n42# a_n163_n139# 0.0182f
C2 a_n221_n42# w_n359_n261# 0.0179f
C3 a_163_n42# a_n163_n139# 0.0182f
C4 a_163_n42# w_n359_n261# 0.0408f
C5 a_163_n42# a_n221_n42# 0.0161f
C6 a_163_n42# VSUBS 0.041f
C7 a_n221_n42# VSUBS 0.056f
C8 a_n163_n139# VSUBS 0.584f
C9 w_n359_n261# VSUBS 1.24f
.ends

.subckt sky130_fd_pr__pfet_01v8_HJHF6N a_n170_n50# w_n308_n269# a_n112_n147# a_112_n50#
+ VSUBS
X0 a_112_n50# a_n112_n147# a_n170_n50# w_n308_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1.12
C0 a_n112_n147# w_n308_n269# 0.378f
C1 a_n170_n50# a_n112_n147# 0.0172f
C2 a_n170_n50# w_n308_n269# 0.0232f
C3 a_112_n50# a_n112_n147# 0.0172f
C4 a_112_n50# w_n308_n269# 0.0232f
C5 a_112_n50# a_n170_n50# 0.0259f
C6 a_112_n50# VSUBS 0.0577f
C7 a_n170_n50# VSUBS 0.0577f
C8 a_n112_n147# VSUBS 0.389f
C9 w_n308_n269# VSUBS 1.14f
.ends

.subckt sky130_fd_pr__nfet_01v8_N39H2X a_n76_n100# a_n33_n188# a_18_n100# a_144_n240#
X0 a_18_n100# a_n33_n188# a_n76_n100# a_144_n240# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.18
C0 a_n76_n100# a_n33_n188# 0.0205f
C1 a_18_n100# a_n76_n100# 0.152f
C2 a_18_n100# a_n33_n188# 0.0205f
C3 a_18_n100# a_144_n240# 0.133f
C4 a_n76_n100# a_144_n240# 0.115f
C5 a_n33_n188# a_144_n240# 0.32f
.ends

.subckt th05 Vp V05 Vin Vn
XXM0 Vn m1_752_n794# Vn Vin sky130_fd_pr__nfet_01v8_Q7AWK3
XXM1 Vp Vin m1_752_n794# Vp Vn sky130_fd_pr__pfet_01v8_EXJYQP
XXM2 Vp Vp m1_752_n794# V05 Vn sky130_fd_pr__pfet_01v8_HJHF6N
XXM3 Vn m1_752_n794# V05 Vn sky130_fd_pr__nfet_01v8_N39H2X
C0 m1_752_n794# Vin 0.2f
C1 V05 m1_752_n794# 0.0855f
C2 Vn Vp 0.0115f
C3 Vn Vin 0.041f
C4 V05 Vn 0.0364f
C5 Vp Vin 0.139f
C6 V05 Vp 0.0548f
C7 V05 Vin 0.00406f
C8 Vn m1_752_n794# 0.136f
C9 Vp m1_752_n794# 0.198f
C10 Vin 0 0.905f
C11 Vp 0 2.28f
C12 V05 0 0.314f
C13 m1_752_n794# 0 0.788f
C14 Vn 0 0.547f
.ends

