magic
tech sky130A
magscale 1 2
timestamp 1706224144
<< nwell >>
rect -359 -261 359 261
<< pmos >>
rect -163 -42 163 42
<< pdiff >>
rect -221 30 -163 42
rect -221 -30 -209 30
rect -175 -30 -163 30
rect -221 -42 -163 -30
rect 163 30 221 42
rect 163 -30 175 30
rect 209 -30 221 30
rect 163 -42 221 -30
<< pdiffc >>
rect -209 -30 -175 30
rect 175 -30 209 30
<< nsubdiff >>
rect 289 129 323 191
rect 289 -191 323 -129
<< nsubdiffcont >>
rect 289 -129 323 129
<< poly >>
rect -163 123 163 139
rect -163 89 -147 123
rect 147 89 163 123
rect -163 42 163 89
rect -163 -89 163 -42
rect -163 -123 -147 -89
rect 147 -123 163 -89
rect -163 -139 163 -123
<< polycont >>
rect -147 89 147 123
rect -147 -123 147 -89
<< locali >>
rect 289 129 323 191
rect -163 89 -147 123
rect 147 89 163 123
rect -209 30 -175 46
rect -209 -46 -175 -30
rect 175 30 209 46
rect 175 -46 209 -30
rect -163 -123 -147 -89
rect 147 -123 163 -89
rect 289 -191 323 -129
<< viali >>
rect -147 89 147 123
rect -209 -30 -175 30
rect 175 -30 209 30
rect -147 -123 147 -89
<< metal1 >>
rect -159 123 159 129
rect -159 89 -147 123
rect 147 89 159 123
rect -159 83 159 89
rect -215 30 -169 42
rect -215 -30 -209 30
rect -175 -30 -169 30
rect -215 -42 -169 -30
rect 169 30 215 42
rect 169 -30 175 30
rect 209 -30 215 30
rect 169 -42 215 -30
rect -159 -89 159 -83
rect -159 -123 -147 -89
rect 147 -123 159 -89
rect -159 -129 159 -123
<< properties >>
string FIXED_BBOX -306 -208 306 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 1.633 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
