** sch_path: /home/exotic/Desktop/ASIC_ADC/xschem/Vth_sch/test_ngspice/test_script1.sch
**.subckt test_script1 Vout
*.opin Vout
R1 VDD Vout 1k m=1
R2 Vout GND 1k m=1
V1 VDD GND 3
**** begin user architecture code


*.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.save all
.op

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
