* NGSPICE file created from preamp.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_4N47A3 w_n231_n369# a_n93_n150# a_35_n150# a_n35_n247#
+ VSUBS
X0 a_35_n150# a_n35_n247# a_n93_n150# w_n231_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.35
C0 a_35_n150# a_n35_n247# 0.0165f
C1 a_n93_n150# a_n35_n247# 0.0165f
C2 a_n93_n150# a_35_n150# 0.166f
C3 a_n35_n247# w_n231_n369# 0.233f
C4 a_35_n150# w_n231_n369# 0.116f
C5 a_n93_n150# w_n231_n369# 0.116f
C6 a_35_n150# VSUBS 0.0757f
C7 a_n93_n150# VSUBS 0.0757f
C8 a_n35_n247# VSUBS 0.141f
C9 w_n231_n369# VSUBS 1.52f
.ends

.subckt sky130_fd_pr__nfet_01v8_48YMBA a_n518_n42# a_460_n42# a_n620_n216# a_n460_n130#
X0 a_460_n42# a_n460_n130# a_n518_n42# a_n620_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=4.6
C0 a_460_n42# a_n518_n42# 0.00624f
C1 a_n518_n42# a_n460_n130# 0.0236f
C2 a_460_n42# a_n460_n130# 0.0236f
C3 a_460_n42# a_n620_n216# 0.0868f
C4 a_n518_n42# a_n620_n216# 0.0868f
C5 a_n460_n130# a_n620_n216# 2.69f
.ends

.subckt preamp Vp Vin Vpamp Vn
XXM0 Vpamp Vn Vpamp Vin Vpamp sky130_fd_pr__pfet_01v8_4N47A3
XXM1 Vp Vpamp Vpamp Vin sky130_fd_pr__nfet_01v8_48YMBA
C0 Vn Vpamp 0.213f
C1 Vpamp Vp 0.0775f
C2 Vin Vpamp 0.488f
C3 Vn Vp 0.0228f
C4 Vin Vn 0.0147f
C5 Vin Vp 0.233f
C6 Vpamp 0 1.57f
C7 Vp 0 0.377f
C8 Vin 0 2.67f
C9 Vn 0 0.247f
.ends

