.subckt th01 Vp Vin Vout Vn
XM1 Vn Vn net2 net2 sky130_fd_pr__pfet_01v8 L=12 W=0.42 nf=1
XM2 Vp Vp net1 net1 sky130_fd_pr__nfet_01v8 L=12 W=0.36 nf=1
XM7 Vout net3 Vp Vp sky130_fd_pr__pfet_01v8 L=0.15000 W=0.42 nf=1
XM10 Vout net3 Vn Vn sky130_fd_pr__nfet_01v8 L=4.5 W=0.42 nf=1
XM3 net3 net4 Vp Vp sky130_fd_pr__pfet_01v8 L=5.00 W=0.42 nf=1
XM4 net3 net4 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15000 W=0.36 nf=1
XM5 net2 Vin net4 net4 sky130_fd_pr__pfet_01v8 L=12 W=0.42 nf=1
XM6 net1 Vin net4 net4 sky130_fd_pr__nfet_01v8 L=12 W=0.36 nf=1
.ends th01


.subckt th02 Vp Vout Vin Vn
XM7 Vout net1 Vp Vp sky130_fd_pr__pfet_01v8 L=0.150 W=24.000 nf=1
XM1 net1 Vin net2 net2 sky130_fd_pr__pfet_01v8 L=23.6000 W=0.42 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=23.6000 nf=1
XM2 Vp Vp net2 net2 sky130_fd_pr__nfet_01v8 L=23.55 W=0.36 nf=1
XM4 Vout net1 net3 net3 sky130_fd_pr__nfet_01v8 L=24.000 W=0.360 nf=1
XM5 net3 net1 Vn Vn sky130_fd_pr__nfet_01v8 L=24.000 W=0.360 nf=1
.ends th02


.subckt th03 Vp Vin Vout Vn
XM7 Vout net1 Vp Vp sky130_fd_pr__pfet_01v8 L=0.150 W=2.3000 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=2.2000 W=0.360 nf=1
XM1 net1 Vin net2 net2 sky130_fd_pr__pfet_01v8 L=5.000 W=0.42 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=5.000 nf=1
XM2 Vp Vp net2 net2 sky130_fd_pr__nfet_01v8 L=5.0 W=0.36 nf=1
.ends th03


.subckt th04 Vp Vout Vin Vn
XM7 Vout net1 Vp Vp sky130_fd_pr__pfet_01v8 L=1.000 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.000 nf=1
XM1 net1 Vin net2 net2 sky130_fd_pr__pfet_01v8 L=1.000 W=0.42 nf=1
XM1 net1 Vin net2 net2 sky130_fd_pr__pfet_01v8 L=1.000 W=0.42 nf=1
XM1 net1 Vin net2 net2 sky130_fd_pr__pfet_01v8 L=1.000 W=0.42 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.000 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.000 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.000 nf=1
XM2 Vp Vp net2 net2 sky130_fd_pr__nfet_01v8 L=0.15 W=0.46300 nf=1
XM2 Vp Vp net2 net2 sky130_fd_pr__nfet_01v8 L=0.15 W=0.46300 nf=1
XM2 Vp Vp net2 net2 sky130_fd_pr__nfet_01v8 L=0.15 W=0.46300 nf=1
.ends th04


.subckt th05 Vp Vout Vin Vn
XM7 Vout net1 Vp Vp sky130_fd_pr__pfet_01v8 L=1.12000 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.12000 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.12000 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.12000 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=2.000 W=0.42 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=2.000 W=0.42 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=2.000 W=0.42 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=2.00 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=2.00 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=2.00 nf=1
.ends th05


.subckt th06 Vp Vout Vin Vn
XM7 Vout net1 Vp Vp sky130_fd_pr__pfet_01v8 L=0.436000 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.46000 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.46000 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.46000 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.47000 W=0.42 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.47000 W=0.42 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.47000 W=0.42 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.3900 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.3900 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.3900 nf=1
.ends th06


.subckt th07 Vp Vout Vin Vn
XM7 Vout net1 Vp Vp sky130_fd_pr__pfet_01v8 L=0.47000 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.46000 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.46000 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.46000 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.151 W=0.42 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.151 W=0.42 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.151 W=0.42 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.155 W=0.36 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.155 W=0.36 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.155 W=0.36 nf=1
.ends th07


.subckt th08 Vp Vout Vin Vn
XM7 Vout net1 Vp Vp sky130_fd_pr__pfet_01v8 L=0.47 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.468 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.468 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.468 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=0.67 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=0.67 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=0.67 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.67 W=0.36 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.67 W=0.36 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.67 W=0.36 nf=1
.ends th08


.subckt th09 Vp Vout Vin Vn
XM7 net2 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=1.58 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=1.58 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=1.58 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=1.58 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.57 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.57 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.57 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=1.58 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=1.58 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=1.58 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=1.58 W=0.36 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=1.58 W=0.36 nf=1
XM3 net1 Vin Vn Vn sky130_fd_pr__nfet_01v8 L=1.58 W=0.36 nf=1
.ends th09


.subckt th10 Vp Vout Vin Vn
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=0.15 W=0.36 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=0.15 W=0.36 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=0.15 W=0.36 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
XM7 net2 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1
XM7 net2 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1
XM7 net2 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1
.ends th10


.subckt th11 Vp Vout Vin Vn
XM7 net2 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=1.42 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=1.42 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=1.42 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=1.42 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1.42 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=1.42 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=1.42 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=1.42 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=1.42 W=0.36 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=1.42 W=0.36 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=1.42 W=0.36 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
.ends th11


.subckt th12 Vp Vout Vin Vn
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=2.92 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=2.92 W=0.36 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=2.92 W=0.36 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=2.92 W=0.36 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
XM7 net2 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=2.92 W=0.42 nf=1
XM7 net2 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=2.92 W=0.42 nf=1
XM7 net2 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=2.92 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=2.92 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=2.92 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=2.92 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=2.92 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=2.92 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=2.92 nf=1
.ends th12


.subckt th13 Vp Vout Vin Vn
XM4 net2 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=13.8 W=0.42 nf=1
XM5 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=13.8 W=0.42 nf=1
XM5 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=13.8 W=0.42 nf=1
XM5 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=13.8 W=0.42 nf=1
XM6 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=13.8 nf=1
XM6 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=13.8 nf=1
XM6 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=13.8 nf=1
XM8 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=5.5 nf=1
XM8 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=5.5 nf=1
XM8 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=5.5 nf=1
XM11 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=5.5 W=0.36 nf=1
XM11 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=5.5 W=0.36 nf=1
XM11 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=5.5 W=0.36 nf=1
XM12 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
XM12 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
XM12 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1
.ends th13


.subckt th14 Vp Vout Vin Vn
XM7 net2 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=25 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=25 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=25 W=0.42 nf=1
XM9 Vout net1 net2 net2 sky130_fd_pr__pfet_01v8 L=25 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=25 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=25 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=25 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=19.5 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=19.5 nf=1
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=19.5 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=19.5 W=0.36 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=19.5 W=0.36 nf=1
XM3 net1 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=19.5 W=0.36 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=0.69 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=0.69 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=0.69 nf=1
.ends th14


.subckt th15 Vp Vout Vin Vn
XM1 net1 Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=25 nf=1
XM3 net2 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=25 W=0.36 nf=1
XM3 net2 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=25 W=0.36 nf=1
XM3 net2 Vin net3 net3 sky130_fd_pr__nfet_01v8 L=25 W=0.36 nf=1
XM4 net1 Vin net2 net2 sky130_fd_pr__nfet_01v8 L=25 W=0.36 nf=1
XM4 net1 Vin net2 net2 sky130_fd_pr__nfet_01v8 L=25 W=0.36 nf=1
XM4 net1 Vin net2 net2 sky130_fd_pr__nfet_01v8 L=25 W=0.36 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.2 W=1 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.2 W=1 nf=1
XM2 Vn Vn net3 net3 sky130_fd_pr__pfet_01v8 L=0.2 W=1 nf=1
XM7 net4 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=25 W=0.42 nf=1
XM7 net4 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=25 W=0.42 nf=1
XM7 net4 net1 Vp Vp sky130_fd_pr__pfet_01v8 L=25 W=0.42 nf=1
XM9 Vout net1 net4 net4 sky130_fd_pr__pfet_01v8 L=25 W=0.42 nf=1
XM9 Vout net1 net4 net4 sky130_fd_pr__pfet_01v8 L=25 W=0.42 nf=1
XM9 Vout net1 net4 net4 sky130_fd_pr__pfet_01v8 L=25 W=0.42 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=25 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=25 nf=1
XM10 Vout net1 Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=25 nf=1
.ends th15


.subckt Analog Vp Vin V1 V2 V3 V4 V5 V6 V7 V8 V9 V10 V11 V12 V13 V14 V15 Vn
x1 Vp Vin V1 Vn th01
x2 Vp V2 Vin Vn th02
x3 Vp Vin V3 Vn th03
x4 Vp V4 Vin Vn th04
x5 Vp V5 Vin Vn th05
x6 Vp V6 Vin Vn th06
x7 Vp V7 Vin Vn th07
x8 Vp V8 Vin Vn th08
x9 Vp V9 Vin Vn th09
x10 Vp V10 Vin Vn th10
x11 Vp V11 Vin Vn th11
x12 Vp V12 Vin Vn th12
x13 Vp V13 Vin Vn th13
x14 Vp V14 Vin Vn th14
x15 Vp V15 Vin Vn th15
.ends Analog


sky130_fd_sc_hd__clkinv_1
sky130_fd_sc_hd__and2_0
sky130_fd_sc_hd__nand3_1
sky130_fd_sc_hd__a22oi_1
sky130_fd_sc_hd__or3_1
sky130_fd_sc_hd__lpflow_inputiso1p_1
sky130_fd_sc_hd__nand2b_1
sky130_fd_sc_hd__nor4b_1
sky130_fd_sc_hd__nor4_1
sky130_fd_sc_hd__or3b_1
sky130_fd_sc_hd__or4_1
sky130_fd_sc_hd__a211oi_1
sky130_fd_sc_hd__a32oi_1 
sky130_fd_sc_hd__o2111ai_1
sky130_fd_sc_hd__nand3b_1
sky130_fd_sc_hd__nor3_1
sky130_fd_sc_hd__nand4_1
sky130_fd_sc_hd__nor2_1
sky130_fd_sc_hd__o21ai_0
sky130_fd_sc_hd__o31ai_1
sky130_fd_sc_hd__nand2_1




.subckt analog_therm b0 Vin b1 b2 b3 Vp Vn
x0 p10 VGND VNB VPB VPWR 1 sky130_fd_sc_hd__clkinv_1
x1 p1 p0 VGND VNB VPB VPWR 2 sky130_fd_sc_hd__nand2_1
x2 p1 p0 p2 VGND VNB VPB VPWR 3 sky130_fd_sc_hd__nand3_1
x3 p1 p0 p3 p2 VGND VNB VPB VPWR 4 sky130_fd_sc_hd__nand4_1
x4 p5 p4 VGND VNB VPB VPWR 5 sky130_fd_sc_hd__nand2_1
x5 p5 p4 p7 p6 VGND VNB VPB VPWR 6 sky130_fd_sc_hd__nand4_1
x6 4 6 VGND VNB VPB VPWR 7 sky130_fd_sc_hd__nor2_1
x7 p8 p9 VGND VNB VPB VPWR 8 sky130_fd_sc_hd__nand2_1
x8 p11 p10 VGND VNB VPB VPWR 9 sky130_fd_sc_hd__nand2_1
x9 4 6 8 9 VGND VNB VPB VPWR 10 sky130_fd_sc_hd__nor4_1
x10 p13 p12 VGND VNB VPB VPWR 11 sky130_fd_sc_hd__and2_0
x11 10 11 VGND VNB VPB VPWR 12 sky130_fd_sc_hd__nand2_1
x12 p14 10 11 VGND VNB VPB VPWR 13 sky130_fd_sc_hd__nand3_1
x13 p7 5 VGND VNB VPB VPWR 14 sky130_fd_sc_hd__nor2_1
x14 p5 p7 p6 VGND VNB VPB VPWR 15 sky130_fd_sc_hd__nor3_1
x15 p6 14 15 p4 VGND VNB VPB VPWR 16 sky130_fd_sc_hd__a22oi_1
x16 p13 p14 VGND VNB VPB VPWR 17 sky130_fd_sc_hd__nor2_1
x17 p13 p12 p14 VGND VNB VPB VPWR 18 sky130_fd_sc_hd__or3_1
x18 p11 p10 VGND VNB VPB VPWR 19 sky130_fd_sc_hd__lpflow_inputiso1p_1
x19 p8 p9 18 19 VGND VNB VPB VPWR 20 sky130_fd_sc_hd__nor4_1
x20 4 20 VGND VNB VPB VPWR 21 sky130_fd_sc_hd__nand2b_1
x21 p9 18 19 p8 VGND VNB VPB VPWR 22 sky130_fd_sc_hd__nor4b_1
x22 p11 8 18 VGND VNB VPB VPWR 23 sky130_fd_sc_hd__nor3_1
x23 p11 1 8 18 VGND VNB VPB VPWR 24 sky130_fd_sc_hd__nor4_1
x24 22 24 7 VGND VNB VPB VPWR 25 sky130_fd_sc_hd__o21ai_0
x25 p1 p2 p0 VGND VNB VPB VPWR 26 sky130_fd_sc_hd__or3b_1
x26 p5 p4 p7 p6 VGND VNB VPB VPWR 27 sky130_fd_sc_hd__or4_1
x27 3 26 27 p3 VGND VNB VPB VPWR 28 sky130_fd_sc_hd__a211oi_1
x28 p12 10 17 20 28 VGND VNB VPB VPWR 29 sky130_fd_sc_hd__a32oi_1
x29 16 21 25 29 13 VGND VNB VPB VPWR b0 sky130_fd_sc_hd__o2111ai_1
x30 4 14 20 VGND VNB VPB VPWR 30 sky130_fd_sc_hd__nand3b_1
x31 7 23 VGND VNB VPB VPWR 31 sky130_fd_sc_hd__nand2_1
x32 p3 2 27 VGND VNB VPB VPWR 32 sky130_fd_sc_hd__nor3_1
x33 20 32 VGND VNB VPB VPWR 33 sky130_fd_sc_hd__nand2_1
x34 12 30 31 33 VGND VNB VPB VPWR b1 sky130_fd_sc_hd__nand4_1
x35 11 17 10 VGND VNB VPB VPWR 34 sky130_fd_sc_hd__o21ai_0
x36 14 15 VGND VNB VPB VPWR 35 sky130_fd_sc_hd__nor2_1
x37 21 35 34 VGND VNB VPB VPWR b2 sky130_fd_sc_hd__o21ai_0
x38 20 22 23 7 VGND VNB VPB VPWR 36 sky130_fd_sc_hd__o31ai_1
x39 34 36 VGND VNB VPB VPWR b3 sky130_fd_sc_hd__nand2_1
x40 Vp Vin p0 p1 p2 p3 p4 p5 p6 p7 p8 p9 p10 p11 p12 p13 p14 Vn Analog
.ends analog_therm
