magic
tech sky130A
magscale 1 2
timestamp 1706629535
<< metal1 >>
rect 1128 9174 1180 9180
rect 1097 9118 1128 9163
rect 1097 9112 1180 9118
rect 1097 7742 1131 9112
rect 1097 7457 1135 7742
rect 1101 3389 1135 7457
rect 4768 6510 4868 6610
rect 4807 6415 4841 6510
rect 4807 6381 4945 6415
rect 3869 6162 3903 6253
rect 5204 6174 6270 6202
rect 3836 6062 3936 6162
rect 1232 5870 1238 5922
rect 1294 5870 1300 5922
rect 4838 5866 4890 5872
rect 4838 5808 4890 5814
rect 5003 5388 5009 5440
rect 5061 5388 5067 5440
rect 5204 5190 5232 6174
rect 5963 5384 5969 5436
rect 6021 5429 6027 5436
rect 6021 5392 6364 5429
rect 6021 5384 6027 5392
rect 4788 5162 5232 5190
rect 4788 4604 4816 5162
rect 5130 4610 6372 4638
rect 1370 4428 1422 4434
rect 1370 4366 1422 4372
rect 5130 3796 5158 4610
rect 6224 4406 6280 4434
rect 4730 3768 5158 3796
rect 4600 3418 4606 3470
rect 4658 3418 4664 3470
rect 1294 3401 1346 3407
rect 1101 3355 1294 3389
rect 1294 3343 1346 3349
rect 2344 3401 2396 3407
rect 2344 3343 2396 3349
rect 4730 3104 4758 3768
rect 5310 3644 5362 3650
rect 5310 3586 5362 3592
rect 4715 3052 4721 3104
rect 4773 3052 4779 3104
rect 5310 2446 5338 3586
rect 4582 2418 5338 2446
rect 3984 2212 3990 2264
rect 4042 2212 4048 2264
rect 3999 1873 4033 2212
rect 3959 1839 4033 1873
rect 1476 1664 1528 1670
rect 1476 1602 1528 1608
rect 4582 726 4610 2418
rect 9268 2286 9320 2292
rect 7442 2230 7448 2286
rect 7504 2275 7510 2286
rect 7504 2241 9268 2275
rect 7504 2230 7510 2241
rect 9268 2224 9320 2230
rect 8654 2126 8706 2132
rect 6674 2064 6680 2116
rect 6736 2115 6742 2116
rect 6736 2081 8654 2115
rect 6736 2064 6742 2081
rect 8654 2064 8706 2070
rect 8020 1928 8072 1934
rect 5831 1914 8020 1917
rect 5782 1862 5788 1914
rect 5844 1883 8020 1914
rect 5844 1862 5850 1883
rect 8020 1866 8072 1872
rect 7844 1786 7896 1792
rect 4446 698 4610 726
rect 4661 1741 7844 1775
rect 4661 -37 4695 1741
rect 7844 1724 7896 1730
rect 7442 1659 7448 1668
rect 7421 1616 7448 1659
rect 7504 1616 7510 1668
rect 5630 1196 5682 1202
rect 5630 1134 5682 1140
rect 6598 768 6604 820
rect 6660 768 6666 820
rect 7421 599 7455 1616
rect 9580 1218 9680 3754
rect 8398 726 8404 778
rect 8460 726 8466 778
rect 9608 610 9660 616
rect 9608 548 9660 554
rect 5327 175 5361 261
rect 5458 175 5558 216
rect 5327 141 5558 175
rect 5458 116 5558 141
rect 2101 -189 2135 -43
rect 2701 -71 4695 -37
rect 2701 -189 2735 -71
rect 2101 -223 2735 -189
<< via1 >>
rect 1128 9118 1180 9174
rect 1238 5870 1294 5922
rect 4838 5814 4890 5866
rect 5009 5388 5061 5440
rect 5969 5384 6021 5436
rect 1370 4372 1422 4428
rect 4606 3418 4658 3470
rect 1294 3349 1346 3401
rect 2344 3349 2396 3401
rect 5310 3592 5362 3644
rect 4721 3052 4773 3104
rect 3990 2212 4042 2264
rect 1476 1608 1528 1664
rect 7448 2230 7504 2286
rect 9268 2230 9320 2286
rect 6680 2064 6736 2116
rect 8654 2070 8706 2126
rect 5788 1862 5844 1914
rect 8020 1872 8072 1928
rect 7844 1730 7896 1786
rect 7448 1616 7504 1668
rect 5630 1140 5682 1196
rect 6604 768 6660 820
rect 8404 726 8460 778
rect 9608 554 9660 610
<< metal2 >>
rect 948 10194 8544 10250
rect 948 4428 1004 10194
rect 1433 9201 1489 9210
rect 1122 9118 1128 9174
rect 1180 9118 1433 9174
rect 1433 9082 1489 9091
rect 5096 7773 5105 7787
rect 4978 7745 5105 7773
rect 1207 5936 1216 5992
rect 1316 5936 1325 5992
rect 1238 5922 1294 5936
rect 1238 5864 1294 5870
rect 4832 5814 4838 5866
rect 4890 5854 4896 5866
rect 4978 5854 5006 7745
rect 5096 7731 5105 7745
rect 5215 7731 5224 7787
rect 4890 5826 5006 5854
rect 4890 5814 4896 5826
rect 5314 5485 5323 5541
rect 5433 5485 5442 5541
rect 5009 5440 5061 5446
rect 5007 5388 5009 5392
rect 5061 5388 5063 5392
rect 5007 5383 5063 5388
rect 5007 5264 5063 5273
rect 5361 4951 5395 5485
rect 5969 5436 6021 5442
rect 5967 5384 5969 5392
rect 6021 5384 6023 5392
rect 5967 5383 6023 5384
rect 5967 5264 6023 5273
rect 5041 4917 5395 4951
rect 948 4372 1370 4428
rect 1422 4372 1428 4428
rect 5041 3723 5075 4917
rect 4615 3689 5075 3723
rect 4615 3476 4649 3689
rect 5304 3592 5310 3644
rect 5362 3632 5368 3644
rect 5362 3604 6690 3632
rect 5362 3592 5368 3604
rect 4606 3470 4658 3476
rect 4606 3412 4658 3418
rect 1288 3349 1294 3401
rect 1346 3392 1352 3401
rect 2338 3392 2344 3401
rect 1346 3358 2344 3392
rect 1346 3349 1352 3358
rect 2338 3349 2344 3358
rect 2396 3349 2402 3401
rect 4721 3104 4773 3110
rect 4721 3046 4773 3052
rect 4730 2645 4764 3046
rect 3999 2611 4764 2645
rect 3999 2270 4033 2611
rect 4730 2602 4764 2611
rect 7448 2286 7504 2292
rect 3990 2264 4042 2270
rect 3990 2206 4042 2212
rect 9262 2230 9268 2286
rect 9320 2230 9832 2286
rect 6680 2116 6736 2122
rect 5788 1914 5844 1920
rect 1196 1608 1476 1664
rect 1528 1608 1534 1664
rect 1196 -360 1252 1608
rect 5788 1492 5844 1862
rect 5694 1436 5844 1492
rect 5694 1196 5750 1436
rect 6680 1412 6736 2064
rect 7448 1668 7504 2230
rect 8648 2070 8654 2126
rect 8706 2070 9188 2126
rect 8014 1872 8020 1928
rect 8072 1872 8544 1928
rect 7838 1730 7844 1786
rect 7896 1730 7902 1786
rect 7200 1534 7256 1658
rect 7448 1610 7504 1616
rect 9904 1598 10476 1654
rect 10728 1604 11120 1660
rect 9904 1534 9960 1598
rect 7200 1478 7566 1534
rect 5624 1140 5630 1196
rect 5682 1140 5750 1196
rect 6604 1356 6736 1412
rect 6604 820 6660 1356
rect 6604 762 6660 768
rect 7510 -360 7566 1478
rect 8404 1478 9960 1534
rect 8404 778 8460 1478
rect 8404 720 8460 726
rect 10728 610 10784 1604
rect 9602 554 9608 610
rect 9660 554 10784 610
rect 1196 -416 7566 -360
<< via2 >>
rect 1433 9091 1489 9201
rect 1216 5936 1316 5992
rect 5105 7731 5215 7787
rect 5323 5485 5433 5541
rect 5007 5273 5063 5383
rect 5967 5273 6023 5383
<< metal3 >>
rect 1428 9201 5404 9206
rect 1428 9091 1433 9201
rect 1489 9091 5404 9201
rect 1428 9086 5404 9091
rect 1211 8411 5473 8521
rect 1211 5992 1321 8411
rect 5100 7787 5370 7846
rect 5100 7731 5105 7787
rect 5215 7731 5370 7787
rect 5100 7726 5370 7731
rect 1211 5936 1216 5992
rect 1316 5936 1321 5992
rect 1211 5931 1321 5936
rect 5318 5541 5438 5806
rect 5318 5485 5323 5541
rect 5433 5485 5438 5541
rect 5318 5480 5438 5485
rect 5002 5383 6028 5388
rect 5002 5273 5007 5383
rect 5063 5273 5967 5383
rect 6023 5273 6028 5383
rect 5002 5268 6028 5273
use Analog  Analog_0
timestamp 1706548588
transform 1 0 -336 0 1 6974
box 1538 -7112 10018 -488
use therm_raw  therm_raw_0
timestamp 1705015937
transform 1 0 5250 0 1 1598
box 0 0 7058 9202
<< labels >>
flabel metal1 5458 116 5558 216 0 FreeSans 256 0 0 0 Vp
port 30 nsew
flabel metal1 4768 6510 4868 6610 0 FreeSans 256 180 0 0 Vn
port 31 nsew
flabel metal1 3836 6062 3936 6162 0 FreeSans 256 0 0 0 Vin
port 32 nsew
<< end >>
