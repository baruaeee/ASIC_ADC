magic
tech sky130A
magscale 1 2
timestamp 1703627557
<< obsli1 >>
rect 1104 2159 5888 6545
<< obsm1 >>
rect 934 2128 5888 6576
<< metal2 >>
rect 3238 8402 3294 9202
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
<< obsm2 >>
rect 938 8346 3182 8402
rect 3350 8346 5868 8402
rect 938 856 5868 8346
rect 938 800 1250 856
rect 1418 800 1894 856
rect 2062 800 2538 856
rect 2706 800 3182 856
rect 3350 800 3826 856
rect 3994 800 4470 856
rect 4638 800 5114 856
rect 5282 800 5758 856
<< metal3 >>
rect 0 7488 800 7608
rect 0 6808 800 6928
rect 0 6128 800 6248
rect 0 5448 800 5568
rect 6258 5448 7058 5568
rect 0 4768 800 4888
rect 6258 4768 7058 4888
rect 0 4088 800 4208
rect 0 3408 800 3528
rect 0 2728 800 2848
<< obsm3 >>
rect 880 7408 6258 7581
rect 800 7008 6258 7408
rect 880 6728 6258 7008
rect 800 6328 6258 6728
rect 880 6048 6258 6328
rect 800 5648 6258 6048
rect 880 5368 6178 5648
rect 800 4968 6258 5368
rect 880 4688 6178 4968
rect 800 4288 6258 4688
rect 880 4008 6258 4288
rect 800 3608 6258 4008
rect 880 3328 6258 3608
rect 800 2928 6258 3328
rect 880 2648 6258 2928
rect 800 2143 6258 2648
<< metal4 >>
rect 2744 2128 3064 6576
rect 3404 2128 3724 6576
<< labels >>
rlabel metal4 s 3404 2128 3724 6576 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2744 2128 3064 6576 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 6258 5448 7058 5568 6 b[0]
port 3 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 b[1]
port 4 nsew signal output
rlabel metal3 s 6258 4768 7058 4888 6 b[2]
port 5 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 b[3]
port 6 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 p[0]
port 7 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 p[10]
port 8 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 p[11]
port 9 nsew signal input
rlabel metal2 s 3238 8402 3294 9202 6 p[12]
port 10 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 p[13]
port 11 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 p[14]
port 12 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 p[1]
port 13 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 p[2]
port 14 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 p[3]
port 15 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 p[4]
port 16 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 p[5]
port 17 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 p[6]
port 18 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 p[7]
port 19 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 p[8]
port 20 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 p[9]
port 21 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 7058 9202
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 287084
string GDS_FILE /openlane/designs/ADC/runs/RUN_2023.12.26_21.49.15/results/signoff/ADC.magic.gds
string GDS_START 160928
<< end >>

