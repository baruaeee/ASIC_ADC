* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : pre_therm                                    *
* Netlisted  : Fri Dec  6 04:50:32 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733457022020                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733457022020 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6.5e-07 W=4.45e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733457022020

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733457022021                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733457022021 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=6.3e-07 W=7.9e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733457022021

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv01f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv01f VDD VSS A Y
** N=9 EP=4 FDC=2
X3 VSS Y A nfet_01v8_CDNS_733457022020 $T=295 475 0 0 $X=-110 $Y=325
X4 VDD Y A pfet_01v8_CDNS_733457022021 $T=295 2820 0 0 $X=-150 $Y=2640
.ends inv01f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733457022022                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733457022022 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 pfet_01v8 L=1.05e-06 W=5.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733457022022

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733457022023                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733457022023 1 2 3 4
** N=10 EP=4 FDC=1
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=1.02e-06 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733457022023

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: preampF                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt preampF VDD VSS A Y
** N=9 EP=4 FDC=2
X5 Y VSS A VDD pfet_01v8_CDNS_733457022022 $T=825 3430 0 270 $X=645 $Y=1935
X6 Y VDD A VSS nfet_01v8_CDNS_733457022023 $T=430 485 1 180 $X=-125 $Y=335
.ends preampF

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pre_therm                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pre_therm
** N=6 EP=0 FDC=4
X4 4 5 2 3 inv01f $T=1740 9060 1 0 $X=1560 $Y=4615
X5 4 5 1 2 preampF $T=0 9060 1 0 $X=-180 $Y=4615
.ends pre_therm
