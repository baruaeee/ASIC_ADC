* NGSPICE file created from th07.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_VGVEGU a_n74_n42# a_n33_n130# a_n176_n216# a_16_n42#
X0 a_16_n42# a_n33_n130# a_n74_n42# a_n176_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.16
C0 a_16_n42# a_n74_n42# 0.0684f
C1 a_16_n42# a_n33_n130# 0.0191f
C2 a_n74_n42# a_n33_n130# 0.0191f
C3 a_16_n42# a_n176_n216# 0.0737f
C4 a_n74_n42# a_n176_n216# 0.0737f
C5 a_n33_n130# a_n176_n216# 0.338f
.ends

.subckt sky130_fd_pr__pfet_01v8_EDPLE3 a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n42# a_n33_n139# 0.0192f
C1 a_n73_n42# w_n211_n261# 0.0463f
C2 a_n73_n42# a_15_n42# 0.0699f
C3 a_n33_n139# w_n211_n261# 0.236f
C4 a_n33_n139# a_15_n42# 0.0192f
C5 w_n211_n261# a_15_n42# 0.0463f
C6 a_15_n42# VSUBS 0.0263f
C7 a_n73_n42# VSUBS 0.0263f
C8 a_n33_n139# VSUBS 0.115f
C9 w_n211_n261# VSUBS 1.03f
.ends

.subckt sky130_fd_pr__pfet_01v8_NZD9V2 w_n243_n261# a_47_n42# a_n47_n139# a_n105_n42#
+ VSUBS
X0 a_47_n42# a_n47_n139# a_n105_n42# w_n243_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.47
C0 a_n105_n42# a_n47_n139# 0.00866f
C1 a_n105_n42# w_n243_n261# 0.0499f
C2 a_n105_n42# a_47_n42# 0.0406f
C3 a_n47_n139# w_n243_n261# 0.27f
C4 a_n47_n139# a_47_n42# 0.00866f
C5 w_n243_n261# a_47_n42# 0.0499f
C6 a_47_n42# VSUBS 0.0297f
C7 a_n105_n42# VSUBS 0.0297f
C8 a_n47_n139# VSUBS 0.168f
C9 w_n243_n261# VSUBS 1.17f
.ends

.subckt sky130_fd_pr__nfet_01v8_97T34Z a_n73_n46# a_n175_n220# a_n33_n134# a_15_n46#
X0 a_15_n46# a_n33_n134# a_n73_n46# a_n175_n220# sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.5 as=0.133 ps=1.5 w=0.46 l=0.15
C0 a_15_n46# a_n73_n46# 0.0763f
C1 a_15_n46# a_n33_n134# 0.0212f
C2 a_n73_n46# a_n33_n134# 0.0212f
C3 a_15_n46# a_n175_n220# 0.0769f
C4 a_n73_n46# a_n175_n220# 0.0769f
C5 a_n33_n134# a_n175_n220# 0.338f
.ends

.subckt th07 Vp Vin V07 Vn
XXM0 m1_400_n1066# Vin Vn Vn sky130_fd_pr__nfet_01v8_VGVEGU
XXM1 m1_400_n1066# Vp Vin Vp Vn sky130_fd_pr__pfet_01v8_EDPLE3
XXM2 Vp V07 m1_400_n1066# Vp Vn sky130_fd_pr__pfet_01v8_NZD9V2
XXM3 Vn Vn m1_400_n1066# V07 sky130_fd_pr__nfet_01v8_97T34Z
C0 m1_400_n1066# Vp 0.32f
C1 Vin V07 6.52e-19
C2 Vp V07 0.102f
C3 m1_400_n1066# V07 0.167f
C4 Vin Vp 0.212f
C5 m1_400_n1066# Vin 0.436f
C6 Vin Vn 0.75f
C7 m1_400_n1066# Vn 0.943f
C8 V07 Vn 0.395f
C9 Vp Vn 2.43f
.ends

