magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 148 29 154
rect -29 114 -17 148
rect -29 108 29 114
rect -29 -114 29 -108
rect -29 -148 -17 -114
rect -29 -154 29 -148
<< nwell >>
rect -211 -286 211 286
<< pmos >>
rect -15 -67 15 67
<< pdiff >>
rect -73 55 -15 67
rect -73 -55 -61 55
rect -27 -55 -15 55
rect -73 -67 -15 -55
rect 15 55 73 67
rect 15 -55 27 55
rect 61 -55 73 55
rect 15 -67 73 -55
<< pdiffc >>
rect -61 -55 -27 55
rect 27 -55 61 55
<< nsubdiff >>
rect -175 216 -79 250
rect 79 216 175 250
rect -175 154 -141 216
rect 141 154 175 216
rect -175 -216 -141 -154
rect 141 -216 175 -154
rect -175 -250 -79 -216
rect 79 -250 175 -216
<< nsubdiffcont >>
rect -79 216 79 250
rect -175 -154 -141 154
rect 141 -154 175 154
rect -79 -250 79 -216
<< poly >>
rect -33 148 33 164
rect -33 114 -17 148
rect 17 114 33 148
rect -33 98 33 114
rect -15 67 15 98
rect -15 -98 15 -67
rect -33 -114 33 -98
rect -33 -148 -17 -114
rect 17 -148 33 -114
rect -33 -164 33 -148
<< polycont >>
rect -17 114 17 148
rect -17 -148 17 -114
<< locali >>
rect -175 216 -79 250
rect 79 216 175 250
rect -175 154 -141 216
rect 141 154 175 216
rect -33 114 -17 148
rect 17 114 33 148
rect -61 55 -27 71
rect -61 -71 -27 -55
rect 27 55 61 71
rect 27 -71 61 -55
rect -33 -148 -17 -114
rect 17 -148 33 -114
rect -175 -216 -141 -154
rect 141 -216 175 -154
rect -175 -250 -79 -216
rect 79 -250 175 -216
<< viali >>
rect -17 114 17 148
rect -61 -55 -27 55
rect 27 -55 61 55
rect -17 -148 17 -114
<< metal1 >>
rect -29 148 29 154
rect -29 114 -17 148
rect 17 114 29 148
rect -29 108 29 114
rect -67 55 -21 67
rect -67 -55 -61 55
rect -27 -55 -21 55
rect -67 -67 -21 -55
rect 21 55 67 67
rect 21 -55 27 55
rect 61 -55 67 55
rect 21 -67 67 -55
rect -29 -114 29 -108
rect -29 -148 -17 -114
rect 17 -148 29 -114
rect -29 -154 29 -148
<< properties >>
string FIXED_BBOX -158 -233 158 233
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.67 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
