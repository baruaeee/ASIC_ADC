magic
tech sky130A
magscale 1 2
timestamp 1704301096
<< error_p >>
rect -29 1131 29 1137
rect -29 1097 -17 1131
rect -29 1091 29 1097
rect -29 -1097 29 -1091
rect -29 -1131 -17 -1097
rect -29 -1137 29 -1131
<< nwell >>
rect -211 -1269 211 1269
<< pmos >>
rect -15 -1050 15 1050
<< pdiff >>
rect -73 1038 -15 1050
rect -73 -1038 -61 1038
rect -27 -1038 -15 1038
rect -73 -1050 -15 -1038
rect 15 1038 73 1050
rect 15 -1038 27 1038
rect 61 -1038 73 1038
rect 15 -1050 73 -1038
<< pdiffc >>
rect -61 -1038 -27 1038
rect 27 -1038 61 1038
<< nsubdiff >>
rect -175 1199 -79 1233
rect 79 1199 175 1233
rect -175 1137 -141 1199
rect 141 1137 175 1199
rect -175 -1199 -141 -1137
rect 141 -1199 175 -1137
rect -175 -1233 -79 -1199
rect 79 -1233 175 -1199
<< nsubdiffcont >>
rect -79 1199 79 1233
rect -175 -1137 -141 1137
rect 141 -1137 175 1137
rect -79 -1233 79 -1199
<< poly >>
rect -33 1131 33 1147
rect -33 1097 -17 1131
rect 17 1097 33 1131
rect -33 1081 33 1097
rect -15 1050 15 1081
rect -15 -1081 15 -1050
rect -33 -1097 33 -1081
rect -33 -1131 -17 -1097
rect 17 -1131 33 -1097
rect -33 -1147 33 -1131
<< polycont >>
rect -17 1097 17 1131
rect -17 -1131 17 -1097
<< locali >>
rect -175 1199 -79 1233
rect 79 1199 175 1233
rect -175 1137 -141 1199
rect 141 1137 175 1199
rect -33 1097 -17 1131
rect 17 1097 33 1131
rect -61 1038 -27 1054
rect -61 -1054 -27 -1038
rect 27 1038 61 1054
rect 27 -1054 61 -1038
rect -33 -1131 -17 -1097
rect 17 -1131 33 -1097
rect -175 -1199 -141 -1137
rect 141 -1199 175 -1137
rect -175 -1233 -79 -1199
rect 79 -1233 175 -1199
<< viali >>
rect -17 1097 17 1131
rect -61 -1038 -27 1038
rect 27 -1038 61 1038
rect -17 -1131 17 -1097
<< metal1 >>
rect -29 1131 29 1137
rect -29 1097 -17 1131
rect 17 1097 29 1131
rect -29 1091 29 1097
rect -67 1038 -21 1050
rect -67 -1038 -61 1038
rect -27 -1038 -21 1038
rect -67 -1050 -21 -1038
rect 21 1038 67 1050
rect 21 -1038 27 1038
rect 61 -1038 67 1038
rect 21 -1050 67 -1038
rect -29 -1097 29 -1091
rect -29 -1131 -17 -1097
rect 17 -1131 29 -1097
rect -29 -1137 29 -1131
<< properties >>
string FIXED_BBOX -158 -1216 158 1216
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
