* NGSPICE file created from th06.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_DD6SHA a_n33_n130# a_15_n42# a_n175_n182# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_15_n42# a_n73_n42# 0.0699f
C1 a_15_n42# a_n33_n130# 0.0209f
C2 a_n73_n42# a_n33_n130# 0.0209f
C3 a_15_n42# a_n175_n182# 0.0637f
C4 a_n73_n42# a_n175_n182# 0.0716f
C5 a_n33_n130# a_n175_n182# 0.314f
.ends

.subckt sky130_fd_pr__pfet_01v8_7DPLFP w_n245_n261# a_n107_n42# a_n49_n139# a_49_n42#
+ VSUBS
X0 a_49_n42# a_n49_n139# a_n107_n42# w_n245_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.49
C0 a_n107_n42# a_n49_n139# 0.00895f
C1 a_n107_n42# w_n245_n261# 0.0224f
C2 a_49_n42# a_n107_n42# 0.0396f
C3 a_n49_n139# w_n245_n261# 0.221f
C4 a_49_n42# a_n49_n139# 0.00895f
C5 a_49_n42# w_n245_n261# 0.0224f
C6 a_49_n42# VSUBS 0.0487f
C7 a_n107_n42# VSUBS 0.0487f
C8 a_n49_n139# VSUBS 0.206f
C9 w_n245_n261# VSUBS 0.876f
.ends

.subckt sky130_fd_pr__pfet_01v8_MDPZBH a_n102_n42# a_44_n42# a_n44_n139# w_n240_n261#
+ VSUBS
X0 a_44_n42# a_n44_n139# a_n102_n42# w_n240_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.44
C0 a_n102_n42# a_n44_n139# 0.00823f
C1 a_n102_n42# w_n240_n261# 0.0224f
C2 a_44_n42# a_n102_n42# 0.0423f
C3 a_n44_n139# w_n240_n261# 0.208f
C4 a_44_n42# a_n44_n139# 0.00823f
C5 a_44_n42# w_n240_n261# 0.0224f
C6 a_44_n42# VSUBS 0.0485f
C7 a_n102_n42# VSUBS 0.0485f
C8 a_n44_n139# VSUBS 0.191f
C9 w_n240_n261# VSUBS 0.858f
.ends

.subckt sky130_fd_pr__nfet_01v8_MYA4RC a_n73_n46# a_n33_n134# a_15_n46# a_n175_n186#
X0 a_15_n46# a_n33_n134# a_n73_n46# a_n175_n186# sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.5 as=0.133 ps=1.5 w=0.46 l=0.15
C0 a_15_n46# a_n73_n46# 0.0763f
C1 a_15_n46# a_n33_n134# 0.0212f
C2 a_n73_n46# a_n33_n134# 0.0212f
C3 a_15_n46# a_n175_n186# 0.0671f
C4 a_n73_n46# a_n175_n186# 0.0756f
C5 a_n33_n134# a_n175_n186# 0.314f
.ends

.subckt th06 Vp Vin V06 Vn
XXM0 Vin m1_904_n796# Vn Vn sky130_fd_pr__nfet_01v8_DD6SHA
XXM1 Vp Vp Vin m1_904_n796# Vn sky130_fd_pr__pfet_01v8_7DPLFP
XXM2 Vp V06 m1_904_n796# Vp Vn sky130_fd_pr__pfet_01v8_MDPZBH
XXM3 Vn m1_904_n796# V06 Vn sky130_fd_pr__nfet_01v8_MYA4RC
C0 Vp Vin 0.113f
C1 m1_904_n796# Vn 0.0382f
C2 m1_904_n796# Vp 0.197f
C3 Vn Vp 0.0214f
C4 m1_904_n796# V06 0.157f
C5 m1_904_n796# Vin 0.203f
C6 V06 Vn 0.00141f
C7 V06 Vp 0.06f
C8 Vn Vin 0.0188f
C9 Vp 0 1.69f
C10 m1_904_n796# 0 0.495f
C11 V06 0 0.217f
C12 Vn 0 0.286f
C13 Vin 0 0.524f
.ends

