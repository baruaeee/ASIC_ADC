* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : preampF_comm_B                               *
* Netlisted  : Tue Dec  3 03:50:38 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733194226940                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733194226940 1 2 3
** N=9 EP=3 FDC=1
M0 1 3 2 2 pfet_01v8 L=1.05e-06 W=5.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733194226940

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733194226941                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733194226941 1 2 3
** N=11 EP=3 FDC=1
M0 1 3 2 2 nfet_01v8 L=1.5e-07 W=1.02e-06 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733194226941

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: preampF_comm_B                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt preampF_comm_B A VDD VSS Y
** N=5 EP=4 FDC=2
X2 VSS Y A pfet_01v8_CDNS_733194226940 $T=130 1720 0 270 $X=-50 $Y=225
X3 VDD Y A nfet_01v8_CDNS_733194226941 $T=485 2750 1 180 $X=-70 $Y=2600
.ends preampF_comm_B
