magic
tech sky130A
magscale 1 2
timestamp 1706454272
<< error_p >>
rect -29 322 29 328
rect -29 288 -17 322
rect -29 282 29 288
rect -29 -288 29 -282
rect -29 -322 -17 -288
rect -29 -328 29 -322
<< pwell >>
rect -211 -460 157 460
<< nmos >>
rect -15 -250 15 250
<< ndiff >>
rect -73 238 -15 250
rect -73 -238 -61 238
rect -27 -238 -15 238
rect -73 -250 -15 -238
rect 15 238 73 250
rect 15 -238 27 238
rect 61 -238 73 238
rect 15 -250 73 -238
<< ndiffc >>
rect -61 -238 -27 238
rect 27 -238 61 238
<< psubdiff >>
rect -141 -424 -79 -390
rect 79 -424 141 -390
<< psubdiffcont >>
rect -79 -424 79 -390
<< poly >>
rect -33 322 33 338
rect -33 288 -17 322
rect 17 288 33 322
rect -33 272 33 288
rect -15 250 15 272
rect -15 -272 15 -250
rect -33 -288 33 -272
rect -33 -322 -17 -288
rect 17 -322 33 -288
rect -33 -338 33 -322
<< polycont >>
rect -17 288 17 322
rect -17 -322 17 -288
<< locali >>
rect -33 288 -17 322
rect 17 288 33 322
rect -61 238 -27 254
rect -61 -254 -27 -238
rect 27 238 61 254
rect 27 -254 61 -238
rect -33 -322 -17 -288
rect 17 -322 33 -288
rect -141 -424 -79 -390
rect 79 -424 141 -390
<< viali >>
rect -17 288 17 322
rect -61 -238 -27 238
rect 27 -238 61 238
rect -17 -322 17 -288
<< metal1 >>
rect -29 322 29 328
rect -29 288 -17 322
rect 17 288 29 322
rect -29 282 29 288
rect -67 238 -21 250
rect -67 -238 -61 238
rect -27 -238 -21 238
rect -67 -250 -21 -238
rect 21 238 67 250
rect 21 -238 27 238
rect 61 -238 67 238
rect 21 -250 67 -238
rect -29 -288 29 -282
rect -29 -322 -17 -288
rect 17 -322 29 -288
rect -29 -328 29 -322
<< properties >>
string FIXED_BBOX -158 -407 158 407
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
