* NGSPICE file created from Analog.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_D7Y3TR a_n63_n101# a_n33_n75# a_n249_n145# a_63_n75#
+ a_n125_n75#
X0 a_63_n75# a_n63_n101# a_n33_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.233 pd=2.12 as=0.124 ps=1.08 w=0.75 l=0.15
X1 a_n33_n75# a_n63_n101# a_n125_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.08 as=0.233 ps=2.12 w=0.75 l=0.15
C0 a_n33_n75# a_63_n75# 0.113f
C1 a_n63_n101# a_n125_n75# 0.00451f
C2 a_63_n75# a_n63_n101# 0.0104f
C3 a_n33_n75# a_n125_n75# 0.113f
C4 a_n33_n75# a_n63_n101# 0.0186f
C5 a_63_n75# a_n249_n145# 0.0963f
C6 a_n33_n75# a_n249_n145# 0.0361f
C7 a_n125_n75# a_n249_n145# 0.105f
C8 a_n63_n101# a_n249_n145# 0.294f
.ends

.subckt sky130_fd_pr__pfet_01v8_2ZD99F w_n349_n261# a_n153_n139# a_n211_n42# a_153_n42#
+ VSUBS
X0 a_153_n42# a_n153_n139# a_n211_n42# w_n349_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.53
C0 a_n211_n42# a_153_n42# 0.0169f
C1 w_n349_n261# a_n153_n139# 0.388f
C2 a_153_n42# a_n153_n139# 0.0177f
C3 a_153_n42# w_n349_n261# 0.0179f
C4 a_n211_n42# a_n153_n139# 0.0177f
C5 a_n211_n42# w_n349_n261# 0.034f
C6 a_153_n42# VSUBS 0.0558f
C7 a_n211_n42# VSUBS 0.0456f
C8 a_n153_n139# VSUBS 0.556f
C9 w_n349_n261# VSUBS 1.16f
.ends

.subckt sky130_fd_pr__nfet_01v8_2BW22M a_154_n42# a_n154_n130# a_n314_n182# a_n212_n42#
X0 a_154_n42# a_n154_n130# a_n212_n42# a_n314_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.54
C0 a_n154_n130# a_n212_n42# 0.0178f
C1 a_154_n42# a_n212_n42# 0.0169f
C2 a_154_n42# a_n154_n130# 0.0178f
C3 a_154_n42# a_n314_n182# 0.0737f
C4 a_n212_n42# a_n314_n182# 0.0816f
C5 a_n154_n130# a_n314_n182# 0.924f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJP3BL a_15_n150# w_n211_n369# a_n73_n150# a_n33_n247#
+ VSUBS
X0 a_15_n150# a_n33_n247# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.15
C0 a_n73_n150# a_15_n150# 0.242f
C1 w_n211_n369# a_n33_n247# 0.19f
C2 a_15_n150# a_n33_n247# 0.0267f
C3 a_n73_n150# a_n33_n247# 0.0267f
C4 a_15_n150# w_n211_n369# 0.0292f
C5 a_n73_n150# w_n211_n369# 0.0292f
C6 a_15_n150# VSUBS 0.126f
C7 a_n73_n150# VSUBS 0.126f
C8 a_n33_n247# VSUBS 0.146f
C9 w_n211_n369# VSUBS 1.02f
.ends

.subckt sky130_fd_pr__nfet_01v8_LH5FDA a_n150_n130# a_276_n182# a_n208_n42# a_150_n42#
X0 a_150_n42# a_n150_n130# a_n208_n42# a_276_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.5
C0 a_n150_n130# a_n208_n42# 0.0176f
C1 a_150_n42# a_n208_n42# 0.0172f
C2 a_150_n42# a_n150_n130# 0.0176f
C3 a_150_n42# a_276_n182# 0.0815f
C4 a_n208_n42# a_276_n182# 0.0736f
C5 a_n150_n130# a_276_n182# 0.904f
.ends

.subckt th02 Vin V02 Vp m1_983_133# m1_571_144# Vn
XXM0 Vin Vn Vn m1_983_133# m1_983_133# sky130_fd_pr__nfet_01v8_D7Y3TR
XXM1 Vp Vin m1_571_144# m1_983_133# Vn sky130_fd_pr__pfet_01v8_2ZD99F
XXM2 m1_571_144# Vp Vn Vp sky130_fd_pr__nfet_01v8_2BW22M
XXM3 V02 Vp Vp m1_983_133# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_983_133# Vn V02 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 V02 Vn 0.00239f
C1 m1_571_144# Vp 0.176f
C2 m1_983_133# m1_571_144# 0.0183f
C3 Vin Vp 0.25f
C4 m1_983_133# Vin 0.279f
C5 V02 m1_571_144# 0.011f
C6 V02 Vin 0.00845f
C7 Vn m1_571_144# 0.00115f
C8 m1_983_133# Vp 0.366f
C9 Vn Vin 0.0263f
C10 V02 Vp 0.118f
C11 m1_983_133# V02 0.155f
C12 Vn Vp 0.0235f
C13 m1_983_133# Vn 0.216f
C14 Vin m1_571_144# 0.332f
C15 Vn 0 0.263f
C16 V02 0 0.334f
C17 m1_983_133# 0 1.44f
C18 Vp 0 3.16f
C19 m1_571_144# 0 0.252f
C20 Vin 0 0.949f
.ends

.subckt sky130_fd_pr__nfet_01v8_2V6S9N a_n216_n42# a_158_n42# a_n158_n130# a_n284_n216#
X0 a_158_n42# a_n158_n130# a_n216_n42# a_n284_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.58
C0 a_158_n42# a_n158_n130# 0.018f
C1 a_n158_n130# a_n216_n42# 0.018f
C2 a_158_n42# a_n216_n42# 0.0165f
C3 a_158_n42# a_n284_n216# 0.0746f
C4 a_n216_n42# a_n284_n216# 0.0746f
C5 a_n158_n130# a_n284_n216# 0.981f
.ends

.subckt sky130_fd_pr__pfet_01v8_XYZSMQ a_n33_n255# a_15_n158# w_n211_n377# a_n73_n158#
+ VSUBS
X0 a_15_n158# a_n33_n255# a_n73_n158# w_n211_n377# sky130_fd_pr__pfet_01v8 ad=0.458 pd=3.74 as=0.458 ps=3.74 w=1.58 l=0.15
C0 a_15_n158# w_n211_n377# 0.0299f
C1 a_n73_n158# w_n211_n377# 0.0299f
C2 a_15_n158# a_n73_n158# 0.254f
C3 w_n211_n377# a_n33_n255# 0.191f
C4 a_15_n158# a_n33_n255# 0.0271f
C5 a_n73_n158# a_n33_n255# 0.0271f
C6 a_15_n158# VSUBS 0.132f
C7 a_n73_n158# VSUBS 0.132f
C8 a_n33_n255# VSUBS 0.146f
C9 w_n211_n377# VSUBS 1.04f
.ends

.subckt sky130_fd_pr__pfet_01v8_AZD9DW w_n353_n261# a_n157_n139# a_n215_n42# a_157_n42#
+ VSUBS
X0 a_157_n42# a_n157_n139# a_n215_n42# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.57
C0 a_157_n42# w_n353_n261# 0.0323f
C1 a_n215_n42# w_n353_n261# 0.0179f
C2 a_157_n42# a_n215_n42# 0.0166f
C3 w_n353_n261# a_n157_n139# 0.396f
C4 a_157_n42# a_n157_n139# 0.0179f
C5 a_n215_n42# a_n157_n139# 0.0179f
C6 a_157_n42# VSUBS 0.0468f
C7 a_n215_n42# VSUBS 0.0559f
C8 a_n157_n139# VSUBS 0.569f
C9 w_n353_n261# VSUBS 1.17f
.ends

.subckt sky130_fd_pr__nfet_01v8_T8HSQ7 a_n175_n297# a_15_n157# a_n33_n245# a_n73_n157#
X0 a_15_n157# a_n33_n245# a_n73_n157# a_n175_n297# sky130_fd_pr__nfet_01v8 ad=0.455 pd=3.72 as=0.455 ps=3.72 w=1.57 l=0.15
C0 a_15_n157# a_n33_n245# 0.0289f
C1 a_n33_n245# a_n73_n157# 0.0289f
C2 a_15_n157# a_n73_n157# 0.253f
C3 a_15_n157# a_n175_n297# 0.161f
C4 a_n73_n157# a_n175_n297# 0.188f
C5 a_n33_n245# a_n175_n297# 0.322f
.ends

.subckt th09 V09 Vin Vn m1_485_n505# Vp m1_962_372#
XXM0 m1_485_n505# Vn Vin Vn sky130_fd_pr__nfet_01v8_2V6S9N
XXM1 Vin m1_485_n505# Vp Vp Vn sky130_fd_pr__pfet_01v8_XYZSMQ
XXM2 Vp m1_485_n505# Vp m1_962_372# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM3 Vp m1_485_n505# V09 m1_962_372# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM4 Vn V09 m1_485_n505# Vn sky130_fd_pr__nfet_01v8_T8HSQ7
C0 m1_962_372# Vn 6.71e-21
C1 V09 Vn 0.00364f
C2 m1_485_n505# m1_962_372# 0.0822f
C3 m1_962_372# Vp 0.0579f
C4 V09 m1_485_n505# 0.104f
C5 V09 Vp 0.0743f
C6 m1_962_372# Vin 0.00821f
C7 m1_485_n505# Vn 0.0846f
C8 Vn Vp 0.0176f
C9 V09 Vin 2.77e-19
C10 m1_485_n505# Vp 0.372f
C11 V09 m1_962_372# 0.00205f
C12 Vn Vin 0.0386f
C13 m1_485_n505# Vin 0.372f
C14 Vin Vp 0.187f
C15 Vin 0 1.1f
C16 m1_485_n505# 0 1.18f
C17 V09 0 0.27f
C18 Vn 0 0.344f
C19 Vp 0 3.27f
C20 m1_962_372# 0 0.118f
.ends

.subckt sky130_fd_pr__pfet_01v8_HPNF99 a_n33_n147# a_23_n50# a_n81_n50# w_n219_n269#
+ VSUBS
X0 a_23_n50# a_n33_n147# a_n81_n50# w_n219_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.23
C0 a_n81_n50# a_n33_n147# 0.00814f
C1 w_n219_n269# a_n33_n147# 0.173f
C2 w_n219_n269# a_n81_n50# 0.0419f
C3 a_n33_n147# a_23_n50# 0.00814f
C4 a_n81_n50# a_23_n50# 0.07f
C5 w_n219_n269# a_23_n50# 0.0185f
C6 a_23_n50# VSUBS 0.0578f
C7 a_n81_n50# VSUBS 0.0428f
C8 a_n33_n147# VSUBS 0.157f
C9 w_n219_n269# VSUBS 0.779f
.ends

.subckt sky130_fd_pr__nfet_01v8_JZU22M a_n213_n42# a_155_n42# a_n155_n130# a_281_n238#
X0 a_155_n42# a_n155_n130# a_n213_n42# a_281_n238# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.55
C0 a_155_n42# a_n213_n42# 0.0168f
C1 a_n155_n130# a_n213_n42# 0.0178f
C2 a_n155_n130# a_155_n42# 0.0178f
C3 a_155_n42# a_281_n238# 0.0816f
C4 a_n213_n42# a_281_n238# 0.0737f
C5 a_n155_n130# a_281_n238# 0.928f
.ends

.subckt sky130_fd_pr__pfet_01v8_TM5S5A a_n80_n147# a_n138_n50# a_80_n50# w_n276_n269#
+ VSUBS
X0 a_80_n50# a_n80_n147# a_n138_n50# w_n276_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.8
C0 a_n138_n50# a_n80_n147# 0.0141f
C1 w_n276_n269# a_n80_n147# 0.297f
C2 w_n276_n269# a_n138_n50# 0.0231f
C3 a_n80_n147# a_80_n50# 0.0141f
C4 a_n138_n50# a_80_n50# 0.0335f
C5 w_n276_n269# a_80_n50# 0.0231f
C6 a_80_n50# VSUBS 0.0565f
C7 a_n138_n50# VSUBS 0.0565f
C8 a_n80_n147# VSUBS 0.296f
C9 w_n276_n269# VSUBS 1.01f
.ends

.subckt sky130_fd_pr__pfet_01v8_AM8GZ5 w_n526_n261# a_n330_n139# a_330_n42# a_n388_n42#
+ VSUBS
X0 a_330_n42# a_n330_n139# a_n388_n42# w_n526_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.3
C0 a_n388_n42# a_n330_n139# 0.0223f
C1 w_n526_n261# a_n330_n139# 0.719f
C2 w_n526_n261# a_n388_n42# 0.0179f
C3 a_n330_n139# a_330_n42# 0.0223f
C4 a_n388_n42# a_330_n42# 0.00853f
C5 w_n526_n261# a_330_n42# 0.0408f
C6 a_330_n42# VSUBS 0.0435f
C7 a_n388_n42# VSUBS 0.0585f
C8 a_n330_n139# VSUBS 1.13f
C9 w_n526_n261# VSUBS 1.76f
.ends

.subckt sky130_fd_pr__nfet_01v8_H7HSAV a_n73_n250# a_15_n250# a_n33_n338# a_n141_n424#
X0 a_15_n250# a_n33_n338# a_n73_n250# a_n141_n424# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.15
C0 a_15_n250# a_n73_n250# 0.401f
C1 a_n33_n338# a_n73_n250# 0.0337f
C2 a_n33_n338# a_15_n250# 0.0337f
C3 a_15_n250# a_n141_n424# 0.24f
C4 a_n73_n250# a_n141_n424# 0.24f
C5 a_n33_n338# a_n141_n424# 0.327f
.ends

.subckt th14 V14 Vin Vn m1_641_n318# Vp m1_891_419#
XXM0 Vn Vn m1_641_n318# Vp Vn sky130_fd_pr__pfet_01v8_HPNF99
XXM1 m1_641_n318# m1_891_419# Vin Vn sky130_fd_pr__nfet_01v8_JZU22M
XXM2 Vin Vp m1_891_419# Vp Vn sky130_fd_pr__pfet_01v8_TM5S5A
XXM3 Vp m1_891_419# V14 Vp Vn sky130_fd_pr__pfet_01v8_AM8GZ5
XXM4 Vn V14 m1_891_419# Vn sky130_fd_pr__nfet_01v8_H7HSAV
C0 Vp V14 0.082f
C1 Vin m1_641_n318# 0.229f
C2 Vin m1_891_419# 0.132f
C3 m1_891_419# m1_641_n318# 0.00289f
C4 Vin V14 0.00516f
C5 m1_891_419# V14 0.249f
C6 Vin Vp 0.201f
C7 Vp m1_641_n318# 0.0629f
C8 Vp m1_891_419# 0.227f
C9 m1_891_419# Vn 1.7f
C10 V14 Vn 0.273f
C11 Vp Vn 3.39f
C12 Vin Vn 1.76f
C13 m1_641_n318# Vn 0.313f
.ends

.subckt sky130_fd_pr__nfet_01v8_VGVEGU a_n142_n216# a_n74_n42# a_n33_n130# a_16_n42#
X0 a_16_n42# a_n33_n130# a_n74_n42# a_n142_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.16
C0 a_n74_n42# a_n33_n130# 0.0191f
C1 a_16_n42# a_n74_n42# 0.0684f
C2 a_16_n42# a_n33_n130# 0.0191f
C3 a_16_n42# a_n142_n216# 0.0652f
C4 a_n74_n42# a_n142_n216# 0.0652f
C5 a_n33_n130# a_n142_n216# 0.317f
.ends

.subckt sky130_fd_pr__pfet_01v8_EDPLE3 a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n33_n139# w_n211_n261# 0.187f
C1 a_n73_n42# a_15_n42# 0.0699f
C2 a_n33_n139# a_15_n42# 0.0192f
C3 a_n73_n42# a_n33_n139# 0.0192f
C4 w_n211_n261# a_15_n42# 0.0197f
C5 a_n73_n42# w_n211_n261# 0.0197f
C6 a_15_n42# VSUBS 0.0445f
C7 a_n73_n42# VSUBS 0.0445f
C8 a_n33_n139# VSUBS 0.143f
C9 w_n211_n261# VSUBS 0.749f
.ends

.subckt sky130_fd_pr__pfet_01v8_JM8GTH a_50_n42# w_n246_n261# a_n50_n139# a_n108_n42#
+ VSUBS
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 a_n50_n139# w_n246_n261# 0.223f
C1 a_n108_n42# a_50_n42# 0.0391f
C2 a_n50_n139# a_50_n42# 0.00909f
C3 a_n108_n42# a_n50_n139# 0.00909f
C4 w_n246_n261# a_50_n42# 0.0224f
C5 a_n108_n42# w_n246_n261# 0.0224f
C6 a_50_n42# VSUBS 0.0488f
C7 a_n108_n42# VSUBS 0.0488f
C8 a_n50_n139# VSUBS 0.209f
C9 w_n246_n261# VSUBS 0.88f
.ends

.subckt sky130_fd_pr__nfet_01v8_MYA4RC a_n73_n46# a_n33_n134# a_15_n46# a_n175_n186#
X0 a_15_n46# a_n33_n134# a_n73_n46# a_n175_n186# sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.5 as=0.133 ps=1.5 w=0.46 l=0.15
C0 a_n73_n46# a_n33_n134# 0.0212f
C1 a_15_n46# a_n73_n46# 0.0763f
C2 a_15_n46# a_n33_n134# 0.0212f
C3 a_15_n46# a_n175_n186# 0.0671f
C4 a_n73_n46# a_n175_n186# 0.0756f
C5 a_n33_n134# a_n175_n186# 0.314f
.ends

.subckt th07 Vin V07 Vp m1_808_n892# Vn
XXM0 Vn m1_808_n892# Vin Vn sky130_fd_pr__nfet_01v8_VGVEGU
XXM1 m1_808_n892# Vp Vin Vp Vn sky130_fd_pr__pfet_01v8_EDPLE3
XXM2 V07 Vp m1_808_n892# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM3 V07 m1_808_n892# Vn Vn sky130_fd_pr__nfet_01v8_MYA4RC
C0 Vin m1_808_n892# 0.365f
C1 Vp V07 0.0569f
C2 Vp m1_808_n892# 0.209f
C3 V07 m1_808_n892# 0.112f
C4 Vp Vin 0.157f
C5 V07 Vin 0.00135f
C6 Vin Vn 0.524f
C7 Vp Vn 1.57f
C8 m1_808_n892# Vn 0.596f
C9 V07 Vn 0.276f
.ends

.subckt sky130_fd_pr__pfet_01v8_P28Q2U a_n33_n232# a_15_n135# w_n211_n354# a_n73_n135#
+ VSUBS
X0 a_15_n135# a_n33_n232# a_n73_n135# w_n211_n354# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.28 as=0.391 ps=3.28 w=1.35 l=0.15
C0 a_n73_n135# a_n33_n232# 0.0258f
C1 a_15_n135# w_n211_n354# 0.0279f
C2 w_n211_n354# a_n33_n232# 0.19f
C3 a_15_n135# a_n33_n232# 0.0258f
C4 a_n73_n135# w_n211_n354# 0.0279f
C5 a_15_n135# a_n73_n135# 0.218f
C6 a_15_n135# VSUBS 0.115f
C7 a_n73_n135# VSUBS 0.115f
C8 a_n33_n232# VSUBS 0.146f
C9 w_n211_n354# VSUBS 0.983f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZMY3VB a_n348_n42# a_n290_n130# a_n450_n182# a_290_n42#
X0 a_290_n42# a_n290_n130# a_n348_n42# a_n450_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.9
C0 a_290_n42# a_n348_n42# 0.00961f
C1 a_n290_n130# a_n348_n42# 0.0217f
C2 a_290_n42# a_n290_n130# 0.0217f
C3 a_290_n42# a_n450_n182# 0.076f
C4 a_n348_n42# a_n450_n182# 0.0839f
C5 a_n290_n130# a_n450_n182# 1.6f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n73_n100# a_n33_n197# 0.0236f
C1 a_15_n100# w_n211_n319# 0.0248f
C2 w_n211_n319# a_n33_n197# 0.189f
C3 a_15_n100# a_n33_n197# 0.0236f
C4 a_n73_n100# w_n211_n319# 0.0248f
C5 a_15_n100# a_n73_n100# 0.162f
C6 a_15_n100# VSUBS 0.0885f
C7 a_n73_n100# VSUBS 0.0885f
C8 a_n33_n197# VSUBS 0.145f
C9 w_n211_n319# VSUBS 0.894f
.ends

.subckt sky130_fd_pr__pfet_01v8_WV9GCW a_n158_n42# w_n296_n261# a_n100_n139# a_100_n42#
+ VSUBS
X0 a_100_n42# a_n100_n139# a_n158_n42# w_n296_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1
C0 a_n158_n42# a_n100_n139# 0.0144f
C1 a_100_n42# w_n296_n261# 0.0224f
C2 w_n296_n261# a_n100_n139# 0.346f
C3 a_100_n42# a_n100_n139# 0.0144f
C4 a_n158_n42# w_n296_n261# 0.0224f
C5 a_100_n42# a_n158_n42# 0.024f
C6 a_100_n42# VSUBS 0.0504f
C7 a_n158_n42# VSUBS 0.0504f
C8 a_n100_n139# VSUBS 0.353f
C9 w_n296_n261# VSUBS 1.06f
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n141_240# a_n33_n188# a_15_n100#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n141_240# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_15_n100# a_n73_n100# 0.162f
C1 a_n33_n188# a_n73_n100# 0.0254f
C2 a_15_n100# a_n33_n188# 0.0254f
C3 a_15_n100# a_n141_240# 0.113f
C4 a_n73_n100# a_n141_240# 0.113f
C5 a_n33_n188# a_n141_240# 0.322f
.ends

.subckt th12 Vp V12 Vin m1_529_n42# m1_394_n856# Vn
XXM0 Vn Vn Vp m1_394_n856# Vn sky130_fd_pr__pfet_01v8_P28Q2U
XXM1 m1_529_n42# Vin Vn m1_394_n856# sky130_fd_pr__nfet_01v8_ZMY3VB
XXM2 m1_529_n42# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM3 Vp Vp m1_529_n42# V12 Vn sky130_fd_pr__pfet_01v8_WV9GCW
XXM4 V12 Vn m1_529_n42# Vn sky130_fd_pr__nfet_01v8_648S5X
C0 Vn m1_394_n856# 0.0338f
C1 m1_529_n42# m1_394_n856# 0.0134f
C2 m1_394_n856# V12 4.74e-19
C3 m1_394_n856# Vp 0.04f
C4 Vin m1_394_n856# 0.321f
C5 m1_529_n42# Vn 0.254f
C6 Vn V12 0.0234f
C7 m1_529_n42# V12 0.0929f
C8 Vn Vp 0.132f
C9 m1_529_n42# Vp 0.322f
C10 V12 Vp 0.0454f
C11 Vin Vn 0.135f
C12 Vin m1_529_n42# 0.0965f
C13 Vin V12 0.00205f
C14 Vin Vp 0.238f
C15 Vn 0 0.29f
C16 Vp 0 2.88f
C17 m1_529_n42# 0 0.861f
C18 V12 0 0.359f
C19 Vin 0 1.9f
C20 m1_394_n856# 0 0.215f
.ends

.subckt sky130_fd_pr__nfet_01v8_Q7AWK3 a_n180_n340# a_20_n200# a_n78_n200# a_n33_n288#
X0 a_20_n200# a_n33_n288# a_n78_n200# a_n180_n340# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
C0 a_20_n200# a_n78_n200# 0.288f
C1 a_n33_n288# a_n78_n200# 0.024f
C2 a_n33_n288# a_20_n200# 0.024f
C3 a_20_n200# a_n180_n340# 0.202f
C4 a_n78_n200# a_n180_n340# 0.237f
C5 a_n33_n288# a_n180_n340# 0.325f
.ends

.subckt sky130_fd_pr__pfet_01v8_EXJYQP w_n359_n261# a_n163_n139# a_n221_n42# a_163_n42#
+ VSUBS
X0 a_163_n42# a_n163_n139# a_n221_n42# w_n359_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.63
C0 a_n221_n42# a_n163_n139# 0.0182f
C1 a_163_n42# a_n163_n139# 0.0182f
C2 w_n359_n261# a_n163_n139# 0.413f
C3 a_163_n42# a_n221_n42# 0.0161f
C4 w_n359_n261# a_n221_n42# 0.0179f
C5 a_163_n42# w_n359_n261# 0.0408f
C6 a_163_n42# VSUBS 0.041f
C7 a_n221_n42# VSUBS 0.056f
C8 a_n163_n139# VSUBS 0.584f
C9 w_n359_n261# VSUBS 1.24f
.ends

.subckt sky130_fd_pr__pfet_01v8_HJHF6N a_n170_n50# w_n308_n269# a_n112_n147# a_112_n50#
+ VSUBS
X0 a_112_n50# a_n112_n147# a_n170_n50# w_n308_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1.12
C0 a_n170_n50# a_n112_n147# 0.0172f
C1 a_112_n50# a_n112_n147# 0.0172f
C2 w_n308_n269# a_n112_n147# 0.378f
C3 a_112_n50# a_n170_n50# 0.0259f
C4 w_n308_n269# a_n170_n50# 0.0232f
C5 a_112_n50# w_n308_n269# 0.0232f
C6 a_112_n50# VSUBS 0.0577f
C7 a_n170_n50# VSUBS 0.0577f
C8 a_n112_n147# VSUBS 0.389f
C9 w_n308_n269# VSUBS 1.14f
.ends

.subckt sky130_fd_pr__nfet_01v8_N39H2X a_n76_n100# a_n33_n188# a_18_n100# a_144_n240#
X0 a_18_n100# a_n33_n188# a_n76_n100# a_144_n240# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.18
C0 a_18_n100# a_n76_n100# 0.152f
C1 a_n33_n188# a_n76_n100# 0.0205f
C2 a_n33_n188# a_18_n100# 0.0205f
C3 a_18_n100# a_144_n240# 0.133f
C4 a_n76_n100# a_144_n240# 0.115f
C5 a_n33_n188# a_144_n240# 0.32f
.ends

.subckt th05 Vp V05 Vin m1_752_n794# Vn
XXM0 Vn m1_752_n794# Vn Vin sky130_fd_pr__nfet_01v8_Q7AWK3
XXM1 Vp Vin m1_752_n794# Vp Vn sky130_fd_pr__pfet_01v8_EXJYQP
XXM2 Vp Vp m1_752_n794# V05 Vn sky130_fd_pr__pfet_01v8_HJHF6N
XXM3 Vn m1_752_n794# V05 Vn sky130_fd_pr__nfet_01v8_N39H2X
C0 Vin Vp 0.139f
C1 Vp Vn 0.0115f
C2 Vin m1_752_n794# 0.2f
C3 Vn m1_752_n794# 0.136f
C4 Vin V05 0.00406f
C5 V05 Vn 0.0364f
C6 Vp m1_752_n794# 0.198f
C7 Vp V05 0.0548f
C8 V05 m1_752_n794# 0.0855f
C9 Vin Vn 0.041f
C10 m1_752_n794# 0 0.788f
C11 Vp 0 2.28f
C12 V05 0 0.314f
C13 Vin 0 0.905f
C14 Vn 0 0.547f
.ends

.subckt sky130_fd_pr__nfet_01v8_4L9AWD a_n206_n182# a_n46_n130# a_n104_n42# a_46_n42#
X0 a_46_n42# a_n46_n130# a_n104_n42# a_n206_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.46
C0 a_n46_n130# a_46_n42# 0.00852f
C1 a_n104_n42# a_46_n42# 0.0412f
C2 a_n104_n42# a_n46_n130# 0.00852f
C3 a_46_n42# a_n206_n182# 0.0705f
C4 a_n104_n42# a_n206_n182# 0.0784f
C5 a_n46_n130# a_n206_n182# 0.388f
.ends

.subckt sky130_fd_pr__pfet_01v8_EZD9Q7 w_n224_n261# a_28_n42# a_n33_n139# a_n86_n42#
+ VSUBS
X0 a_28_n42# a_n33_n139# a_n86_n42# w_n224_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.28
C0 a_n86_n42# a_28_n42# 0.0541f
C1 w_n224_n261# a_28_n42# 0.0224f
C2 w_n224_n261# a_n86_n42# 0.0224f
C3 a_n33_n139# a_28_n42# 0.00625f
C4 a_n33_n139# a_n86_n42# 0.00625f
C5 a_n33_n139# w_n224_n261# 0.183f
C6 a_28_n42# VSUBS 0.0479f
C7 a_n86_n42# VSUBS 0.0479f
C8 a_n33_n139# VSUBS 0.155f
C9 w_n224_n261# VSUBS 0.799f
.ends

.subckt sky130_fd_pr__pfet_01v8_M479BZ a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n42# a_15_n42# 0.0699f
C1 w_n211_n261# a_15_n42# 0.0389f
C2 w_n211_n261# a_n73_n42# 0.016f
C3 a_n33_n139# a_15_n42# 0.0192f
C4 a_n33_n139# a_n73_n42# 0.0192f
C5 a_n33_n139# w_n211_n261# 0.182f
C6 a_15_n42# VSUBS 0.0328f
C7 a_n73_n42# VSUBS 0.0478f
C8 a_n33_n139# VSUBS 0.145f
C9 w_n211_n261# VSUBS 0.785f
.ends

.subckt sky130_fd_pr__nfet_01v8_4BNSKG a_n144_n216# a_18_n42# a_n33_n130# a_n76_n42#
X0 a_18_n42# a_n33_n130# a_n76_n42# a_n144_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.18
C0 a_n33_n130# a_18_n42# 0.0154f
C1 a_n76_n42# a_18_n42# 0.0655f
C2 a_n76_n42# a_n33_n130# 0.0154f
C3 a_18_n42# a_n144_n216# 0.0668f
C4 a_n76_n42# a_n144_n216# 0.0668f
C5 a_n33_n130# a_n144_n216# 0.319f
.ends

.subckt th10 Vp V10 Vin Vn m1_502_n495# m1_536_174#
XXM0 m1_502_n495# Vn Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vn Vin m1_536_174# m1_502_n495# sky130_fd_pr__nfet_01v8_4L9AWD
XXM2 Vp m1_536_174# Vin Vp Vn sky130_fd_pr__pfet_01v8_EZD9Q7
XXM3 Vp Vp m1_536_174# V10 Vn sky130_fd_pr__pfet_01v8_M479BZ
XXM4 Vn V10 m1_536_174# Vn sky130_fd_pr__nfet_01v8_4BNSKG
C0 m1_502_n495# Vin 0.0207f
C1 Vin V10 0.0187f
C2 m1_502_n495# Vn 0.0348f
C3 V10 Vn 0.0577f
C4 m1_536_174# Vp 0.172f
C5 m1_502_n495# V10 0.042f
C6 Vin m1_536_174# 0.0971f
C7 m1_536_174# Vn 0.233f
C8 m1_502_n495# m1_536_174# 0.00612f
C9 m1_536_174# V10 0.177f
C10 Vin Vp 0.175f
C11 Vn Vp 0.102f
C12 m1_502_n495# Vp 0.0256f
C13 V10 Vp 0.0702f
C14 Vin Vn 0.114f
C15 Vin 0 0.664f
C16 m1_536_174# 0 0.825f
C17 Vp 0 2.17f
C18 V10 0 0.249f
C19 Vn 0 0.463f
C20 m1_502_n495# 0 0.146f
.ends

.subckt sky130_fd_pr__nfet_01v8_X33H33 a_n73_n110# a_n175_n250# a_n33_n198# a_15_n110#
X0 a_15_n110# a_n33_n198# a_n73_n110# a_n175_n250# sky130_fd_pr__nfet_01v8 ad=0.319 pd=2.78 as=0.319 ps=2.78 w=1.1 l=0.15
C0 a_15_n110# a_n73_n110# 0.178f
C1 a_15_n110# a_n33_n198# 0.0261f
C2 a_n73_n110# a_n33_n198# 0.0261f
C3 a_15_n110# a_n175_n250# 0.121f
C4 a_n73_n110# a_n175_n250# 0.141f
C5 a_n33_n198# a_n175_n250# 0.32f
.ends

.subckt sky130_fd_pr__pfet_01v8_AMA9E4 a_n194_n44# a_n136_n141# w_n332_n263# a_136_n44#
+ VSUBS
X0 a_136_n44# a_n136_n141# a_n194_n44# w_n332_n263# sky130_fd_pr__pfet_01v8 ad=0.128 pd=1.46 as=0.128 ps=1.46 w=0.44 l=1.36
C0 a_n194_n44# a_n136_n141# 0.0174f
C1 a_n194_n44# w_n332_n263# 0.0226f
C2 a_n194_n44# a_136_n44# 0.0196f
C3 a_n136_n141# w_n332_n263# 0.434f
C4 a_n136_n141# a_136_n44# 0.0174f
C5 a_136_n44# w_n332_n263# 0.0226f
C6 a_136_n44# VSUBS 0.0532f
C7 a_n194_n44# VSUBS 0.0532f
C8 a_n136_n141# VSUBS 0.457f
C9 w_n332_n263# VSUBS 1.2f
.ends

.subckt sky130_fd_pr__pfet_01v8_8DZSNJ a_n74_n100# a_16_n100# w_n212_n319# a_n33_n197#
+ VSUBS
X0 a_16_n100# a_n33_n197# a_n74_n100# w_n212_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.16
C0 a_n74_n100# a_n33_n197# 0.0223f
C1 a_n74_n100# w_n212_n319# 0.0252f
C2 a_n74_n100# a_16_n100# 0.159f
C3 a_n33_n197# w_n212_n319# 0.189f
C4 a_n33_n197# a_16_n100# 0.0223f
C5 a_16_n100# w_n212_n319# 0.0252f
C6 a_16_n100# VSUBS 0.089f
C7 a_n74_n100# VSUBS 0.089f
C8 a_n33_n197# VSUBS 0.146f
C9 w_n212_n319# VSUBS 0.899f
.ends

.subckt th03 V03 Vin Vp m1_890_n844# m1_638_n591# Vn
XXM0 Vn Vn Vin m1_890_n844# sky130_fd_pr__nfet_01v8_X33H33
XXM1 m1_638_n591# Vin Vp m1_890_n844# Vn sky130_fd_pr__pfet_01v8_AMA9E4
XXM2 Vp Vn Vp m1_638_n591# sky130_fd_pr__nfet_01v8_LH5FDA
XXM3 Vp V03 Vp m1_890_n844# Vn sky130_fd_pr__pfet_01v8_8DZSNJ
XXM4 m1_890_n844# Vn Vn V03 sky130_fd_pr__nfet_01v8_LH5FDA
C0 Vn m1_890_n844# 0.183f
C1 Vp m1_890_n844# 0.459f
C2 Vin m1_890_n844# 0.188f
C3 m1_638_n591# m1_890_n844# 0.0187f
C4 V03 m1_890_n844# 0.129f
C5 Vp Vn 0.023f
C6 Vn Vin 0.105f
C7 Vp Vin 0.313f
C8 Vn m1_638_n591# 0.0097f
C9 Vp m1_638_n591# 0.169f
C10 Vin m1_638_n591# 0.0439f
C11 V03 Vn 0.0337f
C12 V03 Vp 0.0492f
C13 V03 Vin 0.0036f
C14 Vp 0 3.07f
C15 V03 0 0.308f
C16 Vn 0 0.446f
C17 m1_890_n844# 0 1.05f
C18 m1_638_n591# 0 0.224f
C19 Vin 0 0.924f
.ends

.subckt sky130_fd_pr__nfet_01v8_SHU4BF a_n73_n353# a_n141_493# a_15_n353# a_n33_n441#
X0 a_15_n353# a_n33_n441# a_n73_n353# a_n141_493# sky130_fd_pr__nfet_01v8 ad=1.02 pd=7.64 as=1.02 ps=7.64 w=3.53 l=0.15
C0 a_n33_n441# a_15_n353# 0.0384f
C1 a_n73_n353# a_15_n353# 0.564f
C2 a_n73_n353# a_n33_n441# 0.0384f
C3 a_15_n353# a_n141_493# 0.327f
C4 a_n73_n353# a_n141_493# 0.327f
C5 a_n33_n441# a_n141_493# 0.329f
.ends

.subckt sky130_fd_pr__pfet_01v8_HE9GT9 a_n408_n42# a_350_n42# w_n546_n261# a_n350_n139#
+ VSUBS
X0 a_350_n42# a_n350_n139# a_n408_n42# w_n546_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 w_n546_n261# a_n408_n42# 0.0408f
C1 a_n350_n139# a_n408_n42# 0.0226f
C2 a_n350_n139# w_n546_n261# 0.756f
C3 a_350_n42# a_n408_n42# 0.00807f
C4 a_350_n42# w_n546_n261# 0.0179f
C5 a_n350_n139# a_350_n42# 0.0226f
C6 a_350_n42# VSUBS 0.0587f
C7 a_n408_n42# VSUBS 0.0437f
C8 a_n350_n139# VSUBS 1.19f
C9 w_n546_n261# VSUBS 1.83f
.ends

.subckt sky130_fd_pr__nfet_01v8_LHD8GA a_n408_n42# a_350_n42# a_n350_n130# a_n510_n182#
X0 a_350_n42# a_n350_n130# a_n408_n42# a_n510_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 a_n350_n130# a_350_n42# 0.0226f
C1 a_n408_n42# a_350_n42# 0.00807f
C2 a_n408_n42# a_n350_n130# 0.0226f
C3 a_350_n42# a_n510_n182# 0.0766f
C4 a_n408_n42# a_n510_n182# 0.0845f
C5 a_n350_n130# a_n510_n182# 1.9f
.ends

.subckt th01 Vp Vin V01 m1_991_n1219# Vn m1_571_n501#
XXM0 Vn Vn m1_991_n1219# Vin sky130_fd_pr__nfet_01v8_SHU4BF
XXM1 m1_571_n501# m1_991_n1219# Vp Vin Vn sky130_fd_pr__pfet_01v8_HE9GT9
XXM2 Vp m1_571_n501# Vp Vn sky130_fd_pr__nfet_01v8_LHD8GA
XXM3 Vp Vp V01 m1_991_n1219# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_991_n1219# Vn V01 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 Vin Vn 0.0582f
C1 V01 Vn 0.0149f
C2 Vin m1_571_n501# 0.274f
C3 Vin m1_991_n1219# 0.208f
C4 V01 m1_571_n501# 2.16e-20
C5 V01 m1_991_n1219# 0.0901f
C6 Vn m1_571_n501# 2.57e-20
C7 m1_991_n1219# Vn 0.0569f
C8 Vp Vin 0.354f
C9 m1_991_n1219# m1_571_n501# 0.0899f
C10 Vp V01 0.0684f
C11 Vp Vn 0.0233f
C12 Vp m1_571_n501# 0.32f
C13 Vp m1_991_n1219# 0.423f
C14 Vin V01 0.00412f
C15 Vn 0 0.633f
C16 m1_991_n1219# 0 1.24f
C17 V01 0 0.373f
C18 Vp 0 4.41f
C19 m1_571_n501# 0 0.194f
C20 Vin 0 1.87f
.ends

.subckt sky130_fd_pr__pfet_01v8_MWHFPY a_n73_n63# a_n33_n160# w_n211_n282# a_15_n63#
+ VSUBS
X0 a_15_n63# a_n33_n160# a_n73_n63# w_n211_n282# sky130_fd_pr__pfet_01v8 ad=0.183 pd=1.84 as=0.183 ps=1.84 w=0.63 l=0.15
C0 w_n211_n282# a_15_n63# 0.0591f
C1 a_n33_n160# a_15_n63# 0.021f
C2 a_n73_n63# a_15_n63# 0.103f
C3 a_n33_n160# w_n211_n282# 0.237f
C4 w_n211_n282# a_n73_n63# 0.0591f
C5 a_n33_n160# a_n73_n63# 0.021f
C6 a_15_n63# VSUBS 0.0348f
C7 a_n73_n63# VSUBS 0.0348f
C8 a_n33_n160# VSUBS 0.116f
C9 w_n211_n282# VSUBS 1.1f
.ends

.subckt sky130_fd_pr__nfet_01v8_DPSGWY a_350_n100# a_n408_n100# a_n350_n188# a_n510_n274#
X0 a_350_n100# a_n350_n188# a_n408_n100# a_n510_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3.5
C0 a_n408_n100# a_n350_n188# 0.0439f
C1 a_n350_n188# a_350_n100# 0.0439f
C2 a_n408_n100# a_350_n100# 0.0188f
C3 a_350_n100# a_n510_n274# 0.159f
C4 a_n408_n100# a_n510_n274# 0.159f
C5 a_n350_n188# a_n510_n274# 2.13f
.ends

.subckt preamp Vp Vin Vpamp Vn
XXM0 Vn Vin Vp Vpamp Vn sky130_fd_pr__pfet_01v8_MWHFPY
XXM1 Vpamp Vp Vin Vn sky130_fd_pr__nfet_01v8_DPSGWY
C0 Vn Vp 0.297f
C1 Vin Vp 0.324f
C2 Vn Vpamp 0.047f
C3 Vin Vpamp 0.0777f
C4 Vin Vn 0.29f
C5 Vpamp Vp 0.0552f
C6 Vn 0 0.193f
C7 Vpamp 0 0.444f
C8 Vp 0 1.53f
C9 Vin 0 2.21f
.ends

.subckt sky130_fd_pr__pfet_01v8_LDQF7K a_n33_n147# a_29_n50# a_n87_n50# w_n225_n269#
+ VSUBS
X0 a_29_n50# a_n33_n147# a_n87_n50# w_n225_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.29
C0 a_n87_n50# a_29_n50# 0.0628f
C1 a_n87_n50# w_n225_n269# 0.0457f
C2 a_n33_n147# a_29_n50# 0.00691f
C3 a_n33_n147# w_n225_n269# 0.176f
C4 a_n33_n147# a_n87_n50# 0.00691f
C5 a_29_n50# w_n225_n269# 0.0186f
C6 a_29_n50# VSUBS 0.0581f
C7 a_n87_n50# VSUBS 0.0403f
C8 a_n33_n147# VSUBS 0.158f
C9 w_n225_n269# VSUBS 0.854f
.ends

.subckt sky130_fd_pr__nfet_01v8_HZA4VB a_326_n230# a_n200_n130# a_200_n42# li_n360_158#
+ a_n258_n42#
X0 a_200_n42# a_n200_n130# a_n258_n42# a_326_n230# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_200_n42# a_n200_n130# 0.0196f
C1 a_n258_n42# a_n200_n130# 0.0196f
C2 a_n258_n42# a_200_n42# 0.0134f
C3 li_n360_158# a_326_n230# 0.0244f
C4 a_200_n42# a_326_n230# 0.0748f
C5 a_n258_n42# a_326_n230# 0.0746f
C6 a_n200_n130# a_326_n230# 1.15f
.ends

.subckt sky130_fd_pr__pfet_01v8_GEY2B5 w_n275_n270# a_n137_n51# a_79_n51# a_n79_n148#
+ VSUBS
X0 a_79_n51# a_n79_n148# a_n137_n51# w_n275_n270# sky130_fd_pr__pfet_01v8 ad=0.148 pd=1.6 as=0.148 ps=1.6 w=0.51 l=0.79
C0 a_n137_n51# a_79_n51# 0.0345f
C1 a_n137_n51# w_n275_n270# 0.0232f
C2 a_n79_n148# a_79_n51# 0.0141f
C3 a_n79_n148# w_n275_n270# 0.294f
C4 a_n79_n148# a_n137_n51# 0.0141f
C5 a_79_n51# w_n275_n270# 0.0232f
C6 a_79_n51# VSUBS 0.0573f
C7 a_n137_n51# VSUBS 0.0573f
C8 a_n79_n148# VSUBS 0.294f
C9 w_n275_n270# VSUBS 1.01f
.ends

.subckt sky130_fd_pr__pfet_01v8_KQKFM4 w_n526_n261# a_n330_n139# a_330_n42# a_n388_n42#
+ VSUBS
X0 a_330_n42# a_n330_n139# a_n388_n42# w_n526_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.3
C0 a_n388_n42# a_330_n42# 0.00853f
C1 a_n388_n42# w_n526_n261# 0.0224f
C2 a_n330_n139# a_330_n42# 0.0223f
C3 a_n330_n139# w_n526_n261# 0.911f
C4 a_n330_n139# a_n388_n42# 0.0223f
C5 a_330_n42# w_n526_n261# 0.0224f
C6 a_330_n42# VSUBS 0.0545f
C7 a_n388_n42# VSUBS 0.0545f
C8 a_n330_n139# VSUBS 1.02f
C9 w_n526_n261# VSUBS 1.89f
.ends

.subckt sky130_fd_pr__nfet_01v8_5NW376 a_n73_n251# a_n141_391# a_15_n251# a_n33_n339#
X0 a_15_n251# a_n33_n339# a_n73_n251# a_n141_391# sky130_fd_pr__nfet_01v8 ad=0.728 pd=5.6 as=0.728 ps=5.6 w=2.51 l=0.15
C0 a_15_n251# a_n33_n339# 0.0337f
C1 a_n73_n251# a_n33_n339# 0.0337f
C2 a_n73_n251# a_15_n251# 0.402f
C3 a_15_n251# a_n141_391# 0.241f
C4 a_n73_n251# a_n141_391# 0.241f
C5 a_n33_n339# a_n141_391# 0.327f
.ends

.subckt th15 V15 Vin m1_597_n912# Vp m1_849_n157# Vn
XXM0 Vn Vn m1_597_n912# Vp Vn sky130_fd_pr__pfet_01v8_LDQF7K
XXM1 Vn Vin m1_849_n157# Vn m1_597_n912# sky130_fd_pr__nfet_01v8_HZA4VB
XXM2 Vp Vp m1_849_n157# Vin Vn sky130_fd_pr__pfet_01v8_GEY2B5
XXM3 Vp m1_849_n157# V15 Vp Vn sky130_fd_pr__pfet_01v8_KQKFM4
XXM4 Vn Vn V15 m1_849_n157# sky130_fd_pr__nfet_01v8_5NW376
C0 Vn Vin 0.38f
C1 V15 Vp 0.0762f
C2 m1_597_n912# Vn 0.175f
C3 V15 m1_849_n157# 0.202f
C4 Vp Vn 0.0678f
C5 m1_849_n157# Vn 0.171f
C6 V15 Vn 2.72e-19
C7 m1_597_n912# Vin 0.211f
C8 Vp Vin 0.166f
C9 m1_849_n157# Vin 0.0977f
C10 Vp m1_597_n912# 0.0557f
C11 V15 Vin 0.00573f
C12 m1_597_n912# m1_849_n157# 0.00715f
C13 Vp m1_849_n157# 0.226f
C14 V15 0 0.332f
C15 Vn 0 0.276f
C16 m1_849_n157# 0 1.28f
C17 Vp 0 3.52f
C18 Vin 0 1.58f
C19 m1_597_n912# 0 0.19f
.ends

.subckt sky130_fd_pr__nfet_01v8_JSJ4VK a_113_n42# a_n239_n216# a_n171_n42# a_n113_n130#
X0 a_113_n42# a_n113_n130# a_n171_n42# a_n239_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.13
C0 a_n171_n42# a_113_n42# 0.0218f
C1 a_n113_n130# a_113_n42# 0.0154f
C2 a_n113_n130# a_n171_n42# 0.0154f
C3 a_113_n42# a_n239_n216# 0.0734f
C4 a_n171_n42# a_n239_n216# 0.0734f
C5 a_n113_n130# a_n239_n216# 0.746f
.ends

.subckt sky130_fd_pr__pfet_01v8_EVXEQ2 a_16_n67# a_n33_n164# a_n74_n67# w_n212_n286#
+ VSUBS
X0 a_16_n67# a_n33_n164# a_n74_n67# w_n212_n286# sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.92 as=0.194 ps=1.92 w=0.67 l=0.16
C0 a_n33_n164# a_n74_n67# 0.0198f
C1 w_n212_n286# a_n74_n67# 0.0184f
C2 a_n33_n164# a_16_n67# 0.0198f
C3 w_n212_n286# a_16_n67# 0.0544f
C4 a_16_n67# a_n74_n67# 0.107f
C5 w_n212_n286# a_n33_n164# 0.183f
C6 a_16_n67# VSUBS 0.0435f
C7 a_n74_n67# VSUBS 0.0673f
C8 a_n33_n164# VSUBS 0.147f
C9 w_n212_n286# VSUBS 0.864f
.ends

.subckt sky130_fd_pr__pfet_01v8_BBE9QE w_n244_n262# a_n106_n43# a_48_n43# a_n48_n140#
+ VSUBS
X0 a_48_n43# a_n48_n140# a_n106_n43# w_n244_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.48
C0 a_n48_n140# a_n106_n43# 0.00893f
C1 w_n244_n262# a_n106_n43# 0.0225f
C2 a_n48_n140# a_48_n43# 0.00893f
C3 w_n244_n262# a_48_n43# 0.0225f
C4 a_48_n43# a_n106_n43# 0.041f
C5 w_n244_n262# a_n48_n140# 0.218f
C6 a_48_n43# VSUBS 0.0495f
C7 a_n106_n43# VSUBS 0.0495f
C8 a_n48_n140# VSUBS 0.203f
C9 w_n244_n262# VSUBS 0.876f
.ends

.subckt sky130_fd_pr__nfet_01v8_NCP4B2 a_n73_n47# a_n141_n221# a_n33_n135# a_15_n47#
X0 a_15_n47# a_n33_n135# a_n73_n47# a_n141_n221# sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.52 as=0.136 ps=1.52 w=0.47 l=0.15
C0 a_n73_n47# a_15_n47# 0.0779f
C1 a_n33_n135# a_15_n47# 0.0213f
C2 a_n33_n135# a_n73_n47# 0.0213f
C3 a_15_n47# a_n141_n221# 0.0686f
C4 a_n73_n47# a_n141_n221# 0.0686f
C5 a_n33_n135# a_n141_n221# 0.317f
.ends

.subckt th08 Vin V08 m1_477_n803# Vp Vn
XXM0 Vn Vn m1_477_n803# Vin sky130_fd_pr__nfet_01v8_JSJ4VK
XXM1 Vp Vin m1_477_n803# Vp Vn sky130_fd_pr__pfet_01v8_EVXEQ2
XXM2 Vp Vp V08 m1_477_n803# Vn sky130_fd_pr__pfet_01v8_BBE9QE
XXM3 Vn Vn m1_477_n803# V08 sky130_fd_pr__nfet_01v8_NCP4B2
C0 V08 Vin 0.00163f
C1 Vp Vin 0.0933f
C2 V08 m1_477_n803# 0.108f
C3 Vp m1_477_n803# 0.154f
C4 V08 Vp 0.0461f
C5 Vin m1_477_n803# 0.356f
C6 m1_477_n803# Vn 0.656f
C7 Vin Vn 1.02f
C8 V08 Vn 0.271f
C9 Vp Vn 1.66f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFRTVB a_n410_n216# a_n250_n130# a_n308_n42# a_250_n42#
X0 a_250_n42# a_n250_n130# a_n308_n42# a_n410_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.5
C0 a_250_n42# a_n250_n130# 0.0209f
C1 a_250_n42# a_n308_n42# 0.011f
C2 a_n308_n42# a_n250_n130# 0.0209f
C3 a_250_n42# a_n410_n216# 0.0852f
C4 a_n308_n42# a_n410_n216# 0.0853f
C5 a_n250_n130# a_n410_n216# 1.48f
.ends

.subckt sky130_fd_pr__pfet_01v8_XQZLDL a_15_n240# w_n211_n459# a_n73_n240# a_n33_n337#
+ VSUBS
X0 a_15_n240# a_n33_n337# a_n73_n240# w_n211_n459# sky130_fd_pr__pfet_01v8 ad=0.696 pd=5.38 as=0.696 ps=5.38 w=2.4 l=0.15
C0 a_n73_n240# a_15_n240# 0.385f
C1 a_n73_n240# w_n211_n459# 0.0371f
C2 a_n73_n240# a_n33_n337# 0.0313f
C3 a_n33_n337# a_15_n240# 0.0313f
C4 a_15_n240# w_n211_n459# 0.163f
C5 a_n33_n337# w_n211_n459# 0.206f
C6 a_15_n240# VSUBS 0.11f
C7 a_n73_n240# VSUBS 0.195f
C8 a_n33_n337# VSUBS 0.139f
C9 w_n211_n459# VSUBS 1.47f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GC6 a_200_n42# w_n396_n261# a_n200_n139# a_n258_n42#
+ VSUBS
X0 a_200_n42# a_n200_n139# a_n258_n42# w_n396_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_n258_n42# a_200_n42# 0.0134f
C1 a_n258_n42# w_n396_n261# 0.0269f
C2 a_n258_n42# a_n200_n139# 0.0196f
C3 a_n200_n139# a_200_n42# 0.0196f
C4 a_200_n42# w_n396_n261# 0.0498f
C5 a_n200_n139# w_n396_n261# 0.73f
C6 a_200_n42# VSUBS 0.0338f
C7 a_n258_n42# VSUBS 0.0488f
C8 a_n200_n139# VSUBS 0.563f
C9 w_n396_n261# VSUBS 1.69f
.ends

.subckt sky130_fd_pr__nfet_01v8_ATLS57 a_15_n200# a_n73_n200# a_n33_n288# a_n141_n374#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n141_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_15_n200# a_n33_n288# 0.0312f
C1 a_15_n200# a_n73_n200# 0.321f
C2 a_n73_n200# a_n33_n288# 0.0312f
C3 a_15_n200# a_n141_n374# 0.233f
C4 a_n73_n200# a_n141_n374# 0.199f
C5 a_n33_n288# a_n141_n374# 0.341f
.ends

.subckt th13 V13 Vin m1_831_275# Vn Vp m1_559_n458#
XXM0 Vn m1_559_n458# Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vn Vin m1_559_n458# m1_831_275# sky130_fd_pr__nfet_01v8_ZFRTVB
XXM2 Vp Vp m1_831_275# Vin Vn sky130_fd_pr__pfet_01v8_XQZLDL
XXM3 V13 Vp m1_831_275# Vp Vn sky130_fd_pr__pfet_01v8_VZ9GC6
XXM4 V13 Vn m1_831_275# Vn sky130_fd_pr__nfet_01v8_ATLS57
C0 m1_831_275# V13 0.184f
C1 Vin m1_831_275# 0.197f
C2 Vin V13 0.0076f
C3 m1_559_n458# Vp 0.0628f
C4 m1_559_n458# Vn 0.152f
C5 Vp Vn 0.206f
C6 m1_559_n458# m1_831_275# 0.0183f
C7 m1_831_275# Vp 0.215f
C8 Vp V13 0.135f
C9 m1_559_n458# Vin 0.181f
C10 Vin Vp 0.176f
C11 m1_831_275# Vn 0.232f
C12 V13 Vn 0.0706f
C13 Vin Vn 0.347f
C14 m1_831_275# 0 1.05f
C15 Vin 0 1.79f
C16 V13 0 0.365f
C17 Vn 0 0.117f
C18 Vp 0 3.98f
C19 m1_559_n458# 0 0.286f
.ends

.subckt sky130_fd_pr__nfet_01v8_DD6SHA a_n33_n130# a_15_n42# a_n175_n182# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n33_n130# a_15_n42# 0.0209f
C1 a_15_n42# a_n73_n42# 0.0699f
C2 a_n33_n130# a_n73_n42# 0.0209f
C3 a_15_n42# a_n175_n182# 0.0637f
C4 a_n73_n42# a_n175_n182# 0.0716f
C5 a_n33_n130# a_n175_n182# 0.314f
.ends

.subckt sky130_fd_pr__pfet_01v8_7DPLFP w_n245_n261# a_n107_n42# a_n49_n139# a_49_n42#
+ VSUBS
X0 a_49_n42# a_n49_n139# a_n107_n42# w_n245_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.49
C0 a_49_n42# a_n107_n42# 0.0396f
C1 w_n245_n261# a_49_n42# 0.0224f
C2 a_49_n42# a_n49_n139# 0.00895f
C3 w_n245_n261# a_n107_n42# 0.0224f
C4 a_n107_n42# a_n49_n139# 0.00895f
C5 w_n245_n261# a_n49_n139# 0.221f
C6 a_49_n42# VSUBS 0.0487f
C7 a_n107_n42# VSUBS 0.0487f
C8 a_n49_n139# VSUBS 0.206f
C9 w_n245_n261# VSUBS 0.876f
.ends

.subckt sky130_fd_pr__pfet_01v8_MDPZBH a_n102_n42# a_44_n42# a_n44_n139# w_n240_n261#
+ VSUBS
X0 a_44_n42# a_n44_n139# a_n102_n42# w_n240_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.44
C0 a_44_n42# a_n102_n42# 0.0423f
C1 w_n240_n261# a_44_n42# 0.0224f
C2 a_44_n42# a_n44_n139# 0.00823f
C3 w_n240_n261# a_n102_n42# 0.0224f
C4 a_n102_n42# a_n44_n139# 0.00823f
C5 w_n240_n261# a_n44_n139# 0.208f
C6 a_44_n42# VSUBS 0.0485f
C7 a_n102_n42# VSUBS 0.0485f
C8 a_n44_n139# VSUBS 0.191f
C9 w_n240_n261# VSUBS 0.858f
.ends

.subckt th06 Vp Vin V06 Vn m1_904_n796#
XXM0 Vin m1_904_n796# Vn Vn sky130_fd_pr__nfet_01v8_DD6SHA
XXM1 Vp Vp Vin m1_904_n796# Vn sky130_fd_pr__pfet_01v8_7DPLFP
XXM2 Vp V06 m1_904_n796# Vp Vn sky130_fd_pr__pfet_01v8_MDPZBH
XXM3 Vn m1_904_n796# V06 Vn sky130_fd_pr__nfet_01v8_MYA4RC
C0 Vn Vp 0.0214f
C1 V06 Vp 0.06f
C2 Vin Vn 0.0188f
C3 m1_904_n796# Vn 0.0382f
C4 m1_904_n796# V06 0.157f
C5 Vin Vp 0.113f
C6 m1_904_n796# Vp 0.197f
C7 V06 Vn 0.00141f
C8 m1_904_n796# Vin 0.203f
C9 Vp 0 1.69f
C10 V06 0 0.217f
C11 Vn 0 0.286f
C12 m1_904_n796# 0 0.495f
C13 Vin 0 0.524f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGAKDL a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
+ VSUBS
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n73_n200# a_15_n200# 0.321f
C1 a_n33_n297# a_15_n200# 0.0293f
C2 a_15_n200# w_n211_n419# 0.0336f
C3 a_n73_n200# a_n33_n297# 0.0293f
C4 a_n73_n200# w_n211_n419# 0.0336f
C5 a_n33_n297# w_n211_n419# 0.191f
C6 a_15_n200# VSUBS 0.164f
C7 a_n73_n200# VSUBS 0.164f
C8 a_n33_n297# VSUBS 0.147f
C9 w_n211_n419# VSUBS 1.14f
.ends

.subckt sky130_fd_pr__nfet_01v8_4X3CDA a_n306_n216# a_n180_n130# a_n238_n42# a_180_n42#
X0 a_180_n42# a_n180_n130# a_n238_n42# a_n306_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.8
C0 a_180_n42# a_n238_n42# 0.0147f
C1 a_180_n42# a_n180_n130# 0.0189f
C2 a_n238_n42# a_n180_n130# 0.0189f
C3 a_180_n42# a_n306_n216# 0.075f
C4 a_n238_n42# a_n306_n216# 0.075f
C5 a_n180_n130# a_n306_n216# 1.1f
.ends

.subckt sky130_fd_pr__pfet_01v8_MWB9BZ a_15_n43# w_n211_n262# a_n73_n43# a_n33_n140#
+ VSUBS
X0 a_15_n43# a_n33_n140# a_n73_n43# w_n211_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.15
C0 a_n73_n43# a_15_n43# 0.0715f
C1 a_n33_n140# a_15_n43# 0.0193f
C2 a_15_n43# w_n211_n262# 0.0198f
C3 a_n73_n43# a_n33_n140# 0.0193f
C4 a_n73_n43# w_n211_n262# 0.0198f
C5 a_n33_n140# w_n211_n262# 0.187f
C6 a_15_n43# VSUBS 0.0453f
C7 a_n73_n43# VSUBS 0.0453f
C8 a_n33_n140# VSUBS 0.143f
C9 w_n211_n262# VSUBS 0.752f
.ends

.subckt sky130_fd_pr__nfet_01v8_L9ESAD a_n175_n190# a_n73_n50# a_n33_n138# a_15_n50#
X0 a_15_n50# a_n33_n138# a_n73_n50# a_n175_n190# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_15_n50# a_n73_n50# 0.0826f
C1 a_15_n50# a_n33_n138# 0.0216f
C2 a_n73_n50# a_n33_n138# 0.0216f
C3 a_15_n50# a_n175_n190# 0.0704f
C4 a_n73_n50# a_n175_n190# 0.0797f
C5 a_n33_n138# a_n175_n190# 0.315f
.ends

.subckt th11 Vp V11 Vin Vn m1_577_n654# m1_705_187#
XXM0 Vn Vp Vn m1_577_n654# Vn sky130_fd_pr__pfet_01v8_XGAKDL
XXM1 Vn Vin m1_577_n654# m1_705_187# sky130_fd_pr__nfet_01v8_4X3CDA
XXM2 m1_705_187# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_MWB9BZ
XXM3 V11 Vp m1_705_187# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM4 Vn Vn m1_705_187# V11 sky130_fd_pr__nfet_01v8_L9ESAD
C0 m1_705_187# V11 0.376f
C1 m1_705_187# Vin 0.0649f
C2 m1_705_187# Vn 0.463f
C3 m1_705_187# Vp 0.286f
C4 V11 Vin 2.69e-19
C5 m1_705_187# m1_577_n654# 0.0258f
C6 Vn V11 0.00327f
C7 Vn Vin 0.135f
C8 Vp V11 0.026f
C9 Vp Vin 0.285f
C10 m1_577_n654# V11 6.11e-19
C11 m1_577_n654# Vin 0.213f
C12 Vp Vn 0.0775f
C13 Vn m1_577_n654# 0.0457f
C14 Vp m1_577_n654# 0.0405f
C15 Vp 0 2.61f
C16 m1_705_187# 0 0.602f
C17 V11 0 0.404f
C18 Vn 0 0.355f
C19 Vin 0 1.27f
C20 m1_577_n654# 0 0.286f
.ends

.subckt sky130_fd_pr__nfet_01v8_42G4RD a_n80_n42# a_n148_n216# a_n33_n130# a_22_n42#
X0 a_22_n42# a_n33_n130# a_n80_n42# a_n148_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_22_n42# a_n80_n42# 0.0604f
C1 a_n33_n130# a_n80_n42# 0.00866f
C2 a_22_n42# a_n33_n130# 0.00866f
C3 a_22_n42# a_n148_n216# 0.0698f
C4 a_n80_n42# a_n148_n216# 0.0698f
C5 a_n33_n130# a_n148_n216# 0.321f
.ends

.subckt sky130_fd_pr__pfet_01v8_DDPLQ8 a_n77_n42# w_n215_n261# a_n33_n139# a_19_n42#
+ VSUBS
X0 a_19_n42# a_n33_n139# a_n77_n42# w_n215_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_19_n42# a_n33_n139# 0.0127f
C1 a_n77_n42# a_19_n42# 0.0641f
C2 w_n215_n261# a_19_n42# 0.0399f
C3 a_n77_n42# a_n33_n139# 0.0127f
C4 w_n215_n261# a_n33_n139# 0.181f
C5 a_n77_n42# w_n215_n261# 0.017f
C6 a_19_n42# VSUBS 0.035f
C7 a_n77_n42# VSUBS 0.05f
C8 a_n33_n139# VSUBS 0.149f
C9 w_n215_n261# VSUBS 0.797f
.ends

.subckt sky130_fd_pr__nfet_01v8_VWP3K3 a_n33_n130# a_15_n42# a_n141_182# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n141_182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_15_n42# a_n73_n42# 0.0699f
C1 a_n33_n130# a_n73_n42# 0.0209f
C2 a_15_n42# a_n33_n130# 0.0209f
C3 a_15_n42# a_n141_182# 0.0643f
C4 a_n73_n42# a_n141_182# 0.0643f
C5 a_n33_n130# a_n141_182# 0.317f
.ends

.subckt sky130_fd_pr__pfet_01v8_LZD9A4 a_n80_n42# a_22_n42# a_n33_n139# w_n218_n261#
+ VSUBS
X0 a_22_n42# a_n33_n139# a_n80_n42# w_n218_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_22_n42# a_n33_n139# 0.0084f
C1 a_n80_n42# a_22_n42# 0.0604f
C2 w_n218_n261# a_22_n42# 0.0222f
C3 a_n80_n42# a_n33_n139# 0.0084f
C4 w_n218_n261# a_n33_n139# 0.185f
C5 a_n80_n42# w_n218_n261# 0.0222f
C6 a_22_n42# VSUBS 0.0474f
C7 a_n80_n42# VSUBS 0.0474f
C8 a_n33_n139# VSUBS 0.149f
C9 w_n218_n261# VSUBS 0.775f
.ends

.subckt sky130_fd_pr__nfet_01v8_VRD6K3 a_n77_n42# a_n145_n214# a_n33_n130# a_19_n42#
X0 a_19_n42# a_n33_n130# a_n77_n42# a_n145_n214# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_19_n42# a_n77_n42# 0.0641f
C1 a_n33_n130# a_n77_n42# 0.0136f
C2 a_19_n42# a_n33_n130# 0.0136f
C3 a_19_n42# a_n145_n214# 0.0677f
C4 a_n77_n42# a_n145_n214# 0.0677f
C5 a_n33_n130# a_n145_n214# 0.32f
.ends

.subckt th04 Vp V04 Vin Vn m1_892_n998# m1_620_n488#
XXM0 m1_892_n998# Vn Vin Vn sky130_fd_pr__nfet_01v8_42G4RD
XXM1 m1_620_n488# Vp Vin m1_892_n998# Vn sky130_fd_pr__pfet_01v8_DDPLQ8
XXM2 Vp m1_620_n488# Vn Vp sky130_fd_pr__nfet_01v8_VWP3K3
XXM3 Vp V04 m1_892_n998# Vp Vn sky130_fd_pr__pfet_01v8_LZD9A4
XXM4 Vn Vn m1_892_n998# V04 sky130_fd_pr__nfet_01v8_VRD6K3
C0 Vin V04 0.00141f
C1 Vp V04 0.0462f
C2 m1_892_n998# V04 0.13f
C3 Vp Vin 0.14f
C4 Vn V04 0.0639f
C5 m1_892_n998# Vin 0.463f
C6 V04 m1_620_n488# 0.00264f
C7 Vp m1_892_n998# 0.383f
C8 Vin Vn 0.0468f
C9 Vin m1_620_n488# 0.0346f
C10 Vp Vn 0.0386f
C11 Vp m1_620_n488# 0.17f
C12 m1_892_n998# Vn 0.1f
C13 m1_892_n998# m1_620_n488# 0.0117f
C14 Vn m1_620_n488# 2.16e-19
C15 Vin 0 0.679f
C16 V04 0 0.287f
C17 Vn 0 0.259f
C18 m1_892_n998# 0 0.832f
C19 Vp 0 2.13f
C20 m1_620_n488# 0 0.0632f
.ends

.subckt Analog Vin Vp V01 V02 V03 V04 V08 V07 V06 V09 V10 V11 V12 V13 V14 V15 V05
+ Vn
Xth02_0 th15_0/Vin V02 Vp th02_0/m1_983_133# th02_0/m1_571_144# Vn th02
Xth09_0 V09 Vin Vn th09_0/m1_485_n505# Vp th09_0/m1_962_372# th09
Xth14_0 V14 th15_0/Vin Vn th14_0/m1_641_n318# Vp th14_0/m1_891_419# th14
Xth07_0 Vin V07 Vp th07_0/m1_808_n892# Vn th07
Xth12_0 Vp V12 Vin th12_0/m1_529_n42# th12_0/m1_394_n856# Vn th12
Xth05_0 Vp V05 Vin th05_0/m1_752_n794# Vn th05
Xth10_0 Vp V10 Vin Vn th10_0/m1_502_n495# th10_0/m1_536_174# th10
Xth03_0 V03 Vin Vp th03_0/m1_890_n844# th03_0/m1_638_n591# Vn th03
Xth01_0 Vp th15_0/Vin V01 th01_0/m1_991_n1219# Vn th01_0/m1_571_n501# th01
Xpreamp_0 Vp Vin th15_0/Vin Vn preamp
Xth15_0 V15 th15_0/Vin th15_0/m1_597_n912# Vp th15_0/m1_849_n157# Vn th15
Xth08_0 Vin V08 th08_0/m1_477_n803# Vp Vn th08
Xth13_0 V13 Vin th13_0/m1_831_275# Vn Vp th13_0/m1_559_n458# th13
Xth06_0 Vp Vin V06 Vn th06_0/m1_904_n796# th06
Xth11_0 Vp V11 Vin Vn th11_0/m1_577_n654# th11_0/m1_705_187# th11
Xth04_0 Vp V04 Vin Vn th04_0/m1_892_n998# th04_0/m1_620_n488# th04
C0 th11_0/m1_705_187# th01_0/m1_571_n501# 9.49e-20
C1 V01 th15_0/Vin 3.18e-19
C2 th13_0/m1_831_275# V13 0.0112f
C3 th08_0/m1_477_n803# th04_0/m1_620_n488# 6.18e-20
C4 Vn V04 0.00815f
C5 Vp V14 0.0751f
C6 th14_0/m1_891_419# V11 0.0143f
C7 V09 th14_0/m1_641_n318# 6.83e-21
C8 Vn th02_0/m1_571_144# 0.0142f
C9 Vn th07_0/m1_808_n892# 0.00532f
C10 Vn th15_0/Vin 1.48f
C11 V15 th15_0/Vin 1.81e-19
C12 th09_0/m1_485_n505# th02_0/m1_983_133# 0.00736f
C13 th01_0/m1_991_n1219# V01 0.00159f
C14 th12_0/m1_394_n856# V12 2.12e-19
C15 th15_0/m1_849_n157# th13_0/m1_831_275# 0.0859f
C16 th11_0/m1_705_187# Vin 0.278f
C17 th12_0/m1_394_n856# th12_0/m1_529_n42# 1.78e-33
C18 Vin th13_0/m1_831_275# 0.0149f
C19 th14_0/m1_891_419# Vn 0.0525f
C20 V08 Vin 0.164f
C21 th11_0/m1_577_n654# V02 3.56e-21
C22 Vn th01_0/m1_991_n1219# 0.00203f
C23 th12_0/m1_394_n856# th14_0/m1_641_n318# 0.00861f
C24 V14 th15_0/Vin 6.88e-20
C25 Vn th10_0/m1_536_174# 0.0537f
C26 V11 th11_0/m1_577_n654# 1.77e-19
C27 V09 th09_0/m1_485_n505# 0.0182f
C28 V06 Vin 0.094f
C29 V07 Vin 0.0909f
C30 th11_0/m1_705_187# Vp 0.0213f
C31 th08_0/m1_477_n803# Vin 0.055f
C32 Vp th13_0/m1_831_275# 0.0414f
C33 th03_0/m1_890_n844# th01_0/m1_571_n501# 0.00797f
C34 V08 Vp 0.0346f
C35 th14_0/m1_891_419# V14 0.0202f
C36 V10 th12_0/m1_529_n42# 2.39e-20
C37 Vn th11_0/m1_577_n654# 0.0365f
C38 V06 Vp 0.025f
C39 V07 Vp 0.0372f
C40 Vp th08_0/m1_477_n803# 0.0268f
C41 V12 Vin 1.77e-19
C42 V03 Vin 4.84e-19
C43 Vn th03_0/m1_638_n591# 0.0534f
C44 th11_0/m1_705_187# th02_0/m1_571_144# 1.03e-19
C45 Vn th10_0/m1_502_n495# 0.00962f
C46 Vn th05_0/m1_752_n794# 0.00258f
C47 th11_0/m1_705_187# th15_0/Vin 0.0359f
C48 V08 V04 2.69e-20
C49 Vin th12_0/m1_529_n42# 0.0104f
C50 th03_0/m1_890_n844# Vin 4.79e-20
C51 th13_0/m1_831_275# th15_0/Vin 0.0168f
C52 Vn V02 0.00543f
C53 V08 th07_0/m1_808_n892# 0.0102f
C54 th13_0/m1_559_n458# th12_0/m1_529_n42# 9.14e-21
C55 Vin th14_0/m1_641_n318# 0.0621f
C56 Vn V11 0.0184f
C57 th08_0/m1_477_n803# V04 4.48e-19
C58 Vp V12 0.0535f
C59 V03 Vp 0.011f
C60 th11_0/m1_705_187# th14_0/m1_891_419# 0.00195f
C61 V06 th07_0/m1_808_n892# 5.69e-20
C62 V07 th07_0/m1_808_n892# 0.00298f
C63 th11_0/m1_705_187# th01_0/m1_991_n1219# 0.00184f
C64 Vn V01 0.00263f
C65 th07_0/m1_808_n892# th08_0/m1_477_n803# 4.41e-19
C66 Vp th12_0/m1_529_n42# 0.0641f
C67 Vp th03_0/m1_890_n844# 0.0291f
C68 Vp th14_0/m1_641_n318# 0.0569f
C69 th06_0/m1_904_n796# V05 1.38e-20
C70 Vn V15 2.4e-20
C71 th09_0/m1_485_n505# Vin 0.0287f
C72 th02_0/m1_983_133# Vin 0.0835f
C73 V12 th15_0/Vin 1.05e-21
C74 V03 th15_0/Vin 1.39e-20
C75 th09_0/m1_485_n505# th13_0/m1_559_n458# 0.00612f
C76 th12_0/m1_529_n42# th15_0/Vin 0.0262f
C77 th03_0/m1_890_n844# th15_0/Vin 0.00307f
C78 Vn V14 0.0201f
C79 th14_0/m1_641_n318# th15_0/Vin 0.0354f
C80 Vp th09_0/m1_485_n505# 0.0355f
C81 th14_0/m1_891_419# V12 2.97e-19
C82 Vp th02_0/m1_983_133# 0.0442f
C83 V09 Vin 0.00465f
C84 Vin th06_0/m1_904_n796# 0.0348f
C85 V09 th13_0/m1_559_n458# 0.00378f
C86 th14_0/m1_891_419# th12_0/m1_529_n42# 0.0381f
C87 V12 th10_0/m1_536_174# 9.23e-19
C88 th11_0/m1_705_187# V11 5.77e-19
C89 V06 th05_0/m1_752_n794# 0.001f
C90 V09 th09_0/m1_962_372# 8.77e-19
C91 th10_0/m1_536_174# th12_0/m1_529_n42# 0.002f
C92 V07 th05_0/m1_752_n794# 4.77e-21
C93 Vin th04_0/m1_892_n998# 0.111f
C94 V09 Vp 0.00542f
C95 th09_0/m1_485_n505# th02_0/m1_571_144# 0.00503f
C96 Vp th06_0/m1_904_n796# 0.0232f
C97 th12_0/m1_394_n856# Vin 0.0013f
C98 th09_0/m1_485_n505# th15_0/Vin 0.113f
C99 th02_0/m1_983_133# th15_0/Vin 0.0246f
C100 th12_0/m1_394_n856# th13_0/m1_559_n458# 3.47e-20
C101 th11_0/m1_705_187# Vn -0.0527f
C102 th04_0/m1_620_n488# Vin 0.00123f
C103 Vp th04_0/m1_892_n998# 0.0374f
C104 th15_0/m1_849_n157# V13 0.0171f
C105 Vn th13_0/m1_831_275# 0.0355f
C106 V08 Vn 7.17e-19
C107 th08_0/m1_477_n803# V01 4.9e-21
C108 Vin V05 0.00116f
C109 th14_0/m1_891_419# th09_0/m1_485_n505# 3.27e-19
C110 Vin V13 0.00669f
C111 Vp th12_0/m1_394_n856# 0.0145f
C112 th12_0/m1_529_n42# th10_0/m1_502_n495# 8.5e-20
C113 V09 th02_0/m1_571_144# 3.21e-19
C114 th01_0/m1_571_n501# Vin 6.06e-19
C115 Vn V06 5.44e-19
C116 V09 th15_0/Vin 0.0644f
C117 Vn V07 0.00179f
C118 Vp th04_0/m1_620_n488# 0.00246f
C119 Vn th08_0/m1_477_n803# 0.00115f
C120 th07_0/m1_808_n892# th06_0/m1_904_n796# 2e-19
C121 th03_0/m1_890_n844# V02 0.00134f
C122 V04 th04_0/m1_892_n998# 1.47e-19
C123 V10 Vin 0.00422f
C124 th15_0/m1_597_n912# Vin 3.87e-19
C125 Vp V05 0.00375f
C126 th07_0/m1_808_n892# th04_0/m1_892_n998# 1.1e-19
C127 th04_0/m1_892_n998# th15_0/Vin 0.00125f
C128 Vp V13 0.00713f
C129 th15_0/m1_849_n157# Vin 0.00238f
C130 th14_0/m1_891_419# V09 3.7e-19
C131 Vp th01_0/m1_571_n501# 0.0265f
C132 th12_0/m1_394_n856# th15_0/Vin 0.0129f
C133 Vn V12 0.0372f
C134 V03 Vn 2.75e-19
C135 th02_0/m1_983_133# th11_0/m1_577_n654# 1.64e-19
C136 Vin th13_0/m1_559_n458# 0.0257f
C137 V10 Vp 0.0332f
C138 th04_0/m1_620_n488# th15_0/Vin 2.61e-19
C139 Vp th15_0/m1_597_n912# -2.84e-32
C140 Vn th12_0/m1_529_n42# 0.0621f
C141 Vn th03_0/m1_890_n844# 0.0101f
C142 th01_0/m1_991_n1219# th04_0/m1_892_n998# 0.0226f
C143 th03_0/m1_638_n591# th02_0/m1_983_133# 0.0193f
C144 Vp th15_0/m1_849_n157# 0.0962f
C145 th09_0/m1_962_372# Vin 6.36e-19
C146 Vn th14_0/m1_641_n318# 0.0401f
C147 th14_0/m1_891_419# th12_0/m1_394_n856# 5.71e-20
C148 V13 th15_0/Vin 1e-23
C149 th02_0/m1_983_133# V02 0.0161f
C150 Vp Vin 1.96f
C151 th01_0/m1_571_n501# th15_0/Vin -5.68e-32
C152 Vp th13_0/m1_559_n458# 0.0105f
C153 th01_0/m1_991_n1219# th04_0/m1_620_n488# 7.52e-20
C154 th12_0/m1_529_n42# V14 1.86e-19
C155 Vp th09_0/m1_962_372# 0.0369f
C156 th15_0/m1_597_n912# th15_0/Vin 0.0049f
C157 th05_0/m1_752_n794# th06_0/m1_904_n796# 0.00251f
C158 th15_0/m1_849_n157# th15_0/Vin 6.18e-19
C159 V04 Vin 0.175f
C160 V08 V07 6.64e-21
C161 V08 th08_0/m1_477_n803# 0.00927f
C162 th02_0/m1_571_144# Vin 0.00869f
C163 Vn th09_0/m1_485_n505# 0.0537f
C164 th07_0/m1_808_n892# Vin 0.0324f
C165 Vn th02_0/m1_983_133# 0.157f
C166 Vin th15_0/Vin 0.87f
C167 th13_0/m1_559_n458# th15_0/Vin 0.11f
C168 V07 V06 5.71e-22
C169 V07 th08_0/m1_477_n803# 9.47e-21
C170 th09_0/m1_962_372# th02_0/m1_571_144# 0.0112f
C171 V10 th10_0/m1_536_174# 0.0035f
C172 th09_0/m1_962_372# th15_0/Vin 0.0637f
C173 Vp V04 0.00153f
C174 th14_0/m1_891_419# Vin 0.0347f
C175 Vp th02_0/m1_571_144# 0.026f
C176 Vp th07_0/m1_808_n892# 0.0183f
C177 Vp th15_0/Vin 1.24f
C178 th01_0/m1_991_n1219# Vin 0.0315f
C179 V01 th04_0/m1_892_n998# 0.0123f
C180 V09 Vn 0.0232f
C181 th05_0/m1_752_n794# V05 1.39e-19
C182 Vn th06_0/m1_904_n796# 0.00332f
C183 th13_0/m1_831_275# th12_0/m1_529_n42# 1.36e-20
C184 th10_0/m1_536_174# Vin 0.0133f
C185 th11_0/m1_705_187# th14_0/m1_641_n318# 5.69e-22
C186 Vn th04_0/m1_892_n998# 4.09e-20
C187 th14_0/m1_891_419# Vp 0.0102f
C188 V01 th04_0/m1_620_n488# 0.00118f
C189 th07_0/m1_808_n892# V04 6.58e-21
C190 th01_0/m1_991_n1219# Vp 0.0315f
C191 Vn th12_0/m1_394_n856# 0.0035f
C192 Vp th10_0/m1_536_174# 0.0514f
C193 th02_0/m1_571_144# th15_0/Vin 0.00185f
C194 Vin th11_0/m1_577_n654# 0.0113f
C195 Vin th10_0/m1_502_n495# 1.09e-19
C196 th05_0/m1_752_n794# Vin 0.00963f
C197 Vn V05 6.36e-19
C198 th01_0/m1_991_n1219# V04 2.28e-19
C199 th09_0/m1_485_n505# th13_0/m1_831_275# 2.23e-19
C200 Vn V13 0.0182f
C201 V12 th12_0/m1_529_n42# 3.26e-19
C202 V03 th03_0/m1_890_n844# 7.56e-19
C203 Vin V02 0.292f
C204 th14_0/m1_891_419# th15_0/Vin 0.00394f
C205 Vn th01_0/m1_571_n501# 0.00241f
C206 Vp th11_0/m1_577_n654# 0.0262f
C207 th01_0/m1_991_n1219# th15_0/Vin 0.00291f
C208 V15 V13 0.00246f
C209 V11 Vin 0.0579f
C210 th10_0/m1_536_174# th15_0/Vin 3.79e-20
C211 Vp th03_0/m1_638_n591# 0.0167f
C212 Vp th10_0/m1_502_n495# 0.035f
C213 Vp th05_0/m1_752_n794# 8.03e-19
C214 V10 Vn 0.0168f
C215 V01 Vin 0.00532f
C216 Vn th15_0/m1_597_n912# 0.106f
C217 Vp V02 0.00255f
C218 th14_0/m1_891_419# th01_0/m1_991_n1219# 0.0018f
C219 Vn th15_0/m1_849_n157# 0.0342f
C220 V15 th15_0/m1_849_n157# 0.0154f
C221 V08 th06_0/m1_904_n796# 9.74e-22
C222 Vp V11 0.0406f
C223 Vn Vin 1.97f
C224 th02_0/m1_571_144# th11_0/m1_577_n654# 0.0183f
C225 th11_0/m1_577_n654# th15_0/Vin 0.016f
C226 Vn th13_0/m1_559_n458# 0.017f
C227 Vp V01 0.116f
C228 V08 th04_0/m1_892_n998# 3.48e-19
C229 V06 th06_0/m1_904_n796# -1.42e-32
C230 V03 th02_0/m1_983_133# 2.47e-20
C231 V07 th06_0/m1_904_n796# 0.00384f
C232 th03_0/m1_638_n591# th15_0/Vin 0.0177f
C233 th11_0/m1_705_187# th12_0/m1_394_n856# 6.45e-22
C234 th05_0/m1_752_n794# th07_0/m1_808_n892# 1.42e-20
C235 th08_0/m1_477_n803# th06_0/m1_904_n796# 2.84e-21
C236 Vn th09_0/m1_962_372# 0.00557f
C237 th12_0/m1_394_n856# th13_0/m1_831_275# 4.06e-20
C238 th02_0/m1_983_133# th03_0/m1_890_n844# 0.00411f
C239 th15_0/Vin V02 0.00312f
C240 Vn Vp 1.69f
C241 th08_0/m1_477_n803# th04_0/m1_892_n998# 0.00506f
C242 th09_0/m1_485_n505# th14_0/m1_641_n318# 6.8e-20
C243 Vin V14 0.00129f
C244 V08 th04_0/m1_620_n488# 3.51e-21
C245 V11 th02_0/m1_571_144# 4.75e-20
C246 Vp V15 0.00307f
C247 V11 th15_0/Vin 0.00172f
C248 V04 V01 1.84e-20
C249 V04 0 0.191f
C250 th04_0/m1_892_n998# 0 0.832f
C251 th04_0/m1_620_n488# 0 0.0632f
C252 th11_0/m1_705_187# 0 0.602f
C253 V11 0 0.349f
C254 Vin 0 15f
C255 th11_0/m1_577_n654# 0 0.286f
C256 V06 0 0.132f
C257 th06_0/m1_904_n796# 0 0.495f
C258 th13_0/m1_831_275# 0 1.05f
C259 V13 0 0.371f
C260 th13_0/m1_559_n458# 0 0.286f
C261 th08_0/m1_477_n803# 0 0.577f
C262 V08 0 0.139f
C263 V15 0 0.356f
C264 th15_0/m1_849_n157# 0 1.28f
C265 th15_0/m1_597_n912# 0 0.19f
C266 Vn 0 6.57f
C267 th01_0/m1_991_n1219# 0 1.24f
C268 V01 0 0.241f
C269 th01_0/m1_571_n501# 0 0.194f
C270 th15_0/Vin 0 5.76f
C271 Vp 0 43.6f
C272 V03 0 0.303f
C273 th03_0/m1_890_n844# 0 1.05f
C274 th03_0/m1_638_n591# 0 0.224f
C275 th10_0/m1_536_174# 0 0.825f
C276 V10 0 0.269f
C277 th10_0/m1_502_n495# 0 0.146f
C278 th05_0/m1_752_n794# 0 0.788f
C279 V05 0 0.321f
C280 th12_0/m1_529_n42# 0 0.861f
C281 V12 0 0.468f
C282 th12_0/m1_394_n856# 0 0.215f
C283 th07_0/m1_808_n892# 0 0.511f
C284 V07 0 0.159f
C285 th14_0/m1_891_419# 0 1.48f
C286 V14 0 0.233f
C287 th14_0/m1_641_n318# 0 0.241f
C288 th09_0/m1_485_n505# 0 1.18f
C289 V09 0 0.213f
C290 th09_0/m1_962_372# 0 0.118f
C291 V02 0 0.211f
C292 th02_0/m1_983_133# 0 1.44f
C293 th02_0/m1_571_144# 0 0.252f
.ends

