magic
tech sky130A
magscale 1 2
timestamp 1702923036
<< error_s >>
rect 996 717 1037 749
rect 1494 669 1535 701
rect 1808 621 1849 653
rect 2306 573 2347 605
rect 2620 525 2657 557
rect 2934 477 2975 509
rect 3248 429 3289 461
rect 3746 381 3787 413
rect 4558 285 4599 317
rect 4964 237 5005 269
rect 5278 189 5315 221
rect 5684 141 5713 173
rect 6274 93 6315 125
rect 6588 45 6625 77
rect 7086 -3 7127 29
rect 8082 -99 8123 -67
rect 9668 -243 9697 -211
rect 10166 -291 10207 -259
rect 11254 -387 11295 -355
rect 11844 -435 11885 -403
rect 13798 -579 13837 -547
rect 14702 -675 14743 -643
rect 15108 -723 15137 -691
rect 15422 -771 15463 -739
rect 15920 -819 15961 -787
rect 16640 -915 16677 -883
rect 17636 -1011 17649 -979
use sky130_fd_sc_hd__clkinv_1  x0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 -240 0 1 800
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 708 0 1 1514
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 628 0 1 504
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 1034 0 1 456
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  x4
timestamp 1696625445
transform 1 0 1532 0 1 408
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  x5
timestamp 1696625445
transform 1 0 1846 0 1 360
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  x6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 2344 0 1 312
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x7
timestamp 1696625445
transform 1 0 2658 0 1 264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x8
timestamp 1696625445
transform 1 0 2972 0 1 216
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  x9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3286 0 1 168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  x10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3784 0 1 120
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  x11
timestamp 1696625445
transform 1 0 4282 0 1 72
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  x12
timestamp 1696625445
transform 1 0 4596 0 1 24
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  x13
timestamp 1696625445
transform 1 0 5002 0 1 -24
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  x14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 5316 0 1 -72
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 5722 0 1 -120
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  x16
timestamp 1696625445
transform 1 0 6312 0 1 -168
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  x17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 6626 0 1 -216
box -38 -48 498 592
use sky130_fd_sc_hd__lpflow_inputiso1p_1  x18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 7124 0 1 -264
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  x19
timestamp 1696625445
transform 1 0 7622 0 1 -312
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  x20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 8120 0 1 -360
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  x21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 8618 0 1 -408
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  x22
timestamp 1696625445
transform 1 0 9300 0 1 -456
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  x23
timestamp 1696625445
transform 1 0 9706 0 1 -504
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_0  x24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 10204 0 1 -552
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  x25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 10610 0 1 -600
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  x26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 11292 0 1 -648
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  x27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 11882 0 1 -696
box -38 -48 590 592
use sky130_fd_sc_hd__a32oi_1  x28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 12472 0 1 -744
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  x29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 13154 0 1 -792
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  x30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 13836 0 1 -840
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  x31
timestamp 1696625445
transform 1 0 14426 0 1 -888
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  x32
timestamp 1696625445
transform 1 0 14740 0 1 -936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  x33
timestamp 1696625445
transform 1 0 15146 0 1 -984
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  x34
timestamp 1696625445
transform 1 0 15460 0 1 -1032
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_0  x35
timestamp 1696625445
transform 1 0 15958 0 1 -1080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  x36
timestamp 1696625445
transform 1 0 16364 0 1 -1128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_0  x37
timestamp 1696625445
transform 1 0 16678 0 1 -1176
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  x38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 17084 0 1 -1224
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  x39
timestamp 1696625445
transform 1 0 17674 0 1 -1272
box -38 -48 314 592
use Analog  x40
timestamp 1702921602
transform 1 0 17988 0 1 5480
box 0 -6800 200 200
<< end >>
