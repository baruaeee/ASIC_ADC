magic
tech sky130A
magscale 1 2
timestamp 1704880657
<< metal1 >>
rect 1931 2029 3471 2063
rect 1931 1641 1969 2029
rect 1931 1373 1965 1641
rect 3102 1523 3137 1551
rect 3102 1488 3337 1523
rect 3102 1387 3137 1488
rect 2945 931 3713 965
use th01  x1
timestamp 1704880472
transform 1 0 2808 0 1 1382
box 450 -452 1562 754
use preamp  x2
timestamp 1704880455
transform 1 0 1562 0 1 1800
box 369 -869 1682 116
<< end >>
