magic
tech sky130A
magscale 1 2
timestamp 1705440137
<< checkpaint >>
rect -1260 -2460 1460 1460
<< pwell >>
rect 1476 -990 1536 -924
rect 1762 -958 1830 -874
rect 1762 -966 1814 -958
rect 1176 -1038 1210 -1004
<< locali >>
rect 654 -474 802 -414
rect 1678 -948 1828 -870
rect 898 -1130 970 -984
<< metal1 >>
rect 0 0 200 200
rect 1474 -185 1674 -180
rect 0 -400 200 -200
rect 736 -219 2105 -185
rect 736 -474 770 -219
rect 1474 -380 1674 -219
rect 2071 -331 2105 -219
rect 1971 -365 2205 -331
rect 1417 -441 1489 -415
rect 1417 -475 1491 -441
rect 724 -538 909 -535
rect 618 -569 909 -538
rect 0 -800 200 -600
rect 618 -738 818 -569
rect 1455 -709 1489 -475
rect 1721 -709 1755 -371
rect 2107 -453 2345 -419
rect 2464 -424 2522 -362
rect 2216 -482 2251 -453
rect 2217 -611 2251 -482
rect 2217 -645 2643 -611
rect 1091 -728 1949 -709
rect 2609 -722 2643 -645
rect 724 -939 758 -738
rect 1090 -743 1949 -728
rect 1090 -895 1125 -743
rect 1915 -789 1949 -743
rect 1857 -823 2033 -789
rect 2464 -872 2664 -722
rect 931 -929 1287 -895
rect 1090 -930 1124 -929
rect 724 -973 791 -939
rect 724 -974 758 -973
rect 0 -1200 200 -1000
rect 1063 -1017 1305 -983
rect 1476 -990 1536 -924
rect 1762 -958 1830 -874
rect 2446 -922 2664 -872
rect 2446 -948 2504 -922
rect 1762 -966 1814 -958
rect 1176 -1097 1211 -1017
rect 1177 -1133 1211 -1097
rect 1596 -1133 1796 -966
rect 1177 -1166 1796 -1133
rect 1177 -1167 1795 -1166
use sky130_fd_pr__pfet_01v8_3QB9EZ  XM2
timestamp 1704962958
transform 1 0 1110 0 1 -445
box -492 -261 492 261
use sky130_fd_pr__nfet_01v8_J2SMPG  XM3
timestamp 1704962958
transform 0 -1 1138 1 0 -957
box -211 -520 211 520
use sky130_fd_pr__nfet_01v8_G45C34  XM4
timestamp 1704962958
transform -1 0 2137 0 -1 -910
box -493 -258 493 258
use sky130_fd_pr__pfet_01v8_XA2NHL  XM5
timestamp 1704962958
transform 0 -1 2115 1 0 -393
box -211 -529 211 529
<< labels >>
flabel metal1 618 -738 818 -538 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 2464 -922 2664 -722 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 1596 -1166 1796 -966 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 1474 -380 1674 -180 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vin
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vout
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
<< end >>
