magic
tech sky130A
magscale 1 2
timestamp 1706270876
<< locali >>
rect 810 -42 870 106
rect 772 -1006 818 -860
<< metal1 >>
rect 1034 146 1134 148
rect 804 112 1143 146
rect 821 -39 855 112
rect 1034 48 1143 112
rect 1109 -87 1143 48
rect 719 -177 753 -125
rect 1109 -161 1179 -87
rect 1429 -91 1463 -85
rect 1429 -125 1557 -91
rect 1429 -161 1463 -125
rect 617 -211 753 -177
rect 474 -529 574 -482
rect 617 -529 651 -211
rect 719 -333 753 -211
rect 1086 -262 1404 -222
rect 474 -563 651 -529
rect 474 -582 574 -563
rect 616 -857 650 -563
rect 820 -576 860 -392
rect 1086 -550 1126 -262
rect 1523 -288 1557 -125
rect 1508 -333 1608 -288
rect 1470 -388 1608 -333
rect 1470 -389 1521 -388
rect 1086 -576 1434 -550
rect 820 -590 1434 -576
rect 820 -616 1126 -590
rect 820 -754 860 -616
rect 1470 -645 1504 -389
rect 752 -794 1024 -754
rect 1118 -858 1174 -794
rect 1305 -819 1373 -645
rect 866 -859 900 -858
rect 735 -893 1035 -859
rect 829 -895 905 -893
rect 865 -1009 905 -895
rect 1305 -1009 1339 -819
rect 1437 -821 1504 -645
rect 1372 -920 1438 -862
rect 1518 -1009 1618 -938
rect 865 -1038 1618 -1009
rect 865 -1043 1541 -1038
use sky130_fd_pr__nfet_01v8_Q7AWK3  XM0
timestamp 1706224144
transform 0 -1 888 1 0 -826
box -216 -410 216 410
use sky130_fd_pr__pfet_01v8_EXJYQP  XM1
timestamp 1706224144
transform 0 -1 841 1 0 -217
box -359 -261 359 261
use sky130_fd_pr__pfet_01v8_HJHF6N  XM2
timestamp 1706224144
transform 1 0 1304 0 1 -123
box -325 -269 308 269
use sky130_fd_pr__nfet_01v8_N39H2X  XM3
timestamp 1706224144
transform 1 0 1406 0 1 -732
box -214 -310 214 310
<< labels >>
flabel metal1 1518 -1038 1618 -938 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 474 -582 574 -482 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 1508 -388 1608 -288 0 FreeSans 256 0 0 0 V05
port 1 nsew
flabel metal1 1034 48 1134 148 0 FreeSans 256 0 0 0 Vp
port 0 nsew
<< end >>
