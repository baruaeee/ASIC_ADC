magic
tech sky130A
magscale 1 2
timestamp 1706454272
<< nwell >>
rect -526 -261 526 261
<< pmos >>
rect -330 -42 330 42
<< pdiff >>
rect -388 30 -330 42
rect -388 -30 -376 30
rect -342 -30 -330 30
rect -388 -42 -330 -30
rect 330 30 388 42
rect 330 -30 342 30
rect 376 -30 388 30
rect 330 -42 388 -30
<< pdiffc >>
rect -376 -30 -342 30
rect 342 -30 376 30
<< nsubdiff >>
rect 456 129 490 191
rect 456 -159 490 -129
<< nsubdiffcont >>
rect 456 -129 490 129
<< poly >>
rect -330 123 330 139
rect -330 89 -314 123
rect 314 89 330 123
rect -330 42 330 89
rect -330 -89 330 -42
rect -330 -123 -314 -89
rect 314 -123 330 -89
rect -330 -139 330 -123
<< polycont >>
rect -314 89 314 123
rect -314 -123 314 -89
<< locali >>
rect 456 129 490 191
rect -330 89 -314 123
rect 314 89 330 123
rect -376 30 -342 46
rect -376 -46 -342 -30
rect 342 30 376 46
rect 342 -46 376 -30
rect -330 -123 -314 -89
rect 314 -123 330 -89
rect 456 -159 490 -129
<< viali >>
rect -314 89 314 123
rect -376 -30 -342 30
rect 342 -30 376 30
rect -314 -123 314 -89
<< metal1 >>
rect -326 123 326 129
rect -326 89 -314 123
rect 314 89 326 123
rect -326 83 326 89
rect -382 30 -336 42
rect -382 -30 -376 30
rect -342 -30 -336 30
rect -382 -42 -336 -30
rect 336 30 382 42
rect 336 -30 342 30
rect 376 -30 382 30
rect 336 -42 382 -30
rect -326 -89 326 -83
rect -326 -123 -314 -89
rect 314 -123 326 -89
rect -326 -129 326 -123
<< properties >>
string FIXED_BBOX -473 -208 473 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 3.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
