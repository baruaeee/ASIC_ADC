* NGSPICE file created from th14.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_HPNF99 a_n33_n147# a_23_n50# a_n81_n50# w_n219_n269#
+ VSUBS
X0 a_23_n50# a_n33_n147# a_n81_n50# w_n219_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.23
C0 w_n219_n269# a_n33_n147# 0.179f
C1 a_23_n50# w_n219_n269# 0.0185f
C2 a_n81_n50# w_n219_n269# 0.0455f
C3 a_23_n50# a_n33_n147# 0.00814f
C4 a_n81_n50# a_n33_n147# 0.00814f
C5 a_23_n50# a_n81_n50# 0.07f
C6 a_23_n50# VSUBS 0.0578f
C7 a_n81_n50# VSUBS 0.04f
C8 a_n33_n147# VSUBS 0.153f
C9 w_n219_n269# VSUBS 0.835f
.ends

.subckt sky130_fd_pr__nfet_01v8_JZU22M a_n213_n42# a_155_n42# a_n155_n130# a_281_n238#
X0 a_155_n42# a_n155_n130# a_n213_n42# a_281_n238# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.55
C0 a_n155_n130# a_n213_n42# 0.0178f
C1 a_155_n42# a_n155_n130# 0.0178f
C2 a_155_n42# a_n213_n42# 0.0168f
C3 a_155_n42# a_281_n238# 0.0816f
C4 a_n213_n42# a_281_n238# 0.0737f
C5 a_n155_n130# a_281_n238# 0.928f
.ends

.subckt sky130_fd_pr__pfet_01v8_TM5S5A a_n80_n147# a_n138_n50# a_80_n50# w_n276_n269#
+ VSUBS
X0 a_80_n50# a_n80_n147# a_n138_n50# w_n276_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.8
C0 w_n276_n269# a_n80_n147# 0.297f
C1 a_80_n50# w_n276_n269# 0.0231f
C2 a_n138_n50# w_n276_n269# 0.0231f
C3 a_80_n50# a_n80_n147# 0.0141f
C4 a_n138_n50# a_n80_n147# 0.0141f
C5 a_80_n50# a_n138_n50# 0.0335f
C6 a_80_n50# VSUBS 0.0565f
C7 a_n138_n50# VSUBS 0.0565f
C8 a_n80_n147# VSUBS 0.296f
C9 w_n276_n269# VSUBS 1.01f
.ends

.subckt sky130_fd_pr__pfet_01v8_AM8GZ5 w_n526_n261# a_n330_n139# a_330_n42# a_n388_n42#
+ VSUBS
X0 a_330_n42# a_n330_n139# a_n388_n42# w_n526_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.3
C0 w_n526_n261# a_n330_n139# 0.719f
C1 a_330_n42# w_n526_n261# 0.0408f
C2 a_n388_n42# w_n526_n261# 0.0179f
C3 a_330_n42# a_n330_n139# 0.0223f
C4 a_n388_n42# a_n330_n139# 0.0223f
C5 a_330_n42# a_n388_n42# 0.00853f
C6 a_330_n42# VSUBS 0.0435f
C7 a_n388_n42# VSUBS 0.0585f
C8 a_n330_n139# VSUBS 1.13f
C9 w_n526_n261# VSUBS 1.76f
.ends

.subckt sky130_fd_pr__nfet_01v8_H7HSAV a_n103_390# a_n73_n250# a_15_n250# a_n33_n338#
X0 a_15_n250# a_n33_n338# a_n73_n250# a_n103_390# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.15
C0 a_n33_n338# a_n73_n250# 0.0337f
C1 a_15_n250# a_n33_n338# 0.0337f
C2 a_15_n250# a_n73_n250# 0.401f
C3 a_15_n250# a_n103_390# 0.24f
C4 a_n73_n250# a_n103_390# 0.24f
C5 a_n33_n338# a_n103_390# 0.327f
.ends

.subckt th14 Vp V14 Vin Vn
XXM0 Vn Vn m1_641_n318# Vp Vn sky130_fd_pr__pfet_01v8_HPNF99
XXM1 m1_641_n318# m1_891_419# Vin Vn sky130_fd_pr__nfet_01v8_JZU22M
XXM2 Vin Vp m1_891_419# Vp Vn sky130_fd_pr__pfet_01v8_TM5S5A
XXM3 Vp m1_891_419# V14 Vp Vn sky130_fd_pr__pfet_01v8_AM8GZ5
XXM4 Vn Vn V14 m1_891_419# sky130_fd_pr__nfet_01v8_H7HSAV
C0 V14 Vp 0.0858f
C1 m1_891_419# V14 0.249f
C2 m1_641_n318# Vp 0.0615f
C3 m1_891_419# m1_641_n318# 0.00289f
C4 Vp Vin 0.201f
C5 m1_891_419# Vin 0.132f
C6 V14 Vin 0.00516f
C7 m1_641_n318# Vin 0.229f
C8 m1_891_419# Vp 0.227f
C9 m1_891_419# Vn 1.69f
C10 V14 Vn 0.273f
C11 Vp Vn 3.44f
C12 Vin Vn 1.76f
C13 m1_641_n318# Vn 0.311f
.ends

