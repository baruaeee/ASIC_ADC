magic
tech sky130A
timestamp 1703732895
<< pwell >>
rect -1073 -126 1073 126
<< nmos >>
rect -975 -21 975 21
<< ndiff >>
rect -1004 15 -975 21
rect -1004 -15 -998 15
rect -981 -15 -975 15
rect -1004 -21 -975 -15
rect 975 15 1004 21
rect 975 -15 981 15
rect 998 -15 1004 15
rect 975 -21 1004 -15
<< ndiffc >>
rect -998 -15 -981 15
rect 981 -15 998 15
<< psubdiff >>
rect -1055 91 -1007 108
rect 1007 91 1055 108
rect -1055 60 -1038 91
rect 1038 60 1055 91
rect -1055 -91 -1038 -60
rect 1038 -91 1055 -60
rect -1055 -108 -1007 -91
rect 1007 -108 1055 -91
<< psubdiffcont >>
rect -1007 91 1007 108
rect -1055 -60 -1038 60
rect 1038 -60 1055 60
rect -1007 -108 1007 -91
<< poly >>
rect -975 57 975 65
rect -975 40 -967 57
rect 967 40 975 57
rect -975 21 975 40
rect -975 -40 975 -21
rect -975 -57 -967 -40
rect 967 -57 975 -40
rect -975 -65 975 -57
<< polycont >>
rect -967 40 967 57
rect -967 -57 967 -40
<< locali >>
rect -1055 91 -1007 108
rect 1007 91 1055 108
rect -1055 60 -1038 91
rect 1038 60 1055 91
rect -975 40 -967 57
rect 967 40 975 57
rect -998 15 -981 23
rect -998 -23 -981 -15
rect 981 15 998 23
rect 981 -23 998 -15
rect -975 -57 -967 -40
rect 967 -57 975 -40
rect -1055 -91 -1038 -60
rect 1038 -91 1055 -60
rect -1055 -108 -1007 -91
rect 1007 -108 1055 -91
<< viali >>
rect -967 40 967 57
rect -998 -15 -981 15
rect 981 -15 998 15
rect -967 -57 967 -40
<< metal1 >>
rect -973 57 973 60
rect -973 40 -967 57
rect 967 40 973 57
rect -973 37 973 40
rect -1001 15 -978 21
rect -1001 -15 -998 15
rect -981 -15 -978 15
rect -1001 -21 -978 -15
rect 978 15 1001 21
rect 978 -15 981 15
rect 998 -15 1001 15
rect 978 -21 1001 -15
rect -973 -40 973 -37
rect -973 -57 -967 -40
rect 967 -57 973 -40
rect -973 -60 973 -57
<< properties >>
string FIXED_BBOX -1046 -99 1046 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 19.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
