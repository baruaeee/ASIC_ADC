magic
tech sky130A
magscale 1 2
timestamp 1704374400
<< pwell >>
rect -263 -252 263 252
<< nmos >>
rect -67 -42 67 42
<< ndiff >>
rect -125 30 -67 42
rect -125 -30 -113 30
rect -79 -30 -67 30
rect -125 -42 -67 -30
rect 67 30 125 42
rect 67 -30 79 30
rect 113 -30 125 30
rect 67 -42 125 -30
<< ndiffc >>
rect -113 -30 -79 30
rect 79 -30 113 30
<< psubdiff >>
rect -227 182 -131 216
rect 131 182 227 216
rect -227 120 -193 182
rect 193 120 227 182
rect -227 -182 -193 -120
rect 193 -182 227 -120
rect -227 -216 -131 -182
rect 131 -216 227 -182
<< psubdiffcont >>
rect -131 182 131 216
rect -227 -120 -193 120
rect 193 -120 227 120
rect -131 -216 131 -182
<< poly >>
rect -67 114 67 130
rect -67 80 -51 114
rect 51 80 67 114
rect -67 42 67 80
rect -67 -80 67 -42
rect -67 -114 -51 -80
rect 51 -114 67 -80
rect -67 -130 67 -114
<< polycont >>
rect -51 80 51 114
rect -51 -114 51 -80
<< locali >>
rect -227 182 -131 216
rect 131 182 227 216
rect -227 120 -193 182
rect 193 120 227 182
rect -67 80 -51 114
rect 51 80 67 114
rect -113 30 -79 46
rect -113 -46 -79 -30
rect 79 30 113 46
rect 79 -46 113 -30
rect -67 -114 -51 -80
rect 51 -114 67 -80
rect -227 -182 -193 -120
rect 193 -182 227 -120
rect -227 -216 -131 -182
rect 131 -216 227 -182
<< viali >>
rect -51 80 51 114
rect -113 -30 -79 30
rect 79 -30 113 30
rect -51 -114 51 -80
<< metal1 >>
rect -63 114 63 120
rect -63 80 -51 114
rect 51 80 63 114
rect -63 74 63 80
rect -119 30 -73 42
rect -119 -30 -113 30
rect -79 -30 -73 30
rect -119 -42 -73 -30
rect 73 30 119 42
rect 73 -30 79 30
rect 113 -30 119 30
rect 73 -42 119 -30
rect -63 -80 63 -74
rect -63 -114 -51 -80
rect 51 -114 63 -80
rect -63 -120 63 -114
<< properties >>
string FIXED_BBOX -210 -199 210 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.67 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
