magic
tech sky130A
magscale 1 2
timestamp 1706216322
<< error_p >>
rect -29 182 29 188
rect -29 148 -17 182
rect -29 142 29 148
rect -29 -148 29 -142
rect -29 -182 -17 -148
rect -29 -188 29 -182
<< pwell >>
rect -211 -320 211 320
<< nmos >>
rect -15 -110 15 110
<< ndiff >>
rect -73 98 -15 110
rect -73 -98 -61 98
rect -27 -98 -15 98
rect -73 -110 -15 -98
rect 15 98 73 110
rect 15 -98 27 98
rect 61 -98 73 98
rect 15 -110 73 -98
<< ndiffc >>
rect -61 -98 -27 98
rect 27 -98 61 98
<< psubdiff >>
rect -175 188 -141 250
rect -175 -250 -141 -188
<< psubdiffcont >>
rect -175 -188 -141 188
<< poly >>
rect -33 182 33 198
rect -33 148 -17 182
rect 17 148 33 182
rect -33 132 33 148
rect -15 110 15 132
rect -15 -132 15 -110
rect -33 -148 33 -132
rect -33 -182 -17 -148
rect 17 -182 33 -148
rect -33 -198 33 -182
<< polycont >>
rect -17 148 17 182
rect -17 -182 17 -148
<< locali >>
rect -175 188 -141 250
rect -33 148 -17 182
rect 17 148 33 182
rect -61 98 -27 114
rect -61 -114 -27 -98
rect 27 98 61 114
rect 27 -114 61 -98
rect -33 -182 -17 -148
rect 17 -182 33 -148
rect -175 -250 -141 -188
<< viali >>
rect -17 148 17 182
rect -61 -98 -27 98
rect 27 -98 61 98
rect -17 -182 17 -148
<< metal1 >>
rect -29 182 29 188
rect -29 148 -17 182
rect 17 148 29 182
rect -29 142 29 148
rect -67 98 -21 110
rect -67 -98 -61 98
rect -27 -98 -21 98
rect -67 -110 -21 -98
rect 21 98 67 110
rect 21 -98 27 98
rect 61 -98 67 98
rect 21 -110 67 -98
rect -29 -148 29 -142
rect -29 -182 -17 -148
rect 17 -182 29 -148
rect -29 -188 29 -182
<< properties >>
string FIXED_BBOX -158 -267 158 267
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.1 l 0.153 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
