VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
  MACRO oaTaper STRING ;
END PROPERTYDEFINITIONS

MACRO pre_therm
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN pre_therm 0 0 ;
  SIZE 11.935 BY 13.98 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y01
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.71 8.205 3.21 8.535 ;
        RECT 2.985 5.51 3.21 8.535 ;
        RECT 2.69 5.51 3.21 6.2 ;
      LAYER met2 ;
        RECT 2.105 8.215 2.97 8.535 ;
        RECT 0.135 14.4 2.365 14.66 ;
        RECT 2.105 8.215 2.365 14.66 ;
        RECT 0 14.825 0.5 15.325 ;
        RECT 0.135 14.4 0.395 15.325 ;
      LAYER via ;
        RECT 2.765 8.3 2.915 8.45 ;
    END
  END Y01
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
        RECT 11.21 4.47 11.93 4.85 ;
        RECT 11.2 4.495 11.93 4.825 ;
        RECT 11.21 13.79 11.93 14.17 ;
        RECT 11.2 13.815 11.93 14.145 ;
        RECT 2.475 4.485 3.205 4.815 ;
        RECT 2.475 4.465 3.195 4.845 ;
        RECT 0.775 13.81 1.505 14.14 ;
        RECT 0.78 13.785 1.5 14.165 ;
      LAYER met1 ;
        RECT 0 4.4 11.935 4.92 ;
        RECT 10.36 4.4 11.74 5.12 ;
        RECT 8.7 4.2 10.08 4.92 ;
        RECT 8.665 4.4 10.045 5.12 ;
        RECT 6.97 4.4 8.35 5.12 ;
        RECT 6.96 4.2 8.34 4.92 ;
        RECT 5.22 4.2 6.6 5.12 ;
        RECT 3.48 4.2 4.86 5.12 ;
        RECT 1.74 4.2 3.12 5.12 ;
        RECT 0 4.195 1.38 5.12 ;
        RECT -0.125 7.54 0.245 8.59 ;
        RECT -0.125 4.68 0.075 8.59 ;
        RECT 0 13.72 11.935 14.24 ;
        RECT 7.43 13.715 10.44 14.24 ;
        RECT 9.06 13.52 10.44 14.24 ;
        RECT 7.43 13.52 8.81 14.24 ;
        RECT 5.735 13.525 7.115 14.24 ;
        RECT 4.04 13.525 5.42 14.24 ;
      LAYER met2 ;
        RECT 11.225 4.475 11.905 4.845 ;
        RECT 11.225 13.795 11.905 14.165 ;
        RECT 2.5 4.465 3.18 4.835 ;
        RECT 0.8 13.79 1.48 14.16 ;
      LAYER met4 ;
        RECT 11.545 4.4 11.935 14.24 ;
        RECT 11.205 13.815 11.935 14.145 ;
        RECT 11.205 4.495 11.935 4.825 ;
        RECT 1.595 4.4 3.24 4.915 ;
        RECT 0.715 13.72 1.98 14.24 ;
        RECT 1.59 4.915 1.98 14.24 ;
      LAYER via ;
        RECT 0.91 13.895 1.06 14.045 ;
        RECT 1.23 13.895 1.38 14.045 ;
        RECT 2.585 4.575 2.735 4.725 ;
        RECT 2.905 4.575 3.055 4.725 ;
        RECT 11.38 13.9 11.53 14.05 ;
        RECT 11.38 4.58 11.53 4.73 ;
        RECT 11.7 13.9 11.85 14.05 ;
        RECT 11.7 4.58 11.85 4.73 ;
      LAYER via2 ;
        RECT 0.84 13.875 1.04 14.075 ;
        RECT 1.24 13.875 1.44 14.075 ;
        RECT 2.54 4.55 2.74 4.75 ;
        RECT 2.94 4.55 3.14 4.75 ;
        RECT 11.265 13.88 11.465 14.08 ;
        RECT 11.265 4.56 11.465 4.76 ;
        RECT 11.665 13.88 11.865 14.08 ;
        RECT 11.665 4.56 11.865 4.76 ;
      LAYER via3 ;
        RECT 0.84 13.875 1.04 14.075 ;
        RECT 1.24 13.875 1.44 14.075 ;
        RECT 2.535 4.555 2.735 4.755 ;
        RECT 2.935 4.555 3.135 4.755 ;
        RECT 11.27 13.88 11.47 14.08 ;
        RECT 11.27 4.56 11.47 4.76 ;
        RECT 11.67 13.88 11.87 14.08 ;
        RECT 11.67 4.56 11.87 4.76 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
        RECT 10.195 9.155 10.925 9.485 ;
        RECT 10.195 -0.165 10.925 0.165 ;
        RECT 10.365 -0.26 10.755 9.58 ;
        RECT 1.49 -0.165 2.22 0.165 ;
        RECT 1.25 9.14 1.98 9.47 ;
        RECT 1.59 -0.165 1.98 9.47 ;
      LAYER met1 ;
        RECT 0 -0.26 11.935 0.26 ;
        RECT 8.7 -0.26 10.08 0.46 ;
        RECT 6.96 -0.26 8.34 0.46 ;
        RECT 5.22 -0.26 6.6 0.46 ;
        RECT 3.48 -0.26 4.86 0.46 ;
        RECT 1.74 -0.26 3.12 0.46 ;
        RECT 0 -0.26 1.38 0.455 ;
        RECT 0 9.06 11.935 9.58 ;
        RECT 10.36 8.86 11.74 9.58 ;
        RECT 9.06 9.06 10.44 9.78 ;
        RECT 8.665 8.86 10.045 9.58 ;
        RECT 7.43 9.06 8.81 9.78 ;
        RECT 6.97 8.86 8.35 9.58 ;
        RECT 5.735 9.06 7.115 9.785 ;
        RECT 5.22 8.86 6.6 9.58 ;
        RECT 4.04 9.06 5.42 9.785 ;
        RECT 3.48 8.86 4.86 9.58 ;
        RECT 1.74 8.86 3.12 9.58 ;
        RECT 0 8.86 1.38 9.78 ;
        RECT 0.275 8.86 0.505 10.31 ;
      LAYER met2 ;
        RECT 10.22 -0.185 10.9 0.185 ;
        RECT 10.22 9.135 10.9 9.505 ;
        RECT 1.515 -0.185 2.195 0.185 ;
        RECT 1.275 9.12 1.955 9.49 ;
      LAYER via ;
        RECT 1.38 9.225 1.53 9.375 ;
        RECT 1.62 -0.08 1.77 0.07 ;
        RECT 1.7 9.225 1.85 9.375 ;
        RECT 1.94 -0.08 2.09 0.07 ;
        RECT 10.325 9.245 10.475 9.395 ;
        RECT 10.325 -0.075 10.475 0.075 ;
        RECT 10.645 9.245 10.795 9.395 ;
        RECT 10.645 -0.075 10.795 0.075 ;
      LAYER via2 ;
        RECT 1.315 9.205 1.515 9.405 ;
        RECT 1.555 -0.1 1.755 0.1 ;
        RECT 1.715 9.205 1.915 9.405 ;
        RECT 1.955 -0.1 2.155 0.1 ;
        RECT 10.26 9.22 10.46 9.42 ;
        RECT 10.26 -0.1 10.46 0.1 ;
        RECT 10.66 9.22 10.86 9.42 ;
        RECT 10.66 -0.1 10.86 0.1 ;
    END
  END VSS
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.95 2.395 9.32 2.765 ;
        RECT 8.975 2.395 9.295 3.025 ;
        RECT 7.33 2.395 7.7 2.765 ;
        RECT 7.355 2.395 7.675 3.025 ;
        RECT 6.805 6.8 7.175 7.17 ;
        RECT 5.19 7.13 5.56 7.5 ;
        RECT 0.46 1.06 1.015 1.43 ;
        RECT -0.555 1.08 1.015 1.41 ;
        RECT -0.815 1.085 1.015 1.405 ;
        RECT 0.23 6.355 0.6 7.205 ;
        RECT -0.095 11.915 0.345 13.295 ;
      LAYER met2 ;
        RECT -0.815 2.765 9.295 3.025 ;
        RECT 6.855 6.355 7.175 7.06 ;
        RECT -1.655 6.355 7.175 6.61 ;
        RECT 5.19 6.355 5.51 7.39 ;
        RECT -1.655 6.355 0.49 6.675 ;
        RECT -0.815 12.385 0.275 12.705 ;
        RECT -0.815 1.08 -0.555 12.705 ;
        RECT -1.655 6.285 -1.155 6.785 ;
      LAYER via ;
        RECT -0.76 1.17 -0.61 1.32 ;
        RECT 0.07 12.47 0.22 12.62 ;
        RECT 0.285 6.44 0.435 6.59 ;
        RECT 5.275 7.185 5.425 7.335 ;
        RECT 6.94 6.855 7.09 7.005 ;
        RECT 7.44 2.82 7.59 2.97 ;
        RECT 9.06 2.82 9.21 2.97 ;
    END
  END IN
  PIN Y02
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.105 8.045 4.835 8.375 ;
        RECT 4.605 5.47 4.835 8.375 ;
        RECT 4.09 5.47 4.835 6.16 ;
      LAYER met2 ;
        RECT 2.565 8.735 4.365 8.995 ;
        RECT 4.105 8.055 4.365 8.995 ;
        RECT 0.9 14.95 2.825 15.21 ;
        RECT 2.565 8.735 2.825 15.21 ;
        RECT 0.9 14.825 1.4 15.325 ;
      LAYER via ;
        RECT 4.16 8.14 4.31 8.29 ;
    END
  END Y02
  PIN preampF1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.545 1.885 5.915 2.255 ;
        RECT 3.87 1.105 4.24 1.475 ;
        RECT 2.065 1.945 2.435 2.585 ;
        RECT 0.61 1.945 2.435 2.265 ;
        RECT 0.615 1.825 0.84 2.725 ;
        RECT 0.61 1.9 0.84 2.55 ;
      LAYER met2 ;
        RECT 2.105 1.945 5.865 2.205 ;
        RECT 3.87 1.105 4.13 2.205 ;
      LAYER via ;
        RECT 2.19 2 2.34 2.15 ;
        RECT 3.925 1.19 4.075 1.34 ;
        RECT 5.63 2 5.78 2.15 ;
    END
  END preampF1
  PIN Y03
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.45 3.33 3.235 3.955 ;
        RECT 3.005 0.875 3.235 3.955 ;
        RECT 2.505 0.875 3.235 1.565 ;
        RECT 2.45 3.305 2.68 3.955 ;
      LAYER met2 ;
        RECT 2.455 -1.785 2.955 -1.285 ;
        RECT 2.575 -1.785 2.835 1.195 ;
      LAYER via ;
        RECT 2.63 0.96 2.78 1.11 ;
    END
  END Y03
  PIN Y04
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.075 2.875 4.955 3.565 ;
        RECT 4.725 0.985 4.955 3.565 ;
        RECT 4.39 0.985 4.955 1.675 ;
      LAYER met2 ;
        RECT 4.275 -1.785 4.775 -1.285 ;
        RECT 4.39 -1.785 4.65 1.305 ;
      LAYER via ;
        RECT 4.445 1.07 4.595 1.22 ;
    END
  END Y04
  PIN Y05
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.755 3.085 6.525 3.775 ;
        RECT 6.295 0.875 6.525 3.775 ;
        RECT 5.96 0.875 6.525 1.565 ;
      LAYER met2 ;
        RECT 5.845 -1.785 6.345 -1.285 ;
        RECT 5.96 -1.785 6.22 1.305 ;
      LAYER via ;
        RECT 6.015 1.07 6.165 1.22 ;
    END
  END Y05
  PIN Y06
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.755 3.38 8.4 3.71 ;
        RECT 8.17 0.95 8.4 3.71 ;
        RECT 7.7 0.95 8.4 1.64 ;
      LAYER met2 ;
        RECT 7.58 -1.785 8.08 -1.285 ;
        RECT 7.7 -1.785 7.96 1.305 ;
      LAYER via ;
        RECT 7.755 1.07 7.905 1.22 ;
    END
  END Y06
  PIN Y07
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 9.24 3.33 10.04 3.66 ;
        RECT 9.81 0.855 10.04 3.66 ;
        RECT 9.34 0.855 10.04 1.545 ;
      LAYER met2 ;
        RECT 9.22 -1.785 9.72 -1.285 ;
        RECT 9.34 -1.785 9.6 1.305 ;
      LAYER via ;
        RECT 9.395 1.07 9.545 1.22 ;
    END
  END Y07
  PIN Y08
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.09 5.545 6.42 7.305 ;
        RECT 5.77 5.545 6.42 6.235 ;
      LAYER met2 ;
        RECT 3.025 9.195 6.375 9.455 ;
        RECT 6.115 6.94 6.375 9.455 ;
        RECT 3.025 14.825 3.525 15.325 ;
        RECT 3.025 9.195 3.285 15.325 ;
      LAYER via ;
        RECT 6.17 7.025 6.32 7.175 ;
    END
  END Y08
  PIN Y09
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.475 6.61 8.405 6.87 ;
        RECT 7.475 6.61 7.805 7.24 ;
        RECT 7.545 5.67 7.775 7.24 ;
      LAYER met2 ;
        RECT 3.485 9.655 7.765 9.915 ;
        RECT 7.505 6.92 7.765 9.915 ;
        RECT 3.87 14.825 4.37 15.325 ;
        RECT 3.99 14.365 4.25 15.325 ;
        RECT 3.485 14.365 4.25 14.625 ;
        RECT 3.485 9.655 3.745 14.625 ;
      LAYER via ;
        RECT 7.56 7.005 7.71 7.155 ;
    END
  END Y09
  PIN Y10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.695 12.33 5.395 13.02 ;
        RECT 5.135 10.275 5.395 13.02 ;
        RECT 4.645 10.275 5.395 10.965 ;
      LAYER met2 ;
        RECT 4.905 14.825 5.405 15.325 ;
        RECT 5.025 12.7 5.285 15.325 ;
      LAYER via ;
        RECT 5.08 12.785 5.23 12.935 ;
    END
  END Y10
  PIN Y11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.37 12.285 7.185 12.975 ;
        RECT 6.925 10.33 7.185 12.975 ;
      LAYER met2 ;
        RECT 6.24 14.825 6.74 15.325 ;
        RECT 6.37 12.655 6.63 15.325 ;
      LAYER via ;
        RECT 6.425 12.74 6.575 12.89 ;
    END
  END Y11
  PIN Y12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.99 12.405 8.615 13.095 ;
        RECT 8.355 10.2 8.615 13.095 ;
        RECT 8.125 10.2 8.615 10.89 ;
      LAYER met2 ;
        RECT 7.86 14.825 8.36 15.325 ;
        RECT 7.99 12.655 8.25 15.325 ;
      LAYER via ;
        RECT 8.045 12.74 8.195 12.89 ;
    END
  END Y12
  PIN Y13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 9.63 12.355 10.225 13.045 ;
        RECT 9.995 10.3 10.225 13.045 ;
      LAYER met2 ;
        RECT 9.5 14.825 10 15.325 ;
        RECT 9.63 12.655 9.89 15.325 ;
      LAYER via ;
        RECT 9.685 12.74 9.835 12.89 ;
    END
  END Y13
  PIN Y14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 9.715 8.02 9.975 8.34 ;
        RECT 9.715 5.62 9.945 8.34 ;
        RECT 9.285 5.62 9.945 6.31 ;
      LAYER met2 ;
        RECT 12.64 10.52 13.14 11.02 ;
        RECT 9.715 10.655 13.14 10.915 ;
        RECT 9.715 8.02 9.975 10.915 ;
      LAYER via ;
        RECT 9.77 8.105 9.92 8.255 ;
    END
  END Y14
  PIN Y15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 11.55 7.21 11.87 7.47 ;
        RECT 11.55 5.645 11.81 8.315 ;
        RECT 11.155 5.645 11.81 6.335 ;
      LAYER met2 ;
        RECT 12.64 7.1 13.14 7.6 ;
        RECT 11.55 7.21 13.14 7.47 ;
      LAYER via ;
        RECT 11.635 7.265 11.785 7.415 ;
    END
  END Y15
  OBS
    LAYER mcon ;
      RECT 11.58 8.065 11.75 8.235 ;
      RECT 11.195 4.835 11.365 5.005 ;
      RECT 11.195 8.975 11.365 9.145 ;
      RECT 11.185 5.725 11.355 5.895 ;
      RECT 11.185 6.085 11.355 6.255 ;
      RECT 10.975 7.21 11.145 7.38 ;
      RECT 10.735 4.835 10.905 5.005 ;
      RECT 10.735 8.975 10.905 9.145 ;
      RECT 10.025 10.41 10.195 10.58 ;
      RECT 9.895 9.495 10.065 9.665 ;
      RECT 9.895 13.635 10.065 13.805 ;
      RECT 9.745 8.06 9.915 8.23 ;
      RECT 9.66 12.435 9.83 12.605 ;
      RECT 9.66 12.795 9.83 12.965 ;
      RECT 9.535 0.175 9.705 0.345 ;
      RECT 9.535 4.315 9.705 4.485 ;
      RECT 9.5 4.835 9.67 5.005 ;
      RECT 9.5 8.975 9.67 9.145 ;
      RECT 9.44 11.285 9.61 11.455 ;
      RECT 9.435 9.495 9.605 9.665 ;
      RECT 9.435 13.635 9.605 13.805 ;
      RECT 9.37 0.935 9.54 1.105 ;
      RECT 9.37 1.295 9.54 1.465 ;
      RECT 9.315 5.7 9.485 5.87 ;
      RECT 9.315 6.06 9.485 6.23 ;
      RECT 9.27 3.41 9.44 3.58 ;
      RECT 9.1 7.23 9.27 7.4 ;
      RECT 9.075 0.175 9.245 0.345 ;
      RECT 9.075 4.315 9.245 4.485 ;
      RECT 9.05 2.495 9.22 2.665 ;
      RECT 9.04 4.835 9.21 5.005 ;
      RECT 9.04 8.975 9.21 9.145 ;
      RECT 8.265 9.495 8.435 9.665 ;
      RECT 8.265 13.635 8.435 13.805 ;
      RECT 8.155 10.28 8.325 10.45 ;
      RECT 8.155 10.64 8.325 10.81 ;
      RECT 8.02 12.465 8.19 12.635 ;
      RECT 8.02 12.825 8.19 12.995 ;
      RECT 7.81 11.68 7.98 11.85 ;
      RECT 7.805 4.835 7.975 5.005 ;
      RECT 7.805 8.975 7.975 9.145 ;
      RECT 7.805 9.495 7.975 9.665 ;
      RECT 7.805 13.635 7.975 13.805 ;
      RECT 7.795 0.175 7.965 0.345 ;
      RECT 7.795 4.315 7.965 4.485 ;
      RECT 7.785 3.46 7.955 3.63 ;
      RECT 7.73 1.03 7.9 1.2 ;
      RECT 7.73 1.39 7.9 1.56 ;
      RECT 7.575 5.75 7.745 5.92 ;
      RECT 7.555 7.04 7.725 7.21 ;
      RECT 7.43 2.495 7.6 2.665 ;
      RECT 7.345 4.835 7.515 5.005 ;
      RECT 7.345 8.975 7.515 9.145 ;
      RECT 7.335 0.175 7.505 0.345 ;
      RECT 7.335 4.315 7.505 4.485 ;
      RECT 6.955 10.41 7.125 10.58 ;
      RECT 6.905 6.9 7.075 7.07 ;
      RECT 6.57 9.5 6.74 9.67 ;
      RECT 6.57 13.64 6.74 13.81 ;
      RECT 6.4 12.365 6.57 12.535 ;
      RECT 6.4 12.725 6.57 12.895 ;
      RECT 6.17 7.105 6.34 7.275 ;
      RECT 6.13 11.265 6.3 11.435 ;
      RECT 6.11 9.5 6.28 9.67 ;
      RECT 6.11 13.64 6.28 13.81 ;
      RECT 6.055 0.175 6.225 0.345 ;
      RECT 6.055 4.315 6.225 4.485 ;
      RECT 6.055 4.835 6.225 5.005 ;
      RECT 6.055 8.975 6.225 9.145 ;
      RECT 5.99 0.955 6.16 1.125 ;
      RECT 5.99 1.315 6.16 1.485 ;
      RECT 5.8 5.625 5.97 5.795 ;
      RECT 5.8 5.985 5.97 6.155 ;
      RECT 5.785 3.165 5.955 3.335 ;
      RECT 5.785 3.525 5.955 3.695 ;
      RECT 5.645 1.985 5.815 2.155 ;
      RECT 5.595 0.175 5.765 0.345 ;
      RECT 5.595 4.315 5.765 4.485 ;
      RECT 5.595 4.835 5.765 5.005 ;
      RECT 5.595 8.975 5.765 9.145 ;
      RECT 5.29 7.23 5.46 7.4 ;
      RECT 4.875 9.5 5.045 9.67 ;
      RECT 4.875 13.64 5.045 13.81 ;
      RECT 4.725 12.41 4.895 12.58 ;
      RECT 4.725 12.77 4.895 12.94 ;
      RECT 4.675 10.355 4.845 10.525 ;
      RECT 4.675 10.715 4.845 10.885 ;
      RECT 4.455 11.36 4.625 11.53 ;
      RECT 4.42 1.065 4.59 1.235 ;
      RECT 4.42 1.425 4.59 1.595 ;
      RECT 4.415 9.5 4.585 9.67 ;
      RECT 4.415 13.64 4.585 13.81 ;
      RECT 4.315 0.175 4.485 0.345 ;
      RECT 4.315 4.315 4.485 4.485 ;
      RECT 4.315 4.835 4.485 5.005 ;
      RECT 4.315 8.975 4.485 9.145 ;
      RECT 4.135 8.125 4.305 8.295 ;
      RECT 4.12 5.55 4.29 5.72 ;
      RECT 4.12 5.91 4.29 6.08 ;
      RECT 4.105 2.955 4.275 3.125 ;
      RECT 4.105 3.315 4.275 3.485 ;
      RECT 3.97 1.205 4.14 1.375 ;
      RECT 3.855 0.175 4.025 0.345 ;
      RECT 3.855 4.315 4.025 4.485 ;
      RECT 3.855 4.835 4.025 5.005 ;
      RECT 3.855 7.345 4.025 7.515 ;
      RECT 3.855 8.975 4.025 9.145 ;
      RECT 2.74 8.28 2.91 8.45 ;
      RECT 2.72 5.59 2.89 5.76 ;
      RECT 2.72 5.95 2.89 6.12 ;
      RECT 2.575 0.175 2.745 0.345 ;
      RECT 2.575 4.315 2.745 4.485 ;
      RECT 2.575 4.835 2.745 5.005 ;
      RECT 2.575 8.975 2.745 9.145 ;
      RECT 2.535 0.955 2.705 1.125 ;
      RECT 2.535 1.315 2.705 1.485 ;
      RECT 2.48 3.365 2.65 3.535 ;
      RECT 2.48 3.725 2.65 3.895 ;
      RECT 2.23 7.345 2.4 7.515 ;
      RECT 2.165 2.045 2.335 2.215 ;
      RECT 2.115 0.175 2.285 0.345 ;
      RECT 2.115 4.315 2.285 4.485 ;
      RECT 2.115 4.835 2.285 5.005 ;
      RECT 2.115 8.975 2.285 9.145 ;
      RECT 1.265 12.185 1.435 12.355 ;
      RECT 1.015 5.405 1.185 5.575 ;
      RECT 0.835 0.17 1.005 0.34 ;
      RECT 0.835 4.31 1.005 4.48 ;
      RECT 0.835 4.835 1.005 5.005 ;
      RECT 0.835 8.975 1.005 9.145 ;
      RECT 0.835 9.495 1.005 9.665 ;
      RECT 0.725 1.16 0.895 1.33 ;
      RECT 0.64 1.96 0.81 2.13 ;
      RECT 0.64 2.32 0.81 2.49 ;
      RECT 0.525 10.705 0.695 10.875 ;
      RECT 0.525 11.065 0.695 11.235 ;
      RECT 0.485 7.62 0.655 7.79 ;
      RECT 0.485 7.98 0.655 8.15 ;
      RECT 0.485 8.34 0.655 8.51 ;
      RECT 0.375 0.17 0.545 0.34 ;
      RECT 0.375 4.31 0.545 4.48 ;
      RECT 0.375 4.835 0.545 5.005 ;
      RECT 0.375 8.975 0.545 9.145 ;
      RECT 0.375 9.495 0.545 9.665 ;
      RECT 0.33 6.84 0.5 7.01 ;
      RECT 0.305 10.08 0.475 10.25 ;
      RECT 0.06 12.29 0.23 12.46 ;
      RECT 0.06 12.75 0.23 12.92 ;
      RECT 0.045 7.62 0.215 7.79 ;
      RECT 0.045 7.98 0.215 8.15 ;
      RECT 0.045 8.34 0.215 8.51 ;
    LAYER met1 ;
      RECT 10.875 7.11 11.135 7.5 ;
      RECT 10.875 7.11 11.245 7.48 ;
      RECT 7.71 11.58 8.08 11.95 ;
      RECT 7.71 11.26 8.03 11.95 ;
      RECT 1.185 10.625 1.515 12.385 ;
      RECT 1.185 11.26 4.725 11.63 ;
      RECT 0.495 10.625 1.515 11.315 ;
      RECT 0.455 7.54 1.245 8.59 ;
      RECT 0.955 5.375 1.245 8.59 ;
      RECT 9.34 11.185 9.71 11.555 ;
      RECT 9 7.13 9.37 7.5 ;
      RECT 6.03 11.165 6.4 11.535 ;
      RECT 3.755 6.86 4.125 7.71 ;
      RECT 2.13 6.86 2.5 7.71 ;
    LAYER via ;
      RECT 10.93 7.265 11.08 7.415 ;
      RECT 9.425 11.315 9.575 11.465 ;
      RECT 9.055 7.265 9.205 7.415 ;
      RECT 7.795 11.315 7.945 11.465 ;
      RECT 6.115 11.315 6.265 11.465 ;
      RECT 4.49 11.315 4.64 11.465 ;
      RECT 3.81 7.475 3.96 7.625 ;
      RECT 2.185 7.475 2.335 7.625 ;
      RECT 1.02 7.475 1.17 7.625 ;
    LAYER met2 ;
      RECT 4.405 11.26 9.66 11.52 ;
      RECT 9 7.18 9.26 11.52 ;
      RECT 9 7.18 11.135 7.5 ;
      RECT 0.965 7.39 4.015 7.71 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END pre_therm

END LIBRARY
