* NGSPICE file created from th01.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_SHU4BF a_n73_n353# a_n141_493# a_15_n353# a_n33_n441#
X0 a_15_n353# a_n33_n441# a_n73_n353# a_n141_493# sky130_fd_pr__nfet_01v8 ad=1.02 pd=7.64 as=1.02 ps=7.64 w=3.53 l=0.15
C0 a_15_n353# a_n33_n441# 0.0384f
C1 a_15_n353# a_n73_n353# 0.564f
C2 a_n33_n441# a_n73_n353# 0.0384f
C3 a_15_n353# a_n141_493# 0.327f
C4 a_n73_n353# a_n141_493# 0.327f
C5 a_n33_n441# a_n141_493# 0.329f
.ends

.subckt sky130_fd_pr__pfet_01v8_HE9GT9 a_n408_n42# a_350_n42# w_n546_n261# a_n350_n139#
+ VSUBS
X0 a_350_n42# a_n350_n139# a_n408_n42# w_n546_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 a_n408_n42# w_n546_n261# 0.0408f
C1 a_350_n42# w_n546_n261# 0.0179f
C2 a_n408_n42# a_n350_n139# 0.0226f
C3 a_350_n42# a_n350_n139# 0.0226f
C4 a_n408_n42# a_350_n42# 0.00807f
C5 w_n546_n261# a_n350_n139# 0.756f
C6 a_350_n42# VSUBS 0.0587f
C7 a_n408_n42# VSUBS 0.0437f
C8 a_n350_n139# VSUBS 1.19f
C9 w_n546_n261# VSUBS 1.83f
.ends

.subckt sky130_fd_pr__nfet_01v8_LHD8GA a_n408_n42# a_350_n42# a_n350_n130# a_n510_n182#
X0 a_350_n42# a_n350_n130# a_n408_n42# a_n510_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 a_350_n42# a_n350_n130# 0.0226f
C1 a_350_n42# a_n408_n42# 0.00807f
C2 a_n350_n130# a_n408_n42# 0.0226f
C3 a_350_n42# a_n510_n182# 0.0766f
C4 a_n408_n42# a_n510_n182# 0.0845f
C5 a_n350_n130# a_n510_n182# 1.9f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJP3BL a_15_n150# w_n211_n369# a_n73_n150# a_n33_n247#
+ VSUBS
X0 a_15_n150# a_n33_n247# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.15
C0 a_n73_n150# w_n211_n369# 0.0292f
C1 a_15_n150# w_n211_n369# 0.0292f
C2 a_n73_n150# a_n33_n247# 0.0267f
C3 a_15_n150# a_n33_n247# 0.0267f
C4 a_n73_n150# a_15_n150# 0.242f
C5 w_n211_n369# a_n33_n247# 0.19f
C6 a_15_n150# VSUBS 0.126f
C7 a_n73_n150# VSUBS 0.126f
C8 a_n33_n247# VSUBS 0.146f
C9 w_n211_n369# VSUBS 1.02f
.ends

.subckt sky130_fd_pr__nfet_01v8_LH5FDA a_n150_n130# a_276_n182# a_n208_n42# a_150_n42#
X0 a_150_n42# a_n150_n130# a_n208_n42# a_276_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.5
C0 a_150_n42# a_n150_n130# 0.0176f
C1 a_150_n42# a_n208_n42# 0.0172f
C2 a_n150_n130# a_n208_n42# 0.0176f
C3 a_150_n42# a_276_n182# 0.0815f
C4 a_n208_n42# a_276_n182# 0.0736f
C5 a_n150_n130# a_276_n182# 0.904f
.ends

.subckt th01 Vp Vin V01 Vn
XXM0 Vn Vn m1_991_n1219# Vin sky130_fd_pr__nfet_01v8_SHU4BF
XXM1 m1_571_n501# m1_991_n1219# Vp Vin Vn sky130_fd_pr__pfet_01v8_HE9GT9
XXM2 Vp m1_571_n501# Vp Vn sky130_fd_pr__nfet_01v8_LHD8GA
XXM3 Vp Vp V01 m1_991_n1219# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_991_n1219# Vn V01 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 m1_571_n501# V01 2.16e-20
C1 m1_991_n1219# Vp 0.423f
C2 Vin m1_991_n1219# 0.208f
C3 Vin Vp 0.354f
C4 m1_571_n501# m1_991_n1219# 0.0899f
C5 m1_571_n501# Vp 0.32f
C6 m1_571_n501# Vin 0.274f
C7 V01 m1_991_n1219# 0.0901f
C8 V01 Vp 0.0684f
C9 Vin V01 0.00412f
C10 V01 Vn 0.388f
C11 m1_991_n1219# Vn 1.3f
C12 m1_571_n501# Vn 0.194f
C13 Vin Vn 1.93f
C14 Vp Vn 4.44f
.ends

