magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_s >>
rect 362 1008 397 1026
rect 362 999 433 1008
rect 363 972 433 999
rect 749 977 802 1008
rect 380 938 451 972
rect 749 943 820 977
rect 380 583 450 938
rect 562 870 620 876
rect 562 836 574 870
rect 562 830 620 836
rect 562 666 620 672
rect 562 632 574 666
rect 562 626 620 632
rect 380 547 433 583
rect 749 530 819 943
rect 1101 892 1135 910
rect 931 875 989 881
rect 931 841 943 875
rect 1101 856 1171 892
rect 931 835 989 841
rect 1118 822 1189 856
rect 931 613 989 619
rect 931 579 943 613
rect 931 573 989 579
rect 749 494 802 530
rect 1118 477 1188 822
rect 1118 441 1171 477
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_M6KFPY  XM1
timestamp 1703732895
transform 1 0 960 0 1 727
box -211 -286 211 286
use sky130_fd_pr__nfet_01v8_LNCAWD  XM3
timestamp 1703732895
transform 1 0 1381 0 1 640
box -263 -252 263 252
use sky130_fd_pr__pfet_01v8_NZD9V2  XM7
timestamp 1703732895
transform 1 0 190 0 1 808
box -243 -261 243 261
use sky130_fd_pr__nfet_01v8_NCP4B2  XM10
timestamp 1703732895
transform 1 0 591 0 1 751
box -211 -257 211 257
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
