* NGSPICE file created from op-amp.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_FM7VE8 a_n35_n1932# a_n165_n2062# a_n35_1500#
X0 a_n35_1500# a_n35_n1932# a_n165_n2062# sky130_fd_pr__res_xhigh_po_0p35 l=15
C0 a_n35_n1932# a_n165_n2062# 0.598f
C1 a_n35_1500# a_n165_n2062# 0.598f
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_7RFGLT a_n165_n1062# a_n35_500# a_n35_n932#
X0 a_n35_500# a_n35_n932# a_n165_n1062# sky130_fd_pr__res_xhigh_po_0p35 l=5
C0 a_n35_500# a_n35_n932# 0.00382f
C1 a_n35_n932# a_n165_n1062# 0.593f
C2 a_n35_500# a_n165_n1062# 0.593f
.ends

.subckt sky130_fd_pr__nfet_01v8_69TQ3K a_n260_n274# a_100_n100# a_n158_n100# a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n260_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_n158_n100# a_100_n100# 0.0556f
C1 a_n158_n100# a_n100_n188# 0.0268f
C2 a_n100_n188# a_100_n100# 0.0268f
C3 a_100_n100# a_n260_n274# 0.146f
C4 a_n158_n100# a_n260_n274# 0.146f
C5 a_n100_n188# a_n260_n274# 0.724f
.ends

.subckt sky130_fd_pr__pfet_01v8_3HMWVM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
+ VSUBS
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_n100_n197# a_100_n100# 0.0268f
C1 a_n100_n197# a_n158_n100# 0.0268f
C2 a_n100_n197# w_n296_n319# 0.434f
C3 a_100_n100# a_n158_n100# 0.0556f
C4 w_n296_n319# a_100_n100# 0.0852f
C5 w_n296_n319# a_n158_n100# 0.0852f
C6 a_100_n100# VSUBS 0.0607f
C7 a_n158_n100# VSUBS 0.0607f
C8 a_n100_n197# VSUBS 0.311f
C9 w_n296_n319# VSUBS 1.65f
.ends

.subckt sky130_fd_pr__nfet_01v8_PSFW3M a_n88_n100# a_n33_n188# a_n190_n274# a_30_n100#
X0 a_30_n100# a_n33_n188# a_n88_n100# a_n190_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n88_n100# a_30_n100# 0.121f
C1 a_n88_n100# a_n33_n188# 0.0111f
C2 a_n33_n188# a_30_n100# 0.0111f
C3 a_30_n100# a_n190_n274# 0.139f
C4 a_n88_n100# a_n190_n274# 0.139f
C5 a_n33_n188# a_n190_n274# 0.346f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_FJFAMD m3_n386_n240# c1_n346_n200# VSUBS
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 c1_n346_n200# m3_n386_n240# 0.507f
C1 c1_n346_n200# VSUBS 0.17f
C2 m3_n386_n240# VSUBS 0.763f
.ends

.subckt op-amp Vp vin Vout Vn
XXR1 Vout Vn m1_109_n237# sky130_fd_pr__res_xhigh_po_0p35_FM7VE8
XXR2 Vn m1_109_n237# Vn sky130_fd_pr__res_xhigh_po_0p35_7RFGLT
XXR3 Vp Vn m1_n55_181# sky130_fd_pr__res_xhigh_po_0p35_FM7VE8
XXM1 Vn Vn m1_2069_183# m1_1581_69# sky130_fd_pr__nfet_01v8_69TQ3K
XXM2 m1_924_890# m1_109_n237# m1_1581_69# m1_924_890# Vn sky130_fd_pr__pfet_01v8_3HMWVM
XXM3 Vn m1_1581_69# Vn m1_1581_69# sky130_fd_pr__nfet_01v8_69TQ3K
XXM4 m1_924_890# vin m1_924_890# m1_2069_183# Vn sky130_fd_pr__pfet_01v8_3HMWVM
XXM5 Vp m1_155_757# m1_924_890# Vp Vn sky130_fd_pr__pfet_01v8_3HMWVM
XXM6 m1_2069_183# Vp Vn m1_2801_185# sky130_fd_pr__nfet_01v8_PSFW3M
XXM7 Vp m1_155_757# Vout Vp Vn sky130_fd_pr__pfet_01v8_3HMWVM
XXM9 Vp m1_155_757# m1_155_757# Vp Vn sky130_fd_pr__pfet_01v8_3HMWVM
XXM8 Vn Vout Vn m1_2069_183# sky130_fd_pr__nfet_01v8_69TQ3K
XXC1 Vout m1_2801_185# Vn sky130_fd_pr__cap_mim_m3_1_FJFAMD
XXM10 Vn m1_155_757# Vn m1_n55_181# sky130_fd_pr__nfet_01v8_69TQ3K
XXM11 Vn Vn m1_n55_181# m1_n55_181# sky130_fd_pr__nfet_01v8_69TQ3K
C0 vin m1_155_757# 0.0746f
C1 Vp m1_2069_183# 0.164f
C2 Vp Vn 0.969f
C3 m1_1581_69# m1_2069_183# 0.271f
C4 m1_1581_69# Vn 0.486f
C5 m1_109_n237# m1_2069_183# 3.07e-19
C6 m1_109_n237# Vn 1.03f
C7 Vout m1_155_757# 0.0582f
C8 m1_n55_181# m1_155_757# 0.334f
C9 Vn m1_2069_183# 0.454f
C10 m1_155_757# Vp 0.801f
C11 m1_1581_69# m1_155_757# 0.0687f
C12 vin m1_924_890# 0.243f
C13 m1_109_n237# m1_155_757# 0.158f
C14 m1_155_757# m1_2069_183# 0.123f
C15 m1_155_757# Vn 0.264f
C16 m1_2801_185# Vout 0.583f
C17 Vout m1_924_890# 0.00373f
C18 m1_n55_181# m1_924_890# 8.44e-20
C19 m1_2801_185# Vp 0.0455f
C20 Vp m1_924_890# 0.844f
C21 Vout vin 0.00109f
C22 m1_2801_185# m1_1581_69# 7.35e-20
C23 m1_1581_69# m1_924_890# 0.129f
C24 m1_2801_185# m1_109_n237# 6.67e-20
C25 m1_109_n237# m1_924_890# 0.238f
C26 vin Vp 0.108f
C27 m1_2801_185# m1_2069_183# 0.017f
C28 m1_924_890# m1_2069_183# 0.114f
C29 vin m1_1581_69# 0.0119f
C30 m1_2801_185# Vn 0.274f
C31 m1_924_890# Vn 0.423f
C32 m1_109_n237# vin 0.0127f
C33 Vout Vp 0.171f
C34 vin m1_2069_183# 0.186f
C35 m1_n55_181# Vp 0.489f
C36 vin Vn 0.0175f
C37 Vout m1_1581_69# 0.00343f
C38 m1_n55_181# m1_1581_69# 0.00446f
C39 m1_109_n237# Vout 1.13e-20
C40 m1_n55_181# m1_109_n237# 0.0477f
C41 m1_155_757# m1_924_890# 0.429f
C42 m1_1581_69# Vp 0.00755f
C43 Vout m1_2069_183# 0.212f
C44 Vout Vn 0.383f
C45 m1_109_n237# Vp 0.0163f
C46 m1_n55_181# Vn 0.537f
C47 m1_109_n237# m1_1581_69# 0.118f
C48 Vp 0 5.89f
C49 Vn 0 -1.05f
C50 m1_n55_181# 0 2.29f
C51 m1_155_757# 0 1.31f
C52 m1_2801_185# 0 1.37f
C53 m1_2069_183# 0 1.06f
C54 m1_924_890# 0 2.64f
C55 vin 0 0.256f
C56 m1_1581_69# 0 1.4f
C57 Vout 0 2.45f
C58 m1_109_n237# 0 1.8f
.ends

