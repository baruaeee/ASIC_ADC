* NGSPICE file created from adc1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X a_208_47# a_75_199#
+ a_544_297# a_315_47# a_201_297#
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_315_47# VGND 0.00427f
C1 C1 VPWR 0.0146f
C2 a_208_47# A3 3.65e-19
C3 a_544_297# VGND 0.00256f
C4 VPB X 0.0107f
C5 VPWR A3 0.0181f
C6 a_201_297# VGND 0.00403f
C7 VPB A2 0.0376f
C8 a_75_199# A1 0.0696f
C9 B1 A1 0.0716f
C10 a_544_297# X 2.35e-19
C11 a_315_47# A2 0.00335f
C12 a_208_47# a_75_199# 0.0159f
C13 a_201_297# X 0.0131f
C14 C1 VGND 0.0181f
C15 a_75_199# VPWR 0.109f
C16 a_201_297# A2 0.0112f
C17 VGND A3 0.0161f
C18 B1 VPWR 0.0125f
C19 C1 X 5.14e-20
C20 X A3 0.00317f
C21 a_201_297# VPB 0.00186f
C22 A3 A2 0.0747f
C23 a_75_199# VGND 0.362f
C24 B1 VGND 0.0171f
C25 a_201_297# a_544_297# 0.00702f
C26 VPB C1 0.0394f
C27 a_75_199# X 0.0959f
C28 B1 X 7.79e-20
C29 VPB A3 0.0268f
C30 a_75_199# A2 0.0621f
C31 a_201_297# C1 0.00243f
C32 a_201_297# A3 0.00642f
C33 VPB a_75_199# 0.0486f
C34 VPB B1 0.0292f
C35 a_315_47# a_75_199# 0.0202f
C36 a_544_297# a_75_199# 0.0176f
C37 a_544_297# B1 1.13e-19
C38 a_201_297# a_75_199# 0.16f
C39 a_201_297# B1 0.00594f
C40 a_75_199# C1 0.0628f
C41 B1 C1 0.066f
C42 a_75_199# A3 0.163f
C43 VPWR A1 0.0151f
C44 a_208_47# VPWR 8.35e-19
C45 a_75_199# B1 0.102f
C46 VGND A1 0.0113f
C47 a_208_47# VGND 0.00302f
C48 X A1 1.2e-19
C49 VPWR VGND 0.0735f
C50 A2 A1 0.0689f
C51 a_208_47# X 1.91e-19
C52 a_208_47# A2 0.00102f
C53 X VPWR 0.0676f
C54 VPWR A2 0.0174f
C55 VPB A1 0.0306f
C56 a_315_47# A1 0.00313f
C57 X VGND 0.0609f
C58 VPB VPWR 0.0749f
C59 a_201_297# A1 0.011f
C60 VGND A2 0.0119f
C61 a_315_47# VPWR 0.00154f
C62 a_544_297# VPWR 0.0105f
C63 X A2 3.01e-19
C64 C1 A1 3.21e-19
C65 a_201_297# VPWR 0.211f
C66 VPB VGND 0.00772f
C67 VGND VNB 0.437f
C68 VPWR VNB 0.365f
C69 X VNB 0.0906f
C70 C1 VNB 0.148f
C71 B1 VNB 0.0947f
C72 A1 VNB 0.101f
C73 A2 VNB 0.11f
C74 A3 VNB 0.0908f
C75 VPB VNB 0.782f
C76 a_201_297# VNB 0.00345f
C77 a_75_199# VNB 0.205f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_181_47# a_109_47# a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
C0 A VPWR 0.0185f
C1 B C 0.0746f
C2 VGND VPWR 0.0475f
C3 A VPB 0.0426f
C4 VGND X 0.0708f
C5 A a_27_47# 0.157f
C6 VGND VPB 0.00604f
C7 VGND a_27_47# 0.134f
C8 VPWR C 0.00464f
C9 X C 0.0149f
C10 VPB C 0.0347f
C11 C a_27_47# 0.186f
C12 a_181_47# VPWR 3.97e-19
C13 VGND A 0.0154f
C14 a_181_47# a_27_47# 0.00401f
C15 VGND C 0.0703f
C16 VGND a_181_47# 0.00261f
C17 a_181_47# C 0.00151f
C18 VPWR a_109_47# 3.29e-19
C19 B VPWR 0.128f
C20 a_27_47# a_109_47# 0.00517f
C21 X B 0.00111f
C22 VPB B 0.0836f
C23 B a_27_47# 0.0625f
C24 A a_109_47# 6.45e-19
C25 X VPWR 0.0766f
C26 VPB VPWR 0.0795f
C27 VGND a_109_47# 0.00123f
C28 VPWR a_27_47# 0.145f
C29 X VPB 0.0121f
C30 A B 0.0869f
C31 X a_27_47# 0.087f
C32 VPB a_27_47# 0.0501f
C33 VGND B 0.00714f
C34 VGND VNB 0.3f
C35 X VNB 0.0923f
C36 C VNB 0.12f
C37 A VNB 0.174f
C38 VPWR VNB 0.274f
C39 B VNB 0.102f
C40 VPB VNB 0.516f
C41 a_27_47# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
C0 VPWR VPB 0.0625f
C1 VPWR VGND 0.353f
C2 VPB VGND 0.0797f
C3 VPWR VNB 0.47f
C4 VGND VNB 0.427f
C5 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VPWR VPB 0.0787f
C1 VPWR VGND 0.546f
C2 VPB VGND 0.116f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_384_47# a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
C0 a_299_297# a_81_21# 0.0821f
C1 A1 a_384_47# 0.00884f
C2 B1 a_81_21# 0.148f
C3 VPWR a_384_47# 4.08e-19
C4 VPB a_81_21# 0.0593f
C5 a_299_297# A2 0.0468f
C6 X VGND 0.0512f
C7 VPB A2 0.0373f
C8 a_81_21# a_384_47# 0.00138f
C9 X VPWR 0.0847f
C10 B1 a_299_297# 0.00863f
C11 X a_81_21# 0.112f
C12 VPB a_299_297# 0.0111f
C13 VPB B1 0.0387f
C14 a_299_297# a_384_47# 1.48e-19
C15 B1 X 3.04e-20
C16 VPB X 0.0108f
C17 A1 VGND 0.0786f
C18 VPWR VGND 0.0579f
C19 A1 VPWR 0.0209f
C20 a_81_21# VGND 0.173f
C21 A1 a_81_21# 0.0568f
C22 A2 VGND 0.0495f
C23 VPWR a_81_21# 0.146f
C24 A1 A2 0.0921f
C25 A2 VPWR 0.0201f
C26 a_299_297# VGND 0.00772f
C27 B1 VGND 0.0181f
C28 A2 a_81_21# 7.47e-19
C29 A1 a_299_297# 0.0585f
C30 VPB VGND 0.00713f
C31 B1 A1 0.0817f
C32 a_299_297# VPWR 0.202f
C33 B1 VPWR 0.0196f
C34 VPB A1 0.0264f
C35 VPB VPWR 0.068f
C36 a_384_47# VGND 0.00366f
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_pr__nfet_01v8_D7Y3TR a_n63_n101# a_n33_n75# a_n249_n145# a_63_n75#
+ a_n125_n75#
X0 a_63_n75# a_n63_n101# a_n33_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.233 pd=2.12 as=0.124 ps=1.08 w=0.75 l=0.15
X1 a_n33_n75# a_n63_n101# a_n125_n75# a_n249_n145# sky130_fd_pr__nfet_01v8 ad=0.124 pd=1.08 as=0.233 ps=2.12 w=0.75 l=0.15
C0 a_n63_n101# a_n33_n75# 0.0186f
C1 a_n33_n75# a_63_n75# 0.113f
C2 a_n33_n75# a_n125_n75# 0.113f
C3 a_n63_n101# a_63_n75# 0.0104f
C4 a_n63_n101# a_n125_n75# 0.00451f
C5 a_63_n75# a_n249_n145# 0.0963f
C6 a_n33_n75# a_n249_n145# 0.0361f
C7 a_n125_n75# a_n249_n145# 0.105f
C8 a_n63_n101# a_n249_n145# 0.294f
.ends

.subckt sky130_fd_pr__pfet_01v8_2ZD99F w_n349_n261# a_n153_n139# a_n211_n42# a_153_n42#
+ VSUBS
X0 a_153_n42# a_n153_n139# a_n211_n42# w_n349_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.53
C0 w_n349_n261# a_n211_n42# 0.034f
C1 a_n211_n42# a_153_n42# 0.0169f
C2 a_n211_n42# a_n153_n139# 0.0177f
C3 w_n349_n261# a_153_n42# 0.0179f
C4 w_n349_n261# a_n153_n139# 0.388f
C5 a_n153_n139# a_153_n42# 0.0177f
C6 a_153_n42# VSUBS 0.0558f
C7 a_n211_n42# VSUBS 0.0456f
C8 a_n153_n139# VSUBS 0.556f
C9 w_n349_n261# VSUBS 1.16f
.ends

.subckt sky130_fd_pr__nfet_01v8_2BW22M a_154_n42# a_n154_n130# a_n314_n182# a_n212_n42#
X0 a_154_n42# a_n154_n130# a_n212_n42# a_n314_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.54
C0 a_n154_n130# a_154_n42# 0.0178f
C1 a_154_n42# a_n212_n42# 0.0169f
C2 a_n154_n130# a_n212_n42# 0.0178f
C3 a_154_n42# a_n314_n182# 0.0737f
C4 a_n212_n42# a_n314_n182# 0.0816f
C5 a_n154_n130# a_n314_n182# 0.924f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJP3BL a_15_n150# w_n211_n369# a_n73_n150# a_n33_n247#
+ VSUBS
X0 a_15_n150# a_n33_n247# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.15
C0 w_n211_n369# a_n73_n150# 0.0292f
C1 a_n73_n150# a_15_n150# 0.242f
C2 a_n73_n150# a_n33_n247# 0.0267f
C3 w_n211_n369# a_15_n150# 0.0292f
C4 w_n211_n369# a_n33_n247# 0.19f
C5 a_n33_n247# a_15_n150# 0.0267f
C6 a_15_n150# VSUBS 0.126f
C7 a_n73_n150# VSUBS 0.126f
C8 a_n33_n247# VSUBS 0.146f
C9 w_n211_n369# VSUBS 1.02f
.ends

.subckt sky130_fd_pr__nfet_01v8_LH5FDA a_n150_n130# a_276_n182# a_n208_n42# a_150_n42#
X0 a_150_n42# a_n150_n130# a_n208_n42# a_276_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.5
C0 a_n150_n130# a_150_n42# 0.0176f
C1 a_150_n42# a_n208_n42# 0.0172f
C2 a_n150_n130# a_n208_n42# 0.0176f
C3 a_150_n42# a_276_n182# 0.0815f
C4 a_n208_n42# a_276_n182# 0.0736f
C5 a_n150_n130# a_276_n182# 0.904f
.ends

.subckt th02 Vin V02 m1_983_133# Vp m1_571_144# Vn
XXM0 Vin Vn Vn m1_983_133# m1_983_133# sky130_fd_pr__nfet_01v8_D7Y3TR
XXM1 Vp Vin m1_571_144# m1_983_133# Vn sky130_fd_pr__pfet_01v8_2ZD99F
XXM2 m1_571_144# Vp Vn Vp sky130_fd_pr__nfet_01v8_2BW22M
XXM3 V02 Vp Vp m1_983_133# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_983_133# Vn V02 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 m1_983_133# Vin 0.279f
C1 m1_983_133# m1_571_144# 0.0183f
C2 m1_983_133# V02 0.155f
C3 m1_983_133# Vn 0.216f
C4 Vin m1_571_144# 0.332f
C5 m1_983_133# Vp 0.366f
C6 Vin V02 0.00845f
C7 V02 m1_571_144# 0.011f
C8 Vin Vn 0.0263f
C9 Vn m1_571_144# 0.00115f
C10 V02 Vn 0.00239f
C11 Vin Vp 0.25f
C12 m1_571_144# Vp 0.176f
C13 V02 Vp 0.118f
C14 Vn Vp 0.0235f
C15 Vn 0 0.263f
C16 V02 0 0.334f
C17 m1_983_133# 0 1.44f
C18 Vp 0 3.16f
C19 m1_571_144# 0 0.252f
C20 Vin 0 0.949f
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 VPB VPWR 0.0521f
C1 VGND Y 0.155f
C2 VGND VPB 0.00649f
C3 Y A 0.0894f
C4 VPB A 0.0742f
C5 VGND VPWR 0.0423f
C6 Y VPB 0.0061f
C7 A VPWR 0.0631f
C8 VGND A 0.0638f
C9 Y VPWR 0.209f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X a_29_53# a_183_297# a_111_297#
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 A VPB 0.0377f
C1 VPWR VPB 0.0649f
C2 B A 0.0787f
C3 A a_111_297# 0.00223f
C4 B VPWR 0.147f
C5 VPWR a_111_297# 5.94e-19
C6 VGND a_183_297# 5.75e-19
C7 A a_29_53# 0.242f
C8 VPWR a_29_53# 0.0833f
C9 VGND C 0.0161f
C10 VGND X 0.036f
C11 C VPB 0.0396f
C12 B C 0.0802f
C13 VGND VPB 0.00724f
C14 a_29_53# a_183_297# 0.00868f
C15 VPB X 0.0109f
C16 VGND B 0.0152f
C17 VPWR A 0.00936f
C18 B X 6.52e-19
C19 VGND a_111_297# 3.96e-19
C20 C a_29_53# 0.0857f
C21 B VPB 0.0962f
C22 VGND a_29_53# 0.217f
C23 a_29_53# X 0.0991f
C24 A a_183_297# 0.00239f
C25 VPB a_29_53# 0.0491f
C26 VPWR a_183_297# 8.13e-19
C27 B a_29_53# 0.121f
C28 a_111_297# a_29_53# 0.005f
C29 C A 0.0343f
C30 VPWR C 0.00457f
C31 VGND A 0.0187f
C32 A X 0.00127f
C33 VGND VPWR 0.0459f
C34 VPWR X 0.0885f
C35 VGND VNB 0.306f
C36 X VNB 0.0882f
C37 A VNB 0.117f
C38 C VNB 0.16f
C39 B VNB 0.117f
C40 VPWR VNB 0.253f
C41 VPB VNB 0.516f
C42 a_29_53# VNB 0.18f
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
C0 VGND VPB 0.161f
C1 VGND VPWR 0.903f
C2 VPWR VPB 0.0858f
C3 VPWR VNB 0.867f
C4 VGND VNB 0.761f
C5 VPB VNB 0.605f
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 Y B 0.0877f
C1 VPB VPWR 0.0449f
C2 VPWR A 0.0528f
C3 Y a_109_297# 0.0113f
C4 VGND Y 0.154f
C5 VGND B 0.0451f
C6 VPB A 0.0415f
C7 Y VPWR 0.0995f
C8 B VPWR 0.0148f
C9 VGND a_109_297# 0.00128f
C10 VPB Y 0.0139f
C11 Y A 0.0471f
C12 a_109_297# VPWR 0.00638f
C13 VGND VPWR 0.0314f
C14 VPB B 0.0367f
C15 B A 0.0584f
C16 VGND VPB 0.00456f
C17 VGND A 0.0486f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X a_193_297# a_465_47#
+ a_205_47# a_109_297# a_27_47#
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
C0 VPB a_109_297# 0.00421f
C1 a_27_47# VGND 0.395f
C2 a_109_297# A1 1.05e-19
C3 a_465_47# A1 7.06e-19
C4 a_193_297# VPB 0.00774f
C5 a_109_297# X 3.99e-19
C6 a_193_297# A1 0.0109f
C7 a_465_47# X 1.56e-19
C8 A2 a_27_47# 0.153f
C9 VPB B2 0.0256f
C10 B1 VGND 0.0133f
C11 a_27_47# C1 0.0792f
C12 a_193_297# X 0.00367f
C13 VPWR VGND 0.0722f
C14 X B2 6.77e-20
C15 A2 VPWR 0.0209f
C16 B1 C1 6.46e-19
C17 a_193_297# a_109_297# 0.0927f
C18 C1 VPWR 0.0139f
C19 a_109_297# B2 0.0133f
C20 VPB a_27_47# 0.0512f
C21 a_27_47# A1 0.0984f
C22 a_193_297# B2 0.00126f
C23 a_27_47# X 0.0921f
C24 VPB B1 0.0321f
C25 B1 A1 0.0609f
C26 VPB VPWR 0.0799f
C27 VPWR A1 0.0161f
C28 A2 VGND 0.0168f
C29 B1 X 9.58e-20
C30 a_27_47# a_109_297# 0.0961f
C31 a_465_47# a_27_47# 0.013f
C32 VPWR X 0.0897f
C33 C1 VGND 0.0196f
C34 a_193_297# a_27_47# 0.144f
C35 a_27_47# B2 0.0959f
C36 B1 a_109_297# 0.00736f
C37 A2 C1 9.03e-21
C38 a_109_297# VPWR 0.15f
C39 a_465_47# VPWR 5.05e-19
C40 a_193_297# B1 0.00869f
C41 a_193_297# VPWR 0.169f
C42 VPB VGND 0.00844f
C43 B1 B2 0.0784f
C44 a_27_47# a_205_47# 0.00762f
C45 A1 VGND 0.0126f
C46 VPWR B2 0.00842f
C47 X VGND 0.061f
C48 A2 VPB 0.027f
C49 A2 A1 0.0692f
C50 VPB C1 0.0367f
C51 C1 A1 1.77e-20
C52 a_205_47# VPWR 1.62e-19
C53 A2 X 0.00157f
C54 a_109_297# VGND 0.00284f
C55 C1 X 5.03e-20
C56 a_465_47# VGND 0.00257f
C57 a_27_47# B1 0.112f
C58 a_27_47# VPWR 0.099f
C59 a_193_297# VGND 0.00438f
C60 VGND B2 0.0174f
C61 C1 a_109_297# 0.00739f
C62 VPB A1 0.0343f
C63 A2 a_193_297# 0.00683f
C64 B1 VPWR 0.00982f
C65 VPB X 0.0113f
C66 X A1 2.77e-19
C67 a_205_47# VGND 0.00156f
C68 C1 B2 0.0726f
C69 VGND VNB 0.437f
C70 X VNB 0.0919f
C71 VPWR VNB 0.364f
C72 A2 VNB 0.0896f
C73 A1 VNB 0.106f
C74 B1 VNB 0.108f
C75 B2 VNB 0.0887f
C76 C1 VNB 0.139f
C77 VPB VNB 0.782f
C78 a_193_297# VNB 0.0011f
C79 a_109_297# VNB 7.11e-19
C80 a_27_47# VNB 0.216f
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X a_256_47# a_584_47#
+ a_93_21# a_250_297# a_346_47#
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
C0 a_250_297# A3 0.00602f
C1 A2 B1 1.44e-20
C2 A2 a_256_47# 0.00256f
C3 VGND B1 0.0344f
C4 B1 a_93_21# 0.0774f
C5 B1 VPWR 0.01f
C6 a_250_297# VPB 0.00616f
C7 VGND a_256_47# 0.00394f
C8 a_256_47# a_93_21# 0.0114f
C9 VPWR a_256_47# 9.47e-19
C10 a_250_297# A1 0.0129f
C11 a_250_297# X 5.42e-19
C12 a_250_297# B2 0.0344f
C13 A3 VPB 0.0291f
C14 A2 VGND 0.0114f
C15 A2 a_93_21# 0.0747f
C16 A3 X 2.45e-19
C17 A2 VPWR 0.0133f
C18 B2 A3 9.12e-20
C19 VGND a_93_21# 0.251f
C20 VGND VPWR 0.076f
C21 B1 a_250_297# 0.0125f
C22 VPWR a_93_21# 0.0907f
C23 B1 a_584_47# 0.00143f
C24 VPB A1 0.0296f
C25 X VPB 0.0108f
C26 B2 VPB 0.0355f
C27 B1 A3 7.88e-22
C28 X A1 6.03e-20
C29 a_346_47# A1 0.00465f
C30 A3 a_256_47# 4.42e-19
C31 B2 A1 3.14e-19
C32 A2 a_250_297# 0.0129f
C33 B1 VPB 0.0276f
C34 VGND a_250_297# 0.0072f
C35 a_250_297# a_93_21# 0.188f
C36 a_250_297# VPWR 0.313f
C37 VGND a_584_47# 0.00683f
C38 a_584_47# a_93_21# 0.00278f
C39 a_584_47# VPWR 9.47e-19
C40 A2 A3 0.0788f
C41 B1 A1 0.0965f
C42 B1 X 3.83e-20
C43 a_346_47# B1 5.39e-20
C44 B1 B2 0.0823f
C45 VGND A3 0.00974f
C46 A3 a_93_21# 0.124f
C47 A3 VPWR 0.0158f
C48 A2 VPB 0.0287f
C49 A2 A1 0.0971f
C50 VGND VPB 0.00788f
C51 A2 X 1.19e-19
C52 VPB a_93_21# 0.0485f
C53 a_346_47# A2 0.00252f
C54 VPWR VPB 0.0756f
C55 B1 a_256_47# 2.07e-20
C56 A2 B2 1.46e-19
C57 a_250_297# a_584_47# 2.43e-19
C58 VGND A1 0.0133f
C59 VGND X 0.06f
C60 A1 a_93_21# 0.0641f
C61 a_346_47# VGND 0.00514f
C62 X a_93_21# 0.0841f
C63 VPWR A1 0.016f
C64 X VPWR 0.0849f
C65 a_346_47# a_93_21# 0.0119f
C66 a_346_47# VPWR 0.00109f
C67 VGND B2 0.0469f
C68 B2 a_93_21# 0.0147f
C69 B2 VPWR 0.0108f
C70 VGND VNB 0.465f
C71 VPWR VNB 0.365f
C72 X VNB 0.0937f
C73 B2 VNB 0.14f
C74 B1 VNB 0.101f
C75 A1 VNB 0.0951f
C76 A2 VNB 0.0921f
C77 A3 VNB 0.0929f
C78 VPB VNB 0.782f
C79 a_250_297# VNB 0.0278f
C80 a_93_21# VNB 0.151f
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X a_277_297# a_205_297# a_27_297#
+ a_109_297#
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 VGND A 0.016f
C1 a_27_297# a_205_297# 0.00412f
C2 a_277_297# B 2.29e-19
C3 VGND a_109_297# 7.58e-19
C4 VPWR a_205_297# 5.16e-19
C5 a_27_297# C 0.158f
C6 VGND a_277_297# 4.65e-19
C7 D A 2.13e-19
C8 VPWR C 0.00723f
C9 C VPB 0.0338f
C10 X A 0.00133f
C11 B C 0.0917f
C12 a_27_297# VPWR 0.084f
C13 a_205_297# VGND 3.36e-19
C14 a_27_297# VPB 0.0517f
C15 a_277_297# X 6.43e-20
C16 VGND C 0.0191f
C17 VPWR VPB 0.075f
C18 a_27_297# B 0.159f
C19 VPWR B 0.193f
C20 a_27_297# VGND 0.235f
C21 D C 0.0954f
C22 a_277_297# A 2.28e-19
C23 B VPB 0.106f
C24 VPWR VGND 0.0546f
C25 VGND VPB 0.00796f
C26 a_27_297# D 0.054f
C27 VGND B 0.0159f
C28 VPWR D 0.00503f
C29 D VPB 0.0405f
C30 a_27_297# X 0.0991f
C31 C A 0.028f
C32 VPWR X 0.0878f
C33 B D 0.00287f
C34 C a_109_297# 0.00356f
C35 X VPB 0.0109f
C36 a_277_297# C 5.54e-19
C37 a_27_297# A 0.163f
C38 VGND D 0.0517f
C39 B X 6.42e-19
C40 a_27_297# a_109_297# 0.00695f
C41 VPWR A 0.00769f
C42 VPB A 0.033f
C43 a_27_297# a_277_297# 0.00876f
C44 VGND X 0.0354f
C45 VPWR a_109_297# 9.23e-19
C46 a_205_297# C 0.00261f
C47 VPWR a_277_297# 7.48e-19
C48 B A 0.0639f
C49 VGND VNB 0.367f
C50 X VNB 0.0883f
C51 A VNB 0.109f
C52 C VNB 0.105f
C53 D VNB 0.175f
C54 B VNB 0.115f
C55 VPWR VNB 0.29f
C56 VPB VNB 0.605f
C57 a_27_297# VNB 0.163f
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
C0 VPWR VGND 1.57f
C1 VPWR VPB 0.137f
C2 VPB VGND 0.35f
C3 VPWR VNB 1.67f
C4 VGND VNB 1.47f
C5 VPB VNB 1.14f
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X a_369_47# a_469_47#
+ a_297_47# a_193_413# a_27_47#
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VGND a_369_47# 0.00505f
C1 VPWR B 0.0186f
C2 A_N VPWR 0.02f
C3 VGND a_297_47# 0.00183f
C4 VPB a_193_413# 0.0644f
C5 D a_193_413# 0.155f
C6 a_193_413# X 0.108f
C7 VGND B 0.037f
C8 a_193_413# C 0.0389f
C9 A_N VGND 0.0205f
C10 B a_27_47# 0.0794f
C11 A_N a_27_47# 0.237f
C12 VPWR a_193_413# 0.281f
C13 a_369_47# B 0.00129f
C14 VPB D 0.0763f
C15 VPB X 0.0108f
C16 VPB C 0.0742f
C17 a_469_47# a_193_413# 0.00109f
C18 D X 0.0168f
C19 D C 0.183f
C20 C X 0.00479f
C21 VPB VPWR 0.0818f
C22 B a_297_47# 0.00353f
C23 VGND a_193_413# 0.0915f
C24 D VPWR 0.0186f
C25 VPWR X 0.0586f
C26 a_27_47# a_193_413# 0.125f
C27 VPWR C 0.0182f
C28 D a_469_47# 0.00183f
C29 a_469_47# X 0.001f
C30 a_469_47# C 0.00202f
C31 a_369_47# a_193_413# 0.00181f
C32 VPB VGND 0.0123f
C33 VPB a_27_47# 0.092f
C34 D VGND 0.0372f
C35 a_469_47# VPWR 7.77e-19
C36 VGND X 0.0588f
C37 VGND C 0.0395f
C38 a_193_413# a_297_47# 0.00137f
C39 VGND VPWR 0.0727f
C40 VPWR a_27_47# 0.106f
C41 a_369_47# C 0.00448f
C42 B a_193_413# 0.144f
C43 A_N a_193_413# 0.00151f
C44 a_469_47# VGND 0.00551f
C45 VPWR a_369_47# 6.65e-19
C46 VPB B 0.089f
C47 A_N VPB 0.0832f
C48 VGND a_27_47# 0.103f
C49 B C 0.164f
C50 VPWR a_297_47# 2.82e-19
C51 VGND VNB 0.456f
C52 X VNB 0.0934f
C53 VPWR VNB 0.368f
C54 D VNB 0.123f
C55 C VNB 0.108f
C56 B VNB 0.12f
C57 A_N VNB 0.198f
C58 VPB VNB 0.782f
C59 a_193_413# VNB 0.136f
C60 a_27_47# VNB 0.224f
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X a_109_93# a_368_53# a_209_311#
+ a_296_53#
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
C0 VGND a_368_53# 0.0031f
C1 C A_N 7.6e-19
C2 VPWR a_368_53# 4.26e-19
C3 X A_N 1.44e-19
C4 B a_109_93# 0.0802f
C5 VGND B 0.00796f
C6 B VPWR 0.131f
C7 a_209_311# A_N 0.00515f
C8 VPB a_109_93# 0.0652f
C9 VGND VPB 0.00909f
C10 VPB VPWR 0.104f
C11 X C 0.0176f
C12 C a_209_311# 0.19f
C13 B A_N 2.03e-19
C14 X a_209_311# 0.0877f
C15 a_296_53# a_209_311# 0.0049f
C16 C a_368_53# 0.00415f
C17 VPB A_N 0.111f
C18 B C 0.0671f
C19 a_368_53# a_209_311# 0.0026f
C20 X B 0.00119f
C21 VGND a_109_93# 0.0784f
C22 VPWR a_109_93# 0.0984f
C23 VPB C 0.0339f
C24 VGND VPWR 0.0657f
C25 B a_209_311# 0.0609f
C26 X VPB 0.0119f
C27 VPB a_209_311# 0.0515f
C28 a_109_93# A_N 0.117f
C29 VGND A_N 0.045f
C30 VPWR A_N 0.0513f
C31 B VPB 0.0914f
C32 C a_109_93# 3.91e-20
C33 VGND C 0.0678f
C34 VPWR C 0.005f
C35 VGND X 0.0647f
C36 a_296_53# a_109_93# 1.84e-19
C37 X VPWR 0.0732f
C38 VGND a_296_53# 6.07e-19
C39 a_109_93# a_209_311# 0.168f
C40 VGND a_209_311# 0.131f
C41 a_296_53# VPWR 1.15e-19
C42 VPWR a_209_311# 0.155f
C43 VGND VNB 0.44f
C44 X VNB 0.0925f
C45 C VNB 0.114f
C46 B VNB 0.101f
C47 VPWR VNB 0.342f
C48 A_N VNB 0.197f
C49 VPB VNB 0.693f
C50 a_209_311# VNB 0.143f
C51 a_109_93# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
C0 VPWR VGND 0.057f
C1 VPB VGND 0.00583f
C2 a_27_47# X 0.328f
C3 A a_27_47# 0.195f
C4 VPB VPWR 0.0632f
C5 VGND a_27_47# 0.148f
C6 VPWR a_27_47# 0.219f
C7 VPB a_27_47# 0.139f
C8 A X 0.014f
C9 VGND X 0.216f
C10 A VGND 0.0431f
C11 VPWR X 0.317f
C12 A VPWR 0.022f
C13 VPB X 0.0122f
C14 A VPB 0.0321f
C15 VGND VNB 0.358f
C16 X VNB 0.067f
C17 VPWR VNB 0.308f
C18 A VNB 0.148f
C19 VPB VNB 0.605f
C20 a_27_47# VNB 0.543f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
C0 VPWR B 0.0117f
C1 a_59_75# A 0.0809f
C2 VPB a_59_75# 0.0563f
C3 B VGND 0.0115f
C4 VPWR a_145_75# 6.31e-19
C5 a_145_75# VGND 0.00468f
C6 B a_59_75# 0.143f
C7 X A 1.68e-19
C8 VPWR VGND 0.0461f
C9 VPB X 0.0127f
C10 a_59_75# a_145_75# 0.00658f
C11 VPWR a_59_75# 0.15f
C12 B X 0.00276f
C13 VPB A 0.0806f
C14 a_59_75# VGND 0.116f
C15 a_145_75# X 5.76e-19
C16 VPWR X 0.111f
C17 B A 0.0971f
C18 VPB B 0.0629f
C19 X VGND 0.0993f
C20 VPWR A 0.0362f
C21 VPB VPWR 0.0729f
C22 a_59_75# X 0.109f
C23 A VGND 0.0147f
C24 VPB VGND 0.008f
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y a_297_297# a_191_297#
+ a_109_297#
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_191_297# VGND 9.29e-19
C1 VGND VPB 0.0048f
C2 B Y 0.0403f
C3 A VPWR 0.0483f
C4 A a_297_297# 3.16e-19
C5 VPWR a_109_297# 0.00576f
C6 a_191_297# C 0.0195f
C7 VPB C 0.0299f
C8 a_191_297# Y 0.00142f
C9 VPB Y 0.0127f
C10 VPWR B 0.0887f
C11 B a_297_297# 0.0132f
C12 VGND C 0.0184f
C13 VGND Y 0.151f
C14 VPWR a_191_297# 0.0049f
C15 A B 0.11f
C16 VPWR VPB 0.0524f
C17 C Y 0.125f
C18 VPB D 0.0376f
C19 VPWR VGND 0.0492f
C20 VGND a_297_297# 8.1e-19
C21 VGND D 0.0456f
C22 A VPB 0.041f
C23 VPWR C 0.0509f
C24 A VGND 0.0526f
C25 VPWR Y 0.0561f
C26 D C 0.0523f
C27 a_297_297# Y 1.24e-19
C28 a_191_297# B 0.00223f
C29 VGND a_109_297# 0.00181f
C30 D Y 0.108f
C31 B VPB 0.0304f
C32 A C 0.00268f
C33 B VGND 0.0191f
C34 A Y 0.0175f
C35 C a_109_297# 0.0062f
C36 VPWR a_297_297# 0.00317f
C37 Y a_109_297# 0.0122f
C38 VPWR D 0.0128f
C39 B C 0.173f
C40 VGND VNB 0.322f
C41 VPWR VNB 0.276f
C42 Y VNB 0.0645f
C43 A VNB 0.174f
C44 B VNB 0.0968f
C45 C VNB 0.0911f
C46 D VNB 0.159f
C47 VPB VNB 0.516f
.ends

.subckt sky130_fd_pr__nfet_01v8_2V6S9N a_n216_n42# a_158_n42# a_n158_n130# a_n284_n216#
X0 a_158_n42# a_n158_n130# a_n216_n42# a_n284_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.58
C0 a_158_n42# a_n158_n130# 0.018f
C1 a_n216_n42# a_158_n42# 0.0165f
C2 a_n216_n42# a_n158_n130# 0.018f
C3 a_158_n42# a_n284_n216# 0.0746f
C4 a_n216_n42# a_n284_n216# 0.0746f
C5 a_n158_n130# a_n284_n216# 0.981f
.ends

.subckt sky130_fd_pr__pfet_01v8_XYZSMQ a_n33_n255# a_15_n158# w_n211_n377# a_n73_n158#
+ VSUBS
X0 a_15_n158# a_n33_n255# a_n73_n158# w_n211_n377# sky130_fd_pr__pfet_01v8 ad=0.458 pd=3.74 as=0.458 ps=3.74 w=1.58 l=0.15
C0 a_n73_n158# w_n211_n377# 0.0299f
C1 a_n73_n158# a_15_n158# 0.254f
C2 a_n33_n255# a_n73_n158# 0.0271f
C3 a_15_n158# w_n211_n377# 0.0299f
C4 a_n33_n255# w_n211_n377# 0.191f
C5 a_n33_n255# a_15_n158# 0.0271f
C6 a_15_n158# VSUBS 0.132f
C7 a_n73_n158# VSUBS 0.132f
C8 a_n33_n255# VSUBS 0.146f
C9 w_n211_n377# VSUBS 1.04f
.ends

.subckt sky130_fd_pr__pfet_01v8_AZD9DW w_n353_n261# a_n157_n139# a_n215_n42# a_157_n42#
+ VSUBS
X0 a_157_n42# a_n157_n139# a_n215_n42# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.57
C0 a_n215_n42# w_n353_n261# 0.0179f
C1 a_n215_n42# a_157_n42# 0.0166f
C2 a_n157_n139# a_n215_n42# 0.0179f
C3 a_157_n42# w_n353_n261# 0.0323f
C4 a_n157_n139# w_n353_n261# 0.396f
C5 a_n157_n139# a_157_n42# 0.0179f
C6 a_157_n42# VSUBS 0.0468f
C7 a_n215_n42# VSUBS 0.0559f
C8 a_n157_n139# VSUBS 0.569f
C9 w_n353_n261# VSUBS 1.17f
.ends

.subckt sky130_fd_pr__nfet_01v8_T8HSQ7 a_n175_n297# a_15_n157# a_n33_n245# a_n73_n157#
X0 a_15_n157# a_n33_n245# a_n73_n157# a_n175_n297# sky130_fd_pr__nfet_01v8 ad=0.455 pd=3.72 as=0.455 ps=3.72 w=1.57 l=0.15
C0 a_15_n157# a_n33_n245# 0.0289f
C1 a_n73_n157# a_15_n157# 0.253f
C2 a_n73_n157# a_n33_n245# 0.0289f
C3 a_15_n157# a_n175_n297# 0.161f
C4 a_n73_n157# a_n175_n297# 0.188f
C5 a_n33_n245# a_n175_n297# 0.322f
.ends

.subckt th09 V09 Vin Vn m1_485_n505# Vp m1_962_372#
XXM0 m1_485_n505# Vn Vin Vn sky130_fd_pr__nfet_01v8_2V6S9N
XXM1 Vin m1_485_n505# Vp Vp Vn sky130_fd_pr__pfet_01v8_XYZSMQ
XXM2 Vp m1_485_n505# Vp m1_962_372# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM3 Vp m1_485_n505# V09 m1_962_372# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM4 Vn V09 m1_485_n505# Vn sky130_fd_pr__nfet_01v8_T8HSQ7
C0 Vp Vin 0.187f
C1 m1_485_n505# V09 0.104f
C2 Vin m1_962_372# 0.00821f
C3 Vn Vp 0.0176f
C4 Vn m1_962_372# 6.71e-21
C5 Vin V09 2.77e-19
C6 Vn V09 0.00364f
C7 m1_485_n505# Vin 0.372f
C8 Vn m1_485_n505# 0.0846f
C9 Vp m1_962_372# 0.0579f
C10 Vp V09 0.0743f
C11 Vn Vin 0.0386f
C12 V09 m1_962_372# 0.00205f
C13 Vp m1_485_n505# 0.372f
C14 m1_485_n505# m1_962_372# 0.0822f
C15 Vin 0 1.1f
C16 m1_485_n505# 0 1.18f
C17 V09 0 0.27f
C18 Vn 0 0.344f
C19 m1_962_372# 0 0.118f
C20 Vp 0 3.27f
.ends

.subckt sky130_fd_pr__pfet_01v8_HPNF99 a_n33_n147# a_23_n50# a_n81_n50# w_n219_n269#
+ VSUBS
X0 a_23_n50# a_n33_n147# a_n81_n50# w_n219_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.23
C0 a_n81_n50# a_23_n50# 0.07f
C1 w_n219_n269# a_n33_n147# 0.173f
C2 a_n81_n50# w_n219_n269# 0.0419f
C3 a_23_n50# w_n219_n269# 0.0185f
C4 a_n81_n50# a_n33_n147# 0.00814f
C5 a_23_n50# a_n33_n147# 0.00814f
C6 a_23_n50# VSUBS 0.0578f
C7 a_n81_n50# VSUBS 0.0428f
C8 a_n33_n147# VSUBS 0.157f
C9 w_n219_n269# VSUBS 0.779f
.ends

.subckt sky130_fd_pr__nfet_01v8_JZU22M a_n213_n42# a_155_n42# a_n155_n130# a_281_n238#
X0 a_155_n42# a_n155_n130# a_n213_n42# a_281_n238# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.55
C0 a_n155_n130# a_n213_n42# 0.0178f
C1 a_155_n42# a_n155_n130# 0.0178f
C2 a_155_n42# a_n213_n42# 0.0168f
C3 a_155_n42# a_281_n238# 0.0816f
C4 a_n213_n42# a_281_n238# 0.0737f
C5 a_n155_n130# a_281_n238# 0.928f
.ends

.subckt sky130_fd_pr__pfet_01v8_TM5S5A a_n80_n147# a_n138_n50# a_80_n50# w_n276_n269#
+ VSUBS
X0 a_80_n50# a_n80_n147# a_n138_n50# w_n276_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.8
C0 a_n138_n50# a_80_n50# 0.0335f
C1 w_n276_n269# a_n80_n147# 0.297f
C2 a_n138_n50# w_n276_n269# 0.0231f
C3 a_80_n50# w_n276_n269# 0.0231f
C4 a_n138_n50# a_n80_n147# 0.0141f
C5 a_80_n50# a_n80_n147# 0.0141f
C6 a_80_n50# VSUBS 0.0565f
C7 a_n138_n50# VSUBS 0.0565f
C8 a_n80_n147# VSUBS 0.296f
C9 w_n276_n269# VSUBS 1.01f
.ends

.subckt sky130_fd_pr__pfet_01v8_AM8GZ5 w_n526_n261# a_n330_n139# a_330_n42# a_n388_n42#
+ VSUBS
X0 a_330_n42# a_n330_n139# a_n388_n42# w_n526_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.3
C0 a_n388_n42# a_330_n42# 0.00853f
C1 w_n526_n261# a_n330_n139# 0.719f
C2 a_n388_n42# w_n526_n261# 0.0179f
C3 a_330_n42# w_n526_n261# 0.0408f
C4 a_n388_n42# a_n330_n139# 0.0223f
C5 a_330_n42# a_n330_n139# 0.0223f
C6 a_330_n42# VSUBS 0.0435f
C7 a_n388_n42# VSUBS 0.0585f
C8 a_n330_n139# VSUBS 1.13f
C9 w_n526_n261# VSUBS 1.76f
.ends

.subckt sky130_fd_pr__nfet_01v8_H7HSAV a_n73_n250# a_15_n250# a_n33_n338# a_n141_n424#
X0 a_15_n250# a_n33_n338# a_n73_n250# a_n141_n424# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.15
C0 a_n33_n338# a_n73_n250# 0.0337f
C1 a_15_n250# a_n33_n338# 0.0337f
C2 a_15_n250# a_n73_n250# 0.401f
C3 a_15_n250# a_n141_n424# 0.24f
C4 a_n73_n250# a_n141_n424# 0.24f
C5 a_n33_n338# a_n141_n424# 0.327f
.ends

.subckt th14 V14 Vin Vn m1_641_n318# Vp m1_891_419#
XXM0 Vn Vn m1_641_n318# Vp Vn sky130_fd_pr__pfet_01v8_HPNF99
XXM1 m1_641_n318# m1_891_419# Vin Vn sky130_fd_pr__nfet_01v8_JZU22M
XXM2 Vin Vp m1_891_419# Vp Vn sky130_fd_pr__pfet_01v8_TM5S5A
XXM3 Vp m1_891_419# V14 Vp Vn sky130_fd_pr__pfet_01v8_AM8GZ5
XXM4 Vn V14 m1_891_419# Vn sky130_fd_pr__nfet_01v8_H7HSAV
C0 Vp Vin 0.201f
C1 Vp V14 0.082f
C2 m1_641_n318# Vp 0.0629f
C3 Vin V14 0.00516f
C4 m1_641_n318# Vin 0.229f
C5 Vp m1_891_419# 0.227f
C6 m1_891_419# Vin 0.132f
C7 m1_891_419# V14 0.249f
C8 m1_641_n318# m1_891_419# 0.00289f
C9 m1_891_419# Vn 1.7f
C10 V14 Vn 0.273f
C11 Vp Vn 3.39f
C12 Vin Vn 1.76f
C13 m1_641_n318# Vn 0.313f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X a_75_212#
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 X VPWR 0.0896f
C1 X a_75_212# 0.107f
C2 VPWR A 0.0217f
C3 VPWR VGND 0.0289f
C4 a_75_212# A 0.178f
C5 VPWR VPB 0.0355f
C6 a_75_212# VGND 0.105f
C7 a_75_212# VPB 0.0571f
C8 X A 8.48e-19
C9 X VGND 0.0545f
C10 X VPB 0.0128f
C11 VGND A 0.0184f
C12 A VPB 0.0525f
C13 VGND VPB 0.00507f
C14 VPWR a_75_212# 0.134f
C15 VGND VNB 0.207f
C16 VPWR VNB 0.176f
C17 X VNB 0.0942f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_75_212# VNB 0.21f
.ends

.subckt sky130_fd_pr__nfet_01v8_VGVEGU a_n142_n216# a_n74_n42# a_n33_n130# a_16_n42#
X0 a_16_n42# a_n33_n130# a_n74_n42# a_n142_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.16
C0 a_n33_n130# a_n74_n42# 0.0191f
C1 a_16_n42# a_n74_n42# 0.0684f
C2 a_n33_n130# a_16_n42# 0.0191f
C3 a_16_n42# a_n142_n216# 0.0652f
C4 a_n74_n42# a_n142_n216# 0.0652f
C5 a_n33_n130# a_n142_n216# 0.317f
.ends

.subckt sky130_fd_pr__pfet_01v8_EDPLE3 a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 w_n211_n261# a_n33_n139# 0.187f
C1 a_15_n42# a_n73_n42# 0.0699f
C2 a_15_n42# a_n33_n139# 0.0192f
C3 a_n73_n42# a_n33_n139# 0.0192f
C4 a_15_n42# w_n211_n261# 0.0197f
C5 w_n211_n261# a_n73_n42# 0.0197f
C6 a_15_n42# VSUBS 0.0445f
C7 a_n73_n42# VSUBS 0.0445f
C8 a_n33_n139# VSUBS 0.143f
C9 w_n211_n261# VSUBS 0.749f
.ends

.subckt sky130_fd_pr__pfet_01v8_JM8GTH a_50_n42# w_n246_n261# a_n50_n139# a_n108_n42#
+ VSUBS
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 w_n246_n261# a_n50_n139# 0.223f
C1 a_50_n42# a_n108_n42# 0.0391f
C2 a_50_n42# a_n50_n139# 0.00909f
C3 a_n108_n42# a_n50_n139# 0.00909f
C4 a_50_n42# w_n246_n261# 0.0224f
C5 w_n246_n261# a_n108_n42# 0.0224f
C6 a_50_n42# VSUBS 0.0488f
C7 a_n108_n42# VSUBS 0.0488f
C8 a_n50_n139# VSUBS 0.209f
C9 w_n246_n261# VSUBS 0.88f
.ends

.subckt sky130_fd_pr__nfet_01v8_MYA4RC a_n73_n46# a_n33_n134# a_15_n46# a_n175_n186#
X0 a_15_n46# a_n33_n134# a_n73_n46# a_n175_n186# sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.5 as=0.133 ps=1.5 w=0.46 l=0.15
C0 a_n33_n134# a_n73_n46# 0.0212f
C1 a_15_n46# a_n73_n46# 0.0763f
C2 a_n33_n134# a_15_n46# 0.0212f
C3 a_15_n46# a_n175_n186# 0.0671f
C4 a_n73_n46# a_n175_n186# 0.0756f
C5 a_n33_n134# a_n175_n186# 0.314f
.ends

.subckt th07 Vp Vin V07 m1_808_n892# Vn
XXM0 Vn m1_808_n892# Vin Vn sky130_fd_pr__nfet_01v8_VGVEGU
XXM1 m1_808_n892# Vp Vin Vp Vn sky130_fd_pr__pfet_01v8_EDPLE3
XXM2 V07 Vp m1_808_n892# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM3 V07 m1_808_n892# Vn Vn sky130_fd_pr__nfet_01v8_MYA4RC
C0 m1_808_n892# Vp 0.209f
C1 Vin V07 0.00135f
C2 V07 Vp 0.0569f
C3 Vin Vp 0.157f
C4 m1_808_n892# V07 0.112f
C5 m1_808_n892# Vin 0.365f
C6 Vin Vn 0.524f
C7 Vp Vn 1.57f
C8 m1_808_n892# Vn 0.596f
C9 V07 Vn 0.276f
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 VPWR A 0.0215f
C1 X VPB 0.0128f
C2 VPWR VGND 0.029f
C3 a_27_47# X 0.107f
C4 VGND A 0.0184f
C5 VPWR VPB 0.0355f
C6 VPWR a_27_47# 0.135f
C7 VPB A 0.0524f
C8 a_27_47# A 0.181f
C9 VGND VPB 0.00505f
C10 a_27_47# VGND 0.105f
C11 a_27_47# VPB 0.0592f
C12 VPWR X 0.0897f
C13 X A 8.48e-19
C14 X VGND 0.0546f
C15 VGND VNB 0.207f
C16 X VNB 0.0941f
C17 VPWR VNB 0.175f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_27_47# VNB 0.208f
.ends

.subckt sky130_fd_pr__pfet_01v8_P28Q2U a_n33_n232# a_15_n135# w_n211_n354# a_n73_n135#
+ VSUBS
X0 a_15_n135# a_n33_n232# a_n73_n135# w_n211_n354# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.28 as=0.391 ps=3.28 w=1.35 l=0.15
C0 a_n33_n232# w_n211_n354# 0.19f
C1 a_15_n135# a_n73_n135# 0.218f
C2 a_15_n135# a_n33_n232# 0.0258f
C3 a_n33_n232# a_n73_n135# 0.0258f
C4 a_15_n135# w_n211_n354# 0.0279f
C5 w_n211_n354# a_n73_n135# 0.0279f
C6 a_15_n135# VSUBS 0.115f
C7 a_n73_n135# VSUBS 0.115f
C8 a_n33_n232# VSUBS 0.146f
C9 w_n211_n354# VSUBS 0.983f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZMY3VB a_n348_n42# a_n290_n130# a_n450_n182# a_290_n42#
X0 a_290_n42# a_n290_n130# a_n348_n42# a_n450_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.9
C0 a_n348_n42# a_n290_n130# 0.0217f
C1 a_n348_n42# a_290_n42# 0.00961f
C2 a_n290_n130# a_290_n42# 0.0217f
C3 a_290_n42# a_n450_n182# 0.076f
C4 a_n348_n42# a_n450_n182# 0.0839f
C5 a_n290_n130# a_n450_n182# 1.6f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n33_n197# w_n211_n319# 0.189f
C1 a_15_n100# a_n73_n100# 0.162f
C2 a_15_n100# a_n33_n197# 0.0236f
C3 a_n33_n197# a_n73_n100# 0.0236f
C4 a_15_n100# w_n211_n319# 0.0248f
C5 w_n211_n319# a_n73_n100# 0.0248f
C6 a_15_n100# VSUBS 0.0885f
C7 a_n73_n100# VSUBS 0.0885f
C8 a_n33_n197# VSUBS 0.145f
C9 w_n211_n319# VSUBS 0.894f
.ends

.subckt sky130_fd_pr__pfet_01v8_WV9GCW a_n158_n42# w_n296_n261# a_n100_n139# a_100_n42#
+ VSUBS
X0 a_100_n42# a_n100_n139# a_n158_n42# w_n296_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1
C0 a_n100_n139# w_n296_n261# 0.346f
C1 a_100_n42# a_n158_n42# 0.024f
C2 a_100_n42# a_n100_n139# 0.0144f
C3 a_n100_n139# a_n158_n42# 0.0144f
C4 a_100_n42# w_n296_n261# 0.0224f
C5 w_n296_n261# a_n158_n42# 0.0224f
C6 a_100_n42# VSUBS 0.0504f
C7 a_n158_n42# VSUBS 0.0504f
C8 a_n100_n139# VSUBS 0.353f
C9 w_n296_n261# VSUBS 1.06f
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n141_240# a_n33_n188# a_15_n100#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n141_240# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n73_n100# a_n33_n188# 0.0254f
C1 a_n73_n100# a_15_n100# 0.162f
C2 a_n33_n188# a_15_n100# 0.0254f
C3 a_15_n100# a_n141_240# 0.113f
C4 a_n73_n100# a_n141_240# 0.113f
C5 a_n33_n188# a_n141_240# 0.322f
.ends

.subckt th12 V12 Vin m1_394_n856# m1_529_n42# Vp Vn
XXM0 Vn Vn Vp m1_394_n856# Vn sky130_fd_pr__pfet_01v8_P28Q2U
XXM1 m1_529_n42# Vin Vn m1_394_n856# sky130_fd_pr__nfet_01v8_ZMY3VB
XXM2 m1_529_n42# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM3 Vp Vp m1_529_n42# V12 Vn sky130_fd_pr__pfet_01v8_WV9GCW
XXM4 V12 Vn m1_529_n42# Vn sky130_fd_pr__nfet_01v8_648S5X
C0 m1_529_n42# m1_394_n856# 0.0134f
C1 m1_529_n42# V12 0.0929f
C2 m1_529_n42# Vp 0.322f
C3 V12 m1_394_n856# 4.74e-19
C4 Vp m1_394_n856# 0.04f
C5 V12 Vp 0.0454f
C6 m1_529_n42# Vin 0.0965f
C7 m1_529_n42# Vn 0.254f
C8 Vin m1_394_n856# 0.321f
C9 V12 Vin 0.00205f
C10 Vn m1_394_n856# 0.0338f
C11 Vp Vin 0.238f
C12 V12 Vn 0.0234f
C13 Vn Vp 0.132f
C14 Vn Vin 0.135f
C15 Vn 0 0.29f
C16 Vp 0 2.88f
C17 m1_529_n42# 0 0.861f
C18 V12 0 0.359f
C19 Vin 0 1.9f
C20 m1_394_n856# 0 0.215f
.ends

.subckt sky130_fd_pr__nfet_01v8_Q7AWK3 a_n180_n340# a_20_n200# a_n78_n200# a_n33_n288#
X0 a_20_n200# a_n33_n288# a_n78_n200# a_n180_n340# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
C0 a_20_n200# a_n78_n200# 0.288f
C1 a_n33_n288# a_20_n200# 0.024f
C2 a_n33_n288# a_n78_n200# 0.024f
C3 a_20_n200# a_n180_n340# 0.202f
C4 a_n78_n200# a_n180_n340# 0.237f
C5 a_n33_n288# a_n180_n340# 0.325f
.ends

.subckt sky130_fd_pr__pfet_01v8_EXJYQP w_n359_n261# a_n163_n139# a_n221_n42# a_163_n42#
+ VSUBS
X0 a_163_n42# a_n163_n139# a_n221_n42# w_n359_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.63
C0 a_n221_n42# a_n163_n139# 0.0182f
C1 a_163_n42# w_n359_n261# 0.0408f
C2 a_163_n42# a_n221_n42# 0.0161f
C3 a_163_n42# a_n163_n139# 0.0182f
C4 w_n359_n261# a_n221_n42# 0.0179f
C5 w_n359_n261# a_n163_n139# 0.413f
C6 a_163_n42# VSUBS 0.041f
C7 a_n221_n42# VSUBS 0.056f
C8 a_n163_n139# VSUBS 0.584f
C9 w_n359_n261# VSUBS 1.24f
.ends

.subckt sky130_fd_pr__pfet_01v8_HJHF6N a_n170_n50# w_n308_n269# a_n112_n147# a_112_n50#
+ VSUBS
X0 a_112_n50# a_n112_n147# a_n170_n50# w_n308_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1.12
C0 a_n170_n50# a_n112_n147# 0.0172f
C1 a_112_n50# w_n308_n269# 0.0232f
C2 a_112_n50# a_n170_n50# 0.0259f
C3 a_112_n50# a_n112_n147# 0.0172f
C4 w_n308_n269# a_n170_n50# 0.0232f
C5 w_n308_n269# a_n112_n147# 0.378f
C6 a_112_n50# VSUBS 0.0577f
C7 a_n170_n50# VSUBS 0.0577f
C8 a_n112_n147# VSUBS 0.389f
C9 w_n308_n269# VSUBS 1.14f
.ends

.subckt sky130_fd_pr__nfet_01v8_N39H2X a_n76_n100# a_n33_n188# a_18_n100# a_144_n240#
X0 a_18_n100# a_n33_n188# a_n76_n100# a_144_n240# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.18
C0 a_18_n100# a_n76_n100# 0.152f
C1 a_n33_n188# a_18_n100# 0.0205f
C2 a_n33_n188# a_n76_n100# 0.0205f
C3 a_18_n100# a_144_n240# 0.133f
C4 a_n76_n100# a_144_n240# 0.115f
C5 a_n33_n188# a_144_n240# 0.32f
.ends

.subckt th05 Vp V05 Vin m1_752_n794# Vn
XXM0 Vn m1_752_n794# Vn Vin sky130_fd_pr__nfet_01v8_Q7AWK3
XXM1 Vp Vin m1_752_n794# Vp Vn sky130_fd_pr__pfet_01v8_EXJYQP
XXM2 Vp Vp m1_752_n794# V05 Vn sky130_fd_pr__pfet_01v8_HJHF6N
XXM3 Vn m1_752_n794# V05 Vn sky130_fd_pr__nfet_01v8_N39H2X
C0 Vn m1_752_n794# 0.136f
C1 m1_752_n794# V05 0.0855f
C2 Vin Vp 0.139f
C3 Vn V05 0.0364f
C4 Vin m1_752_n794# 0.2f
C5 Vin Vn 0.041f
C6 Vin V05 0.00406f
C7 Vp m1_752_n794# 0.198f
C8 Vp Vn 0.0115f
C9 Vp V05 0.0548f
C10 V05 0 0.314f
C11 m1_752_n794# 0 0.788f
C12 Vp 0 2.28f
C13 Vin 0 0.905f
C14 Vn 0 0.547f
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X a_664_47# a_841_47#
+ a_381_47# a_62_47# a_558_47#
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPB X 0.126f
C1 VGND a_381_47# 0.125f
C2 X a_62_47# 0.156f
C3 VPB A 0.105f
C4 a_62_47# A 0.244f
C5 a_841_47# VPWR 0.0614f
C6 VPB a_664_47# 0.043f
C7 X A 0.0142f
C8 VPWR a_381_47# 0.134f
C9 VPB a_558_47# 0.115f
C10 VPWR VGND 0.0902f
C11 X a_664_47# 6.67e-19
C12 VPB a_841_47# 0.0108f
C13 a_558_47# X 0.0144f
C14 VPB a_381_47# 0.0447f
C15 a_558_47# a_664_47# 0.314f
C16 VPB VGND 0.008f
C17 VGND a_62_47# 0.144f
C18 X a_381_47# 0.318f
C19 a_841_47# a_664_47# 0.134f
C20 a_381_47# A 5.42e-19
C21 a_841_47# a_558_47# 0.00368f
C22 VGND X 0.106f
C23 VPB VPWR 0.103f
C24 VGND A 0.0176f
C25 VPWR a_62_47# 0.149f
C26 a_558_47# a_381_47# 0.16f
C27 VGND a_664_47# 0.125f
C28 VPWR X 0.108f
C29 a_558_47# VGND 0.0816f
C30 VPWR A 0.0174f
C31 VPB a_62_47# 0.0515f
C32 VPWR a_664_47# 0.131f
C33 a_841_47# VGND 0.0585f
C34 VPWR a_558_47# 0.084f
C35 VGND VNB 0.537f
C36 VPWR VNB 0.439f
C37 X VNB 0.163f
C38 A VNB 0.198f
C39 VPB VNB 0.959f
C40 a_841_47# VNB 0.0929f
C41 a_664_47# VNB 0.13f
C42 a_558_47# VNB 0.164f
C43 a_381_47# VNB 0.11f
C44 a_62_47# VNB 0.169f
.ends

.subckt sky130_fd_pr__nfet_01v8_4L9AWD a_n206_n182# a_n46_n130# a_n104_n42# a_46_n42#
X0 a_46_n42# a_n46_n130# a_n104_n42# a_n206_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.46
C0 a_n46_n130# a_n104_n42# 0.00852f
C1 a_46_n42# a_n104_n42# 0.0412f
C2 a_46_n42# a_n46_n130# 0.00852f
C3 a_46_n42# a_n206_n182# 0.0705f
C4 a_n104_n42# a_n206_n182# 0.0784f
C5 a_n46_n130# a_n206_n182# 0.388f
.ends

.subckt sky130_fd_pr__pfet_01v8_EZD9Q7 w_n224_n261# a_28_n42# a_n33_n139# a_n86_n42#
+ VSUBS
X0 a_28_n42# a_n33_n139# a_n86_n42# w_n224_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.28
C0 a_n86_n42# a_28_n42# 0.0541f
C1 w_n224_n261# a_n33_n139# 0.183f
C2 a_n33_n139# a_28_n42# 0.00625f
C3 w_n224_n261# a_28_n42# 0.0224f
C4 a_n86_n42# a_n33_n139# 0.00625f
C5 a_n86_n42# w_n224_n261# 0.0224f
C6 a_28_n42# VSUBS 0.0479f
C7 a_n86_n42# VSUBS 0.0479f
C8 a_n33_n139# VSUBS 0.155f
C9 w_n224_n261# VSUBS 0.799f
.ends

.subckt sky130_fd_pr__pfet_01v8_M479BZ a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n42# a_15_n42# 0.0699f
C1 w_n211_n261# a_n33_n139# 0.182f
C2 a_n33_n139# a_15_n42# 0.0192f
C3 w_n211_n261# a_15_n42# 0.0389f
C4 a_n73_n42# a_n33_n139# 0.0192f
C5 a_n73_n42# w_n211_n261# 0.016f
C6 a_15_n42# VSUBS 0.0328f
C7 a_n73_n42# VSUBS 0.0478f
C8 a_n33_n139# VSUBS 0.145f
C9 w_n211_n261# VSUBS 0.785f
.ends

.subckt sky130_fd_pr__nfet_01v8_4BNSKG a_n144_n216# a_18_n42# a_n33_n130# a_n76_n42#
X0 a_18_n42# a_n33_n130# a_n76_n42# a_n144_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.18
C0 a_n33_n130# a_n76_n42# 0.0154f
C1 a_18_n42# a_n76_n42# 0.0655f
C2 a_18_n42# a_n33_n130# 0.0154f
C3 a_18_n42# a_n144_n216# 0.0668f
C4 a_n76_n42# a_n144_n216# 0.0668f
C5 a_n33_n130# a_n144_n216# 0.319f
.ends

.subckt th10 V10 Vin m1_502_n495# m1_536_174# Vn Vp
XXM0 m1_502_n495# Vn Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vn Vin m1_536_174# m1_502_n495# sky130_fd_pr__nfet_01v8_4L9AWD
XXM2 Vp m1_536_174# Vin Vp Vn sky130_fd_pr__pfet_01v8_EZD9Q7
XXM3 Vp Vp m1_536_174# V10 Vn sky130_fd_pr__pfet_01v8_M479BZ
XXM4 Vn V10 m1_536_174# Vn sky130_fd_pr__nfet_01v8_4BNSKG
C0 Vin m1_502_n495# 0.0207f
C1 Vin Vp 0.175f
C2 m1_536_174# Vn 0.233f
C3 m1_502_n495# Vp 0.0256f
C4 Vn V10 0.0577f
C5 m1_536_174# V10 0.177f
C6 Vin Vn 0.114f
C7 Vin m1_536_174# 0.0971f
C8 Vin V10 0.0187f
C9 m1_502_n495# Vn 0.0348f
C10 m1_536_174# m1_502_n495# 0.00612f
C11 Vp Vn 0.102f
C12 m1_536_174# Vp 0.172f
C13 m1_502_n495# V10 0.042f
C14 Vp V10 0.0702f
C15 Vin 0 0.664f
C16 V10 0 0.249f
C17 Vn 0 0.463f
C18 m1_536_174# 0 0.825f
C19 Vp 0 2.17f
C20 m1_502_n495# 0 0.146f
.ends

.subckt sky130_fd_pr__nfet_01v8_X33H33 a_n73_n110# a_n175_n250# a_n33_n198# a_15_n110#
X0 a_15_n110# a_n33_n198# a_n73_n110# a_n175_n250# sky130_fd_pr__nfet_01v8 ad=0.319 pd=2.78 as=0.319 ps=2.78 w=1.1 l=0.15
C0 a_15_n110# a_n73_n110# 0.178f
C1 a_15_n110# a_n33_n198# 0.0261f
C2 a_n33_n198# a_n73_n110# 0.0261f
C3 a_15_n110# a_n175_n250# 0.121f
C4 a_n73_n110# a_n175_n250# 0.141f
C5 a_n33_n198# a_n175_n250# 0.32f
.ends

.subckt sky130_fd_pr__pfet_01v8_AMA9E4 a_n194_n44# a_n136_n141# w_n332_n263# a_136_n44#
+ VSUBS
X0 a_136_n44# a_n136_n141# a_n194_n44# w_n332_n263# sky130_fd_pr__pfet_01v8 ad=0.128 pd=1.46 as=0.128 ps=1.46 w=0.44 l=1.36
C0 a_n194_n44# a_n136_n141# 0.0174f
C1 a_n194_n44# a_136_n44# 0.0196f
C2 a_136_n44# a_n136_n141# 0.0174f
C3 a_n194_n44# w_n332_n263# 0.0226f
C4 w_n332_n263# a_n136_n141# 0.434f
C5 a_136_n44# w_n332_n263# 0.0226f
C6 a_136_n44# VSUBS 0.0532f
C7 a_n194_n44# VSUBS 0.0532f
C8 a_n136_n141# VSUBS 0.457f
C9 w_n332_n263# VSUBS 1.2f
.ends

.subckt sky130_fd_pr__pfet_01v8_8DZSNJ a_n74_n100# a_16_n100# w_n212_n319# a_n33_n197#
+ VSUBS
X0 a_16_n100# a_n33_n197# a_n74_n100# w_n212_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.16
C0 a_n74_n100# a_n33_n197# 0.0223f
C1 a_n74_n100# a_16_n100# 0.159f
C2 a_16_n100# a_n33_n197# 0.0223f
C3 a_n74_n100# w_n212_n319# 0.0252f
C4 w_n212_n319# a_n33_n197# 0.189f
C5 a_16_n100# w_n212_n319# 0.0252f
C6 a_16_n100# VSUBS 0.089f
C7 a_n74_n100# VSUBS 0.089f
C8 a_n33_n197# VSUBS 0.146f
C9 w_n212_n319# VSUBS 0.899f
.ends

.subckt th03 V03 Vin Vp m1_890_n844# m1_638_n591# Vn
XXM0 Vn Vn Vin m1_890_n844# sky130_fd_pr__nfet_01v8_X33H33
XXM1 m1_638_n591# Vin Vp m1_890_n844# Vn sky130_fd_pr__pfet_01v8_AMA9E4
XXM2 Vp Vn Vp m1_638_n591# sky130_fd_pr__nfet_01v8_LH5FDA
XXM3 Vp V03 Vp m1_890_n844# Vn sky130_fd_pr__pfet_01v8_8DZSNJ
XXM4 m1_890_n844# Vn Vn V03 sky130_fd_pr__nfet_01v8_LH5FDA
C0 Vin Vp 0.313f
C1 Vn Vin 0.105f
C2 V03 m1_890_n844# 0.129f
C3 m1_638_n591# m1_890_n844# 0.0187f
C4 Vn Vp 0.023f
C5 Vin m1_890_n844# 0.188f
C6 V03 Vin 0.0036f
C7 Vp m1_890_n844# 0.459f
C8 Vn m1_890_n844# 0.183f
C9 Vin m1_638_n591# 0.0439f
C10 V03 Vp 0.0492f
C11 Vn V03 0.0337f
C12 Vp m1_638_n591# 0.169f
C13 Vn m1_638_n591# 0.0097f
C14 Vp 0 3.07f
C15 V03 0 0.308f
C16 Vn 0 0.446f
C17 m1_890_n844# 0 1.05f
C18 m1_638_n591# 0 0.224f
C19 Vin 0 0.924f
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y a_129_47# a_47_47# a_285_47#
+ a_377_297#
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VGND a_285_47# 0.211f
C1 Y VGND 0.0381f
C2 VPWR a_285_47# 0.00255f
C3 VPB A 0.0822f
C4 Y VPWR 0.107f
C5 a_377_297# a_47_47# 0.00899f
C6 B A 0.236f
C7 VGND A 0.0635f
C8 VPWR A 0.0349f
C9 B a_129_47# 0.00236f
C10 a_285_47# a_47_47# 0.0175f
C11 Y a_377_297# 0.00188f
C12 VPB B 0.0643f
C13 Y a_47_47# 0.143f
C14 VGND a_129_47# 0.00547f
C15 VPB VGND 0.00568f
C16 VPWR a_129_47# 9.47e-19
C17 VPB VPWR 0.0718f
C18 B VGND 0.0389f
C19 Y a_285_47# 0.0439f
C20 A a_47_47# 0.0307f
C21 B VPWR 0.0408f
C22 VGND VPWR 0.0665f
C23 a_129_47# a_47_47# 0.00369f
C24 VPB a_47_47# 0.0444f
C25 A a_285_47# 0.0353f
C26 Y A 0.00181f
C27 B a_377_297# 0.00254f
C28 B a_47_47# 0.356f
C29 VGND a_377_297# 0.00125f
C30 VGND a_47_47# 0.104f
C31 VPB a_285_47# 5.53e-19
C32 a_377_297# VPWR 0.00559f
C33 Y VPB 0.00878f
C34 VPWR a_47_47# 0.273f
C35 B a_285_47# 0.067f
C36 Y B 0.00334f
C37 VGND VNB 0.4f
C38 Y VNB 0.0783f
C39 VPWR VNB 0.352f
C40 A VNB 0.217f
C41 B VNB 0.212f
C42 VPB VNB 0.693f
C43 a_285_47# VNB 0.0174f
C44 a_47_47# VNB 0.199f
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X a_472_297# a_80_21#
+ a_300_47# a_217_297#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
C0 B1 VGND 0.0175f
C1 a_217_297# a_472_297# 0.00517f
C2 a_80_21# A2 0.128f
C3 VGND A2 0.0191f
C4 A1 VPWR 0.0149f
C5 B1 A1 0.0834f
C6 a_217_297# a_80_21# 0.127f
C7 C1 a_80_21# 0.079f
C8 a_217_297# VGND 0.00342f
C9 a_300_47# VPWR 8.53e-19
C10 A1 A2 0.0881f
C11 VGND C1 0.0176f
C12 a_217_297# A1 0.0124f
C13 B1 VPWR 0.0129f
C14 VPB X 0.0118f
C15 VPWR A2 0.0161f
C16 a_217_297# VPWR 0.197f
C17 VPB a_80_21# 0.0661f
C18 VPWR C1 0.0137f
C19 a_217_297# B1 0.00651f
C20 B1 C1 0.0846f
C21 VGND VPB 0.00775f
C22 a_472_297# X 2.6e-19
C23 a_217_297# A2 0.0135f
C24 A1 VPB 0.0266f
C25 a_80_21# X 0.118f
C26 a_217_297# C1 0.00262f
C27 VGND X 0.0654f
C28 a_472_297# a_80_21# 0.0164f
C29 VGND a_472_297# 0.00188f
C30 A1 X 3.62e-19
C31 VGND a_80_21# 0.293f
C32 VPWR VPB 0.0754f
C33 B1 VPB 0.0267f
C34 a_300_47# X 5.31e-19
C35 VPB A2 0.0384f
C36 A1 a_80_21# 0.111f
C37 VGND A1 0.0147f
C38 VPWR X 0.0884f
C39 a_217_297# VPB 0.00494f
C40 B1 X 1.18e-19
C41 a_300_47# a_80_21# 0.00997f
C42 VPWR a_472_297# 0.00703f
C43 C1 VPB 0.0379f
C44 VGND a_300_47# 0.00536f
C45 B1 a_472_297# 1.87e-19
C46 X A2 6.82e-19
C47 VPWR a_80_21# 0.119f
C48 B1 a_80_21# 0.0964f
C49 a_217_297# X 0.00271f
C50 VGND VPWR 0.0665f
C51 A1 a_300_47# 5.95e-19
C52 C1 X 7.15e-20
C53 VGND VNB 0.385f
C54 VPWR VNB 0.325f
C55 X VNB 0.0899f
C56 C1 VNB 0.144f
C57 B1 VNB 0.0899f
C58 A1 VNB 0.0905f
C59 A2 VNB 0.108f
C60 VPB VNB 0.693f
C61 a_217_297# VNB 0.00117f
C62 a_80_21# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
C0 X D 0.00746f
C1 X VPB 0.0111f
C2 B VGND 0.0453f
C3 A VGND 0.0151f
C4 D VGND 0.0898f
C5 VPB VGND 0.00852f
C6 VGND a_197_47# 0.00387f
C7 A B 0.0839f
C8 a_27_47# a_303_47# 0.00119f
C9 B VPB 0.0643f
C10 B a_197_47# 0.00623f
C11 A VPB 0.0907f
C12 a_303_47# C 0.00527f
C13 D VPB 0.0782f
C14 a_27_47# C 0.0516f
C15 a_303_47# VPWR 4.83e-19
C16 a_27_47# VPWR 0.326f
C17 a_27_47# a_109_47# 0.00578f
C18 C VPWR 0.021f
C19 C a_109_47# 1.72e-20
C20 a_109_47# VPWR 4.66e-19
C21 a_27_47# X 0.0754f
C22 a_303_47# VGND 0.00381f
C23 a_27_47# VGND 0.132f
C24 C VGND 0.0408f
C25 X VPWR 0.0945f
C26 a_27_47# B 0.13f
C27 a_303_47# D 0.00119f
C28 a_27_47# A 0.153f
C29 VGND VPWR 0.0662f
C30 a_27_47# D 0.107f
C31 a_109_47# VGND 0.00223f
C32 a_27_47# VPB 0.082f
C33 C B 0.161f
C34 a_27_47# a_197_47# 0.00167f
C35 C D 0.18f
C36 C VPB 0.0609f
C37 B VPWR 0.0231f
C38 a_109_47# B 0.00153f
C39 C a_197_47# 0.00123f
C40 A VPWR 0.044f
C41 D VPWR 0.0207f
C42 VPB VPWR 0.077f
C43 X VGND 0.0903f
C44 a_197_47# VPWR 5.24e-19
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt sky130_fd_pr__nfet_01v8_SHU4BF a_n73_n353# a_n141_493# a_15_n353# a_n33_n441#
X0 a_15_n353# a_n33_n441# a_n73_n353# a_n141_493# sky130_fd_pr__nfet_01v8 ad=1.02 pd=7.64 as=1.02 ps=7.64 w=3.53 l=0.15
C0 a_15_n353# a_n33_n441# 0.0384f
C1 a_15_n353# a_n73_n353# 0.564f
C2 a_n33_n441# a_n73_n353# 0.0384f
C3 a_15_n353# a_n141_493# 0.327f
C4 a_n73_n353# a_n141_493# 0.327f
C5 a_n33_n441# a_n141_493# 0.329f
.ends

.subckt sky130_fd_pr__pfet_01v8_HE9GT9 a_n408_n42# a_350_n42# w_n546_n261# a_n350_n139#
+ VSUBS
X0 a_350_n42# a_n350_n139# a_n408_n42# w_n546_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 a_n408_n42# w_n546_n261# 0.0408f
C1 w_n546_n261# a_350_n42# 0.0179f
C2 a_n408_n42# a_n350_n139# 0.0226f
C3 a_350_n42# a_n350_n139# 0.0226f
C4 w_n546_n261# a_n350_n139# 0.756f
C5 a_n408_n42# a_350_n42# 0.00807f
C6 a_350_n42# VSUBS 0.0587f
C7 a_n408_n42# VSUBS 0.0437f
C8 a_n350_n139# VSUBS 1.19f
C9 w_n546_n261# VSUBS 1.83f
.ends

.subckt sky130_fd_pr__nfet_01v8_LHD8GA a_n408_n42# a_350_n42# a_n350_n130# a_n510_n182#
X0 a_350_n42# a_n350_n130# a_n408_n42# a_n510_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.5
C0 a_350_n42# a_n350_n130# 0.0226f
C1 a_350_n42# a_n408_n42# 0.00807f
C2 a_n350_n130# a_n408_n42# 0.0226f
C3 a_350_n42# a_n510_n182# 0.0766f
C4 a_n408_n42# a_n510_n182# 0.0845f
C5 a_n350_n130# a_n510_n182# 1.9f
.ends

.subckt th01 V01 Vn m1_991_n1219# m1_571_n501# Vp Vin
XXM0 Vn Vn m1_991_n1219# Vin sky130_fd_pr__nfet_01v8_SHU4BF
XXM1 m1_571_n501# m1_991_n1219# Vp Vin Vn sky130_fd_pr__pfet_01v8_HE9GT9
XXM2 Vp m1_571_n501# Vp Vn sky130_fd_pr__nfet_01v8_LHD8GA
XXM3 Vp Vp V01 m1_991_n1219# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 m1_991_n1219# Vn V01 Vn sky130_fd_pr__nfet_01v8_LH5FDA
C0 Vn V01 0.0149f
C1 Vp V01 0.0684f
C2 m1_571_n501# m1_991_n1219# 0.0899f
C3 m1_991_n1219# Vin 0.208f
C4 m1_571_n501# Vin 0.274f
C5 Vn m1_991_n1219# 0.0569f
C6 m1_991_n1219# Vp 0.423f
C7 m1_571_n501# Vn 2.57e-20
C8 Vn Vin 0.0582f
C9 m1_571_n501# Vp 0.32f
C10 Vp Vin 0.354f
C11 m1_991_n1219# V01 0.0901f
C12 m1_571_n501# V01 2.16e-20
C13 V01 Vin 0.00412f
C14 Vn Vp 0.0233f
C15 Vn 0 0.633f
C16 V01 0 0.373f
C17 m1_991_n1219# 0 1.24f
C18 Vp 0 4.41f
C19 m1_571_n501# 0 0.194f
C20 Vin 0 1.87f
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X a_489_413# a_226_47#
+ a_556_47# a_226_297# a_76_199#
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPB a_76_199# 0.0817f
C1 VPWR a_489_413# 0.143f
C2 VPWR X 0.0589f
C3 VGND B1 0.0471f
C4 VGND B2 0.0335f
C5 A1_N A2_N 0.11f
C6 VPWR a_556_47# 7.24e-19
C7 VGND A2_N 0.0174f
C8 A1_N X 0.00211f
C9 a_76_199# VPWR 0.2f
C10 VGND a_489_413# 0.0058f
C11 a_76_199# a_226_297# 0.00354f
C12 VGND X 0.0627f
C13 B1 B2 0.182f
C14 VPB a_226_47# 0.111f
C15 a_76_199# A1_N 0.119f
C16 VGND a_556_47# 0.00639f
C17 VGND a_76_199# 0.108f
C18 a_489_413# B2 0.0541f
C19 B1 a_489_413# 0.0382f
C20 a_226_47# VPWR 0.0187f
C21 a_556_47# B2 0.00291f
C22 VPB VPWR 0.0951f
C23 a_226_47# a_226_297# 0.00128f
C24 X A2_N 2.55e-19
C25 a_76_199# B1 0.00185f
C26 a_76_199# B2 0.0626f
C27 a_226_47# A1_N 0.0209f
C28 VPB A1_N 0.0339f
C29 VGND a_226_47# 0.149f
C30 a_76_199# A2_N 0.0125f
C31 VPB VGND 0.0128f
C32 a_76_199# a_489_413# 0.0473f
C33 VPWR a_226_297# 8.54e-19
C34 a_76_199# X 0.0995f
C35 a_76_199# a_556_47# 0.0017f
C36 A1_N VPWR 0.00672f
C37 a_226_47# B2 0.0975f
C38 A1_N a_226_297# 0.00184f
C39 VGND VPWR 0.0743f
C40 VPB B2 0.0645f
C41 VPB B1 0.0803f
C42 VGND a_226_297# 5.63e-19
C43 a_226_47# A2_N 0.141f
C44 VPB A2_N 0.0327f
C45 a_226_47# a_489_413# 0.00579f
C46 VGND A1_N 0.0261f
C47 a_226_47# X 0.0108f
C48 VPB a_489_413# 0.015f
C49 VPB X 0.0113f
C50 VPWR B1 0.0188f
C51 VPWR B2 0.0161f
C52 a_76_199# a_226_47# 0.188f
C53 VPWR A2_N 0.00449f
C54 VGND VNB 0.462f
C55 A2_N VNB 0.103f
C56 A1_N VNB 0.111f
C57 VPWR VNB 0.369f
C58 X VNB 0.0975f
C59 B1 VNB 0.206f
C60 B2 VNB 0.106f
C61 VPB VNB 0.782f
C62 a_489_413# VNB 0.0254f
C63 a_226_47# VNB 0.162f
C64 a_76_199# VNB 0.141f
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X a_515_93# a_223_47#
+ a_615_93# a_343_93# a_429_93# a_27_47#
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
C0 VPWR VGND 0.0906f
C1 VPWR a_429_93# 5.19e-19
C2 B_N A_N 0.117f
C3 a_223_47# C 0.151f
C4 a_343_93# a_223_47# 0.269f
C5 VPWR a_615_93# 8.49e-19
C6 a_515_93# VGND 0.00408f
C7 VPWR D 0.0143f
C8 a_223_47# VGND 0.199f
C9 a_429_93# a_223_47# 0.00492f
C10 A_N VGND 0.0146f
C11 VPWR a_27_47# 0.0897f
C12 a_223_47# D 4.03e-19
C13 B_N VPB 0.0646f
C14 VPB X 0.0103f
C15 VPWR a_515_93# 7.86e-19
C16 VPB C 0.0686f
C17 a_27_47# a_223_47# 0.267f
C18 a_343_93# VPB 0.0857f
C19 VPWR a_223_47# 0.114f
C20 a_27_47# A_N 0.0906f
C21 VPB VGND 0.0167f
C22 VPWR A_N 0.0318f
C23 a_223_47# a_515_93# 0.00482f
C24 B_N X 4.64e-20
C25 B_N C 9.56e-20
C26 B_N a_343_93# 0.00112f
C27 a_343_93# X 0.126f
C28 VPB D 0.081f
C29 a_343_93# C 0.0397f
C30 a_223_47# A_N 0.00833f
C31 B_N VGND 0.0427f
C32 X VGND 0.0609f
C33 a_27_47# VPB 0.154f
C34 C VGND 0.025f
C35 a_343_93# VGND 0.0548f
C36 VPWR VPB 0.106f
C37 a_429_93# a_343_93# 0.00484f
C38 B_N D 6.67e-20
C39 a_615_93# C 0.00407f
C40 a_615_93# a_343_93# 0.00103f
C41 X D 0.0193f
C42 a_429_93# VGND 0.00122f
C43 D C 0.163f
C44 a_343_93# D 0.114f
C45 a_223_47# VPB 0.0799f
C46 B_N a_27_47# 0.138f
C47 VPWR B_N 0.0168f
C48 a_615_93# VGND 0.0044f
C49 VPWR X 0.0582f
C50 VPB A_N 0.0848f
C51 D VGND 0.0414f
C52 a_343_93# a_27_47# 0.0406f
C53 VPWR C 0.012f
C54 VPWR a_343_93# 0.255f
C55 a_615_93# D 0.00564f
C56 B_N a_223_47# 0.0431f
C57 a_27_47# VGND 0.0715f
C58 a_515_93# C 0.00389f
C59 a_343_93# a_515_93# 0.00115f
C60 VGND VNB 0.553f
C61 X VNB 0.0908f
C62 VPWR VNB 0.453f
C63 D VNB 0.124f
C64 C VNB 0.107f
C65 B_N VNB 0.134f
C66 A_N VNB 0.144f
C67 VPB VNB 0.959f
C68 a_343_93# VNB 0.172f
C69 a_223_47# VNB 0.141f
C70 a_27_47# VNB 0.259f
.ends

.subckt sky130_fd_pr__pfet_01v8_MWHFPY a_n73_n63# a_n33_n160# w_n211_n282# a_15_n63#
+ VSUBS
X0 a_15_n63# a_n33_n160# a_n73_n63# w_n211_n282# sky130_fd_pr__pfet_01v8 ad=0.183 pd=1.84 as=0.183 ps=1.84 w=0.63 l=0.15
C0 a_15_n63# a_n73_n63# 0.103f
C1 w_n211_n282# a_n33_n160# 0.237f
C2 w_n211_n282# a_n73_n63# 0.0591f
C3 a_n73_n63# a_n33_n160# 0.021f
C4 a_15_n63# w_n211_n282# 0.0591f
C5 a_15_n63# a_n33_n160# 0.021f
C6 a_15_n63# VSUBS 0.0348f
C7 a_n73_n63# VSUBS 0.0348f
C8 a_n33_n160# VSUBS 0.116f
C9 w_n211_n282# VSUBS 1.1f
.ends

.subckt sky130_fd_pr__nfet_01v8_DPSGWY a_350_n100# a_n408_n100# a_n350_n188# a_n510_n274#
X0 a_350_n100# a_n350_n188# a_n408_n100# a_n510_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3.5
C0 a_n350_n188# a_n408_n100# 0.0439f
C1 a_n350_n188# a_350_n100# 0.0439f
C2 a_350_n100# a_n408_n100# 0.0188f
C3 a_350_n100# a_n510_n274# 0.159f
C4 a_n408_n100# a_n510_n274# 0.159f
C5 a_n350_n188# a_n510_n274# 2.13f
.ends

.subckt preamp Vin Vpamp Vn Vp
XXM0 Vn Vin Vp Vpamp Vn sky130_fd_pr__pfet_01v8_MWHFPY
XXM1 Vpamp Vp Vin Vn sky130_fd_pr__nfet_01v8_DPSGWY
C0 Vp Vin 0.324f
C1 Vp Vn 0.297f
C2 Vpamp Vin 0.0777f
C3 Vpamp Vn 0.047f
C4 Vpamp Vp 0.0552f
C5 Vn Vin 0.29f
C6 Vn 0 0.193f
C7 Vpamp 0 0.444f
C8 Vp 0 1.53f
C9 Vin 0 2.21f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 X a_117_297# 2.25e-19
C1 a_285_47# X 0.00206f
C2 X a_285_297# 0.0712f
C3 X VGND 0.173f
C4 a_35_297# A 0.0633f
C5 VPB a_285_297# 0.0133f
C6 VPB VGND 0.00696f
C7 VGND a_117_297# 0.00177f
C8 A B 0.221f
C9 a_35_297# B 0.203f
C10 a_285_47# VGND 0.00552f
C11 VGND a_285_297# 0.00394f
C12 A VPWR 0.0348f
C13 a_35_297# VPWR 0.096f
C14 VPWR B 0.0703f
C15 A X 0.00166f
C16 a_35_297# X 0.166f
C17 X B 0.0149f
C18 A VPB 0.051f
C19 X VPWR 0.0537f
C20 a_35_297# VPB 0.0699f
C21 a_35_297# a_117_297# 0.00641f
C22 VPB B 0.0697f
C23 B a_117_297# 0.00777f
C24 A a_285_297# 0.00749f
C25 A VGND 0.0325f
C26 a_35_297# a_285_47# 0.00723f
C27 a_35_297# a_285_297# 0.025f
C28 a_35_297# VGND 0.177f
C29 VPWR VPB 0.0689f
C30 a_285_47# B 3.98e-19
C31 B a_285_297# 0.0553f
C32 VGND B 0.0304f
C33 VPWR a_117_297# 0.00852f
C34 a_285_47# VPWR 8.6e-19
C35 X VPB 0.0154f
C36 VPWR a_285_297# 0.246f
C37 VPWR VGND 0.0643f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt sky130_fd_pr__pfet_01v8_LDQF7K a_n33_n147# a_29_n50# a_n87_n50# w_n225_n269#
+ VSUBS
X0 a_29_n50# a_n33_n147# a_n87_n50# w_n225_n269# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.29
C0 w_n225_n269# a_n33_n147# 0.176f
C1 a_n87_n50# a_n33_n147# 0.00691f
C2 w_n225_n269# a_29_n50# 0.0186f
C3 a_n87_n50# a_29_n50# 0.0628f
C4 a_n87_n50# w_n225_n269# 0.0457f
C5 a_n33_n147# a_29_n50# 0.00691f
C6 a_29_n50# VSUBS 0.0581f
C7 a_n87_n50# VSUBS 0.0403f
C8 a_n33_n147# VSUBS 0.158f
C9 w_n225_n269# VSUBS 0.854f
.ends

.subckt sky130_fd_pr__nfet_01v8_HZA4VB a_326_n230# a_n200_n130# a_200_n42# li_n360_158#
+ a_n258_n42#
X0 a_200_n42# a_n200_n130# a_n258_n42# a_326_n230# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_n200_n130# a_n258_n42# 0.0196f
C1 a_200_n42# a_n258_n42# 0.0134f
C2 a_200_n42# a_n200_n130# 0.0196f
C3 li_n360_158# a_326_n230# 0.0244f
C4 a_200_n42# a_326_n230# 0.0748f
C5 a_n258_n42# a_326_n230# 0.0746f
C6 a_n200_n130# a_326_n230# 1.15f
.ends

.subckt sky130_fd_pr__pfet_01v8_GEY2B5 w_n275_n270# a_n137_n51# a_79_n51# a_n79_n148#
+ VSUBS
X0 a_79_n51# a_n79_n148# a_n137_n51# w_n275_n270# sky130_fd_pr__pfet_01v8 ad=0.148 pd=1.6 as=0.148 ps=1.6 w=0.51 l=0.79
C0 w_n275_n270# a_n79_n148# 0.294f
C1 a_n137_n51# a_n79_n148# 0.0141f
C2 w_n275_n270# a_79_n51# 0.0232f
C3 a_n137_n51# a_79_n51# 0.0345f
C4 a_n137_n51# w_n275_n270# 0.0232f
C5 a_n79_n148# a_79_n51# 0.0141f
C6 a_79_n51# VSUBS 0.0573f
C7 a_n137_n51# VSUBS 0.0573f
C8 a_n79_n148# VSUBS 0.294f
C9 w_n275_n270# VSUBS 1.01f
.ends

.subckt sky130_fd_pr__pfet_01v8_KQKFM4 w_n526_n261# a_n330_n139# a_330_n42# a_n388_n42#
+ VSUBS
X0 a_330_n42# a_n330_n139# a_n388_n42# w_n526_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.3
C0 w_n526_n261# a_n330_n139# 0.911f
C1 a_n388_n42# a_n330_n139# 0.0223f
C2 w_n526_n261# a_330_n42# 0.0224f
C3 a_n388_n42# a_330_n42# 0.00853f
C4 a_n388_n42# w_n526_n261# 0.0224f
C5 a_n330_n139# a_330_n42# 0.0223f
C6 a_330_n42# VSUBS 0.0545f
C7 a_n388_n42# VSUBS 0.0545f
C8 a_n330_n139# VSUBS 1.02f
C9 w_n526_n261# VSUBS 1.89f
.ends

.subckt sky130_fd_pr__nfet_01v8_5NW376 a_n73_n251# a_n141_391# a_15_n251# a_n33_n339#
X0 a_15_n251# a_n33_n339# a_n73_n251# a_n141_391# sky130_fd_pr__nfet_01v8 ad=0.728 pd=5.6 as=0.728 ps=5.6 w=2.51 l=0.15
C0 a_n33_n339# a_n73_n251# 0.0337f
C1 a_15_n251# a_n73_n251# 0.402f
C2 a_15_n251# a_n33_n339# 0.0337f
C3 a_15_n251# a_n141_391# 0.241f
C4 a_n73_n251# a_n141_391# 0.241f
C5 a_n33_n339# a_n141_391# 0.327f
.ends

.subckt th15 V15 Vin m1_597_n912# m1_849_n157# Vp Vn
XXM0 Vn Vn m1_597_n912# Vp Vn sky130_fd_pr__pfet_01v8_LDQF7K
XXM1 Vn Vin m1_849_n157# Vn m1_597_n912# sky130_fd_pr__nfet_01v8_HZA4VB
XXM2 Vp Vp m1_849_n157# Vin Vn sky130_fd_pr__pfet_01v8_GEY2B5
XXM3 Vp m1_849_n157# V15 Vp Vn sky130_fd_pr__pfet_01v8_KQKFM4
XXM4 Vn Vn V15 m1_849_n157# sky130_fd_pr__nfet_01v8_5NW376
C0 m1_849_n157# V15 0.202f
C1 m1_849_n157# Vn 0.171f
C2 Vn V15 2.72e-19
C3 m1_849_n157# m1_597_n912# 0.00715f
C4 m1_849_n157# Vp 0.226f
C5 Vp V15 0.0762f
C6 Vn m1_597_n912# 0.175f
C7 Vn Vp 0.0678f
C8 m1_849_n157# Vin 0.0977f
C9 Vin V15 0.00573f
C10 Vp m1_597_n912# 0.0557f
C11 Vin Vn 0.38f
C12 Vin m1_597_n912# 0.211f
C13 Vin Vp 0.166f
C14 V15 0 0.332f
C15 Vn 0 0.276f
C16 m1_849_n157# 0 1.28f
C17 Vp 0 3.52f
C18 m1_597_n912# 0 0.19f
C19 Vin 0 1.58f
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X a_465_297# a_297_297#
+ a_215_297# a_392_297# a_109_53#
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 C a_215_297# 0.161f
C1 a_109_53# a_297_297# 7.06e-21
C2 a_109_53# a_215_297# 0.0807f
C3 C A 0.0281f
C4 D_N a_109_53# 0.0889f
C5 a_297_297# VPWR 8.59e-19
C6 a_109_53# A 1.19e-19
C7 VPWR a_215_297# 0.0871f
C8 VPB B 0.116f
C9 D_N VPWR 0.0412f
C10 C a_392_297# 0.00267f
C11 VPB X 0.011f
C12 A VPWR 0.0073f
C13 a_297_297# a_215_297# 0.00659f
C14 D_N a_215_297# 3.19e-19
C15 C VGND 0.0202f
C16 VPWR a_392_297# 5.29e-19
C17 A a_215_297# 0.157f
C18 a_109_53# VGND 0.118f
C19 a_392_297# a_215_297# 0.00419f
C20 VPWR VGND 0.075f
C21 C B 0.0893f
C22 a_297_297# VGND 6.5e-19
C23 a_109_53# B 0.0246f
C24 VGND a_215_297# 0.237f
C25 D_N VGND 0.0531f
C26 C a_465_297# 6.89e-19
C27 B VPWR 0.255f
C28 A VGND 0.0158f
C29 X VPWR 0.0885f
C30 VPB C 0.0337f
C31 VGND a_392_297# 3.44e-19
C32 VPWR a_465_297# 7.08e-19
C33 B a_215_297# 0.159f
C34 VPB a_109_53# 0.0547f
C35 X a_215_297# 0.0991f
C36 A B 0.0666f
C37 VPB VPWR 0.122f
C38 a_215_297# a_465_297# 0.00827f
C39 X A 0.00127f
C40 A a_465_297# 5.42e-19
C41 VPB a_215_297# 0.0508f
C42 VPB D_N 0.0461f
C43 VPB A 0.0325f
C44 B VGND 0.0161f
C45 a_109_53# C 0.0984f
C46 X VGND 0.0359f
C47 VGND a_465_297# 5.02e-19
C48 C VPWR 0.00753f
C49 a_109_53# VPWR 0.0418f
C50 VPB VGND 0.0115f
C51 C a_297_297# 0.00375f
C52 X B 6.65e-19
C53 VGND VNB 0.469f
C54 X VNB 0.0884f
C55 A VNB 0.108f
C56 C VNB 0.101f
C57 D_N VNB 0.185f
C58 B VNB 0.101f
C59 VPWR VNB 0.399f
C60 VPB VNB 0.782f
C61 a_109_53# VNB 0.159f
C62 a_215_297# VNB 0.142f
.ends

.subckt sky130_fd_pr__nfet_01v8_JSJ4VK a_113_n42# a_n239_n216# a_n171_n42# a_n113_n130#
X0 a_113_n42# a_n113_n130# a_n171_n42# a_n239_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.13
C0 a_n113_n130# a_n171_n42# 0.0154f
C1 a_n171_n42# a_113_n42# 0.0218f
C2 a_n113_n130# a_113_n42# 0.0154f
C3 a_113_n42# a_n239_n216# 0.0734f
C4 a_n171_n42# a_n239_n216# 0.0734f
C5 a_n113_n130# a_n239_n216# 0.746f
.ends

.subckt sky130_fd_pr__pfet_01v8_EVXEQ2 a_16_n67# a_n33_n164# a_n74_n67# w_n212_n286#
+ VSUBS
X0 a_16_n67# a_n33_n164# a_n74_n67# w_n212_n286# sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.92 as=0.194 ps=1.92 w=0.67 l=0.16
C0 w_n212_n286# a_n33_n164# 0.183f
C1 a_n33_n164# a_n74_n67# 0.0198f
C2 w_n212_n286# a_n74_n67# 0.0184f
C3 a_16_n67# a_n33_n164# 0.0198f
C4 w_n212_n286# a_16_n67# 0.0544f
C5 a_16_n67# a_n74_n67# 0.107f
C6 a_16_n67# VSUBS 0.0435f
C7 a_n74_n67# VSUBS 0.0673f
C8 a_n33_n164# VSUBS 0.147f
C9 w_n212_n286# VSUBS 0.864f
.ends

.subckt sky130_fd_pr__pfet_01v8_BBE9QE w_n244_n262# a_n106_n43# a_48_n43# a_n48_n140#
+ VSUBS
X0 a_48_n43# a_n48_n140# a_n106_n43# w_n244_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.48
C0 w_n244_n262# a_n48_n140# 0.218f
C1 a_n48_n140# a_n106_n43# 0.00893f
C2 w_n244_n262# a_n106_n43# 0.0225f
C3 a_48_n43# a_n48_n140# 0.00893f
C4 w_n244_n262# a_48_n43# 0.0225f
C5 a_48_n43# a_n106_n43# 0.041f
C6 a_48_n43# VSUBS 0.0495f
C7 a_n106_n43# VSUBS 0.0495f
C8 a_n48_n140# VSUBS 0.203f
C9 w_n244_n262# VSUBS 0.876f
.ends

.subckt sky130_fd_pr__nfet_01v8_NCP4B2 a_n73_n47# a_n141_n221# a_n33_n135# a_15_n47#
X0 a_15_n47# a_n33_n135# a_n73_n47# a_n141_n221# sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.52 as=0.136 ps=1.52 w=0.47 l=0.15
C0 a_n33_n135# a_n73_n47# 0.0213f
C1 a_n73_n47# a_15_n47# 0.0779f
C2 a_n33_n135# a_15_n47# 0.0213f
C3 a_15_n47# a_n141_n221# 0.0686f
C4 a_n73_n47# a_n141_n221# 0.0686f
C5 a_n33_n135# a_n141_n221# 0.317f
.ends

.subckt th08 Vp Vin V08 m1_477_n803# Vn
XXM0 Vn Vn m1_477_n803# Vin sky130_fd_pr__nfet_01v8_JSJ4VK
XXM1 Vp Vin m1_477_n803# Vp Vn sky130_fd_pr__pfet_01v8_EVXEQ2
XXM2 Vp Vp V08 m1_477_n803# Vn sky130_fd_pr__pfet_01v8_BBE9QE
XXM3 Vn Vn m1_477_n803# V08 sky130_fd_pr__nfet_01v8_NCP4B2
C0 Vp V08 0.0461f
C1 Vp Vin 0.0933f
C2 m1_477_n803# V08 0.108f
C3 m1_477_n803# Vin 0.356f
C4 m1_477_n803# Vp 0.154f
C5 V08 Vin 0.00163f
C6 Vp Vn 1.66f
C7 m1_477_n803# Vn 0.656f
C8 Vin Vn 1.02f
C9 V08 Vn 0.271f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFRTVB a_n410_n216# a_n250_n130# a_n308_n42# a_250_n42#
X0 a_250_n42# a_n250_n130# a_n308_n42# a_n410_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.5
C0 a_n308_n42# a_250_n42# 0.011f
C1 a_n308_n42# a_n250_n130# 0.0209f
C2 a_250_n42# a_n250_n130# 0.0209f
C3 a_250_n42# a_n410_n216# 0.0852f
C4 a_n308_n42# a_n410_n216# 0.0853f
C5 a_n250_n130# a_n410_n216# 1.48f
.ends

.subckt sky130_fd_pr__pfet_01v8_XQZLDL a_15_n240# w_n211_n459# a_n73_n240# a_n33_n337#
+ VSUBS
X0 a_15_n240# a_n33_n337# a_n73_n240# w_n211_n459# sky130_fd_pr__pfet_01v8 ad=0.696 pd=5.38 as=0.696 ps=5.38 w=2.4 l=0.15
C0 a_n33_n337# a_n73_n240# 0.0313f
C1 a_n33_n337# w_n211_n459# 0.206f
C2 a_n73_n240# a_15_n240# 0.385f
C3 w_n211_n459# a_15_n240# 0.163f
C4 a_n33_n337# a_15_n240# 0.0313f
C5 a_n73_n240# w_n211_n459# 0.0371f
C6 a_15_n240# VSUBS 0.11f
C7 a_n73_n240# VSUBS 0.195f
C8 a_n33_n337# VSUBS 0.139f
C9 w_n211_n459# VSUBS 1.47f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GC6 a_200_n42# w_n396_n261# a_n200_n139# a_n258_n42#
+ VSUBS
X0 a_200_n42# a_n200_n139# a_n258_n42# w_n396_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_n200_n139# a_n258_n42# 0.0196f
C1 a_n200_n139# w_n396_n261# 0.73f
C2 a_n258_n42# a_200_n42# 0.0134f
C3 w_n396_n261# a_200_n42# 0.0498f
C4 a_n200_n139# a_200_n42# 0.0196f
C5 a_n258_n42# w_n396_n261# 0.0269f
C6 a_200_n42# VSUBS 0.0338f
C7 a_n258_n42# VSUBS 0.0488f
C8 a_n200_n139# VSUBS 0.563f
C9 w_n396_n261# VSUBS 1.69f
.ends

.subckt sky130_fd_pr__nfet_01v8_ATLS57 a_15_n200# a_n73_n200# a_n33_n288# a_n141_n374#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n141_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n73_n200# a_15_n200# 0.321f
C1 a_n73_n200# a_n33_n288# 0.0312f
C2 a_15_n200# a_n33_n288# 0.0312f
C3 a_15_n200# a_n141_n374# 0.233f
C4 a_n73_n200# a_n141_n374# 0.199f
C5 a_n33_n288# a_n141_n374# 0.341f
.ends

.subckt th13 V13 Vin m1_831_275# Vn m1_559_n458# Vp
XXM0 Vn m1_559_n458# Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vn Vin m1_559_n458# m1_831_275# sky130_fd_pr__nfet_01v8_ZFRTVB
XXM2 Vp Vp m1_831_275# Vin Vn sky130_fd_pr__pfet_01v8_XQZLDL
XXM3 V13 Vp m1_831_275# Vp Vn sky130_fd_pr__pfet_01v8_VZ9GC6
XXM4 V13 Vn m1_831_275# Vn sky130_fd_pr__nfet_01v8_ATLS57
C0 Vp Vn 0.206f
C1 Vp V13 0.135f
C2 m1_559_n458# Vn 0.152f
C3 Vin m1_831_275# 0.197f
C4 V13 Vn 0.0706f
C5 Vp m1_831_275# 0.215f
C6 m1_559_n458# m1_831_275# 0.0183f
C7 Vp Vin 0.176f
C8 m1_559_n458# Vin 0.181f
C9 m1_831_275# Vn 0.232f
C10 V13 m1_831_275# 0.184f
C11 m1_559_n458# Vp 0.0628f
C12 Vin Vn 0.347f
C13 Vin V13 0.0076f
C14 m1_831_275# 0 1.05f
C15 Vin 0 1.79f
C16 V13 0 0.365f
C17 Vn 0 0.117f
C18 Vp 0 3.98f
C19 m1_559_n458# 0 0.286f
.ends

.subckt sky130_fd_pr__nfet_01v8_DD6SHA a_n33_n130# a_15_n42# a_n175_n182# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n33_n130# a_n73_n42# 0.0209f
C1 a_n33_n130# a_15_n42# 0.0209f
C2 a_15_n42# a_n73_n42# 0.0699f
C3 a_15_n42# a_n175_n182# 0.0637f
C4 a_n73_n42# a_n175_n182# 0.0716f
C5 a_n33_n130# a_n175_n182# 0.314f
.ends

.subckt sky130_fd_pr__pfet_01v8_7DPLFP w_n245_n261# a_n107_n42# a_n49_n139# a_49_n42#
+ VSUBS
X0 a_49_n42# a_n49_n139# a_n107_n42# w_n245_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.49
C0 a_49_n42# a_n107_n42# 0.0396f
C1 w_n245_n261# a_n49_n139# 0.221f
C2 w_n245_n261# a_n107_n42# 0.0224f
C3 a_49_n42# w_n245_n261# 0.0224f
C4 a_n107_n42# a_n49_n139# 0.00895f
C5 a_49_n42# a_n49_n139# 0.00895f
C6 a_49_n42# VSUBS 0.0487f
C7 a_n107_n42# VSUBS 0.0487f
C8 a_n49_n139# VSUBS 0.206f
C9 w_n245_n261# VSUBS 0.876f
.ends

.subckt sky130_fd_pr__pfet_01v8_MDPZBH a_n102_n42# a_44_n42# a_n44_n139# w_n240_n261#
+ VSUBS
X0 a_44_n42# a_n44_n139# a_n102_n42# w_n240_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.44
C0 a_44_n42# a_n102_n42# 0.0423f
C1 w_n240_n261# a_n44_n139# 0.208f
C2 w_n240_n261# a_n102_n42# 0.0224f
C3 a_44_n42# w_n240_n261# 0.0224f
C4 a_n102_n42# a_n44_n139# 0.00823f
C5 a_44_n42# a_n44_n139# 0.00823f
C6 a_44_n42# VSUBS 0.0485f
C7 a_n102_n42# VSUBS 0.0485f
C8 a_n44_n139# VSUBS 0.191f
C9 w_n240_n261# VSUBS 0.858f
.ends

.subckt th06 Vp Vin V06 m1_904_n796# Vn
XXM0 Vin m1_904_n796# Vn Vn sky130_fd_pr__nfet_01v8_DD6SHA
XXM1 Vp Vp Vin m1_904_n796# Vn sky130_fd_pr__pfet_01v8_7DPLFP
XXM2 Vp V06 m1_904_n796# Vp Vn sky130_fd_pr__pfet_01v8_MDPZBH
XXM3 Vn m1_904_n796# V06 Vn sky130_fd_pr__nfet_01v8_MYA4RC
C0 Vn Vin 0.0188f
C1 Vp V06 0.06f
C2 Vn V06 0.00141f
C3 Vp Vn 0.0214f
C4 m1_904_n796# Vin 0.203f
C5 m1_904_n796# V06 0.157f
C6 Vp m1_904_n796# 0.197f
C7 Vp Vin 0.113f
C8 Vn m1_904_n796# 0.0382f
C9 Vp 0 1.69f
C10 m1_904_n796# 0 0.495f
C11 V06 0 0.217f
C12 Vn 0 0.286f
C13 Vin 0 0.524f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGAKDL a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
+ VSUBS
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n73_n200# a_n33_n297# 0.0293f
C1 w_n211_n419# a_n33_n297# 0.191f
C2 a_n73_n200# a_15_n200# 0.321f
C3 w_n211_n419# a_15_n200# 0.0336f
C4 a_15_n200# a_n33_n297# 0.0293f
C5 w_n211_n419# a_n73_n200# 0.0336f
C6 a_15_n200# VSUBS 0.164f
C7 a_n73_n200# VSUBS 0.164f
C8 a_n33_n297# VSUBS 0.147f
C9 w_n211_n419# VSUBS 1.14f
.ends

.subckt sky130_fd_pr__nfet_01v8_4X3CDA a_n306_n216# a_n180_n130# a_n238_n42# a_180_n42#
X0 a_180_n42# a_n180_n130# a_n238_n42# a_n306_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.8
C0 a_180_n42# a_n238_n42# 0.0147f
C1 a_n180_n130# a_n238_n42# 0.0189f
C2 a_n180_n130# a_180_n42# 0.0189f
C3 a_180_n42# a_n306_n216# 0.075f
C4 a_n238_n42# a_n306_n216# 0.075f
C5 a_n180_n130# a_n306_n216# 1.1f
.ends

.subckt sky130_fd_pr__pfet_01v8_MWB9BZ a_15_n43# w_n211_n262# a_n73_n43# a_n33_n140#
+ VSUBS
X0 a_15_n43# a_n33_n140# a_n73_n43# w_n211_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.15
C0 a_n73_n43# a_n33_n140# 0.0193f
C1 w_n211_n262# a_n33_n140# 0.187f
C2 a_n73_n43# a_15_n43# 0.0715f
C3 w_n211_n262# a_15_n43# 0.0198f
C4 a_15_n43# a_n33_n140# 0.0193f
C5 w_n211_n262# a_n73_n43# 0.0198f
C6 a_15_n43# VSUBS 0.0453f
C7 a_n73_n43# VSUBS 0.0453f
C8 a_n33_n140# VSUBS 0.143f
C9 w_n211_n262# VSUBS 0.752f
.ends

.subckt sky130_fd_pr__nfet_01v8_L9ESAD a_n175_n190# a_n73_n50# a_n33_n138# a_15_n50#
X0 a_15_n50# a_n33_n138# a_n73_n50# a_n175_n190# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_15_n50# a_n73_n50# 0.0826f
C1 a_n33_n138# a_n73_n50# 0.0216f
C2 a_n33_n138# a_15_n50# 0.0216f
C3 a_15_n50# a_n175_n190# 0.0704f
C4 a_n73_n50# a_n175_n190# 0.0797f
C5 a_n33_n138# a_n175_n190# 0.315f
.ends

.subckt th11 V11 Vin Vp m1_705_187# Vn m1_577_n654#
XXM0 Vn Vp Vn m1_577_n654# Vn sky130_fd_pr__pfet_01v8_XGAKDL
XXM1 Vn Vin m1_577_n654# m1_705_187# sky130_fd_pr__nfet_01v8_4X3CDA
XXM2 m1_705_187# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_MWB9BZ
XXM3 V11 Vp m1_705_187# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM4 Vn Vn m1_705_187# V11 sky130_fd_pr__nfet_01v8_L9ESAD
C0 Vp m1_705_187# 0.286f
C1 Vn Vp 0.0775f
C2 m1_577_n654# V11 5.55e-19
C3 Vn m1_705_187# 0.463f
C4 Vp Vin 0.285f
C5 Vin m1_705_187# 0.0649f
C6 Vn Vin 0.135f
C7 Vp m1_577_n654# 0.0405f
C8 m1_577_n654# m1_705_187# 0.0258f
C9 Vn m1_577_n654# 0.0457f
C10 m1_577_n654# Vin 0.213f
C11 Vp V11 0.026f
C12 m1_705_187# V11 0.377f
C13 Vn V11 0.00287f
C14 Vin V11 2.69e-19
C15 Vin 0 1.27f
C16 m1_705_187# 0 0.602f
C17 V11 0 0.346f
C18 Vn 0 0.355f
C19 Vp 0 2.61f
C20 m1_577_n654# 0 0.286f
.ends

.subckt sky130_fd_pr__nfet_01v8_42G4RD a_n80_n42# a_n148_n216# a_n33_n130# a_22_n42#
X0 a_22_n42# a_n33_n130# a_n80_n42# a_n148_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_n33_n130# a_22_n42# 0.00866f
C1 a_n33_n130# a_n80_n42# 0.00866f
C2 a_n80_n42# a_22_n42# 0.0604f
C3 a_22_n42# a_n148_n216# 0.0698f
C4 a_n80_n42# a_n148_n216# 0.0698f
C5 a_n33_n130# a_n148_n216# 0.321f
.ends

.subckt sky130_fd_pr__pfet_01v8_DDPLQ8 a_n77_n42# w_n215_n261# a_n33_n139# a_19_n42#
+ VSUBS
X0 a_19_n42# a_n33_n139# a_n77_n42# w_n215_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 w_n215_n261# a_n77_n42# 0.017f
C1 w_n215_n261# a_n33_n139# 0.181f
C2 a_n33_n139# a_n77_n42# 0.0127f
C3 w_n215_n261# a_19_n42# 0.0399f
C4 a_19_n42# a_n77_n42# 0.0641f
C5 a_19_n42# a_n33_n139# 0.0127f
C6 a_19_n42# VSUBS 0.035f
C7 a_n77_n42# VSUBS 0.05f
C8 a_n33_n139# VSUBS 0.149f
C9 w_n215_n261# VSUBS 0.797f
.ends

.subckt sky130_fd_pr__nfet_01v8_VWP3K3 a_n33_n130# a_15_n42# a_n141_182# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n141_182# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n33_n130# a_15_n42# 0.0209f
C1 a_n33_n130# a_n73_n42# 0.0209f
C2 a_n73_n42# a_15_n42# 0.0699f
C3 a_15_n42# a_n141_182# 0.0643f
C4 a_n73_n42# a_n141_182# 0.0643f
C5 a_n33_n130# a_n141_182# 0.317f
.ends

.subckt sky130_fd_pr__pfet_01v8_LZD9A4 a_n80_n42# a_22_n42# a_n33_n139# w_n218_n261#
+ VSUBS
X0 a_22_n42# a_n33_n139# a_n80_n42# w_n218_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 w_n218_n261# a_n80_n42# 0.0222f
C1 w_n218_n261# a_n33_n139# 0.185f
C2 a_n33_n139# a_n80_n42# 0.0084f
C3 w_n218_n261# a_22_n42# 0.0222f
C4 a_22_n42# a_n80_n42# 0.0604f
C5 a_22_n42# a_n33_n139# 0.0084f
C6 a_22_n42# VSUBS 0.0474f
C7 a_n80_n42# VSUBS 0.0474f
C8 a_n33_n139# VSUBS 0.149f
C9 w_n218_n261# VSUBS 0.775f
.ends

.subckt sky130_fd_pr__nfet_01v8_VRD6K3 a_n77_n42# a_n145_n214# a_n33_n130# a_19_n42#
X0 a_19_n42# a_n33_n130# a_n77_n42# a_n145_n214# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_n33_n130# a_19_n42# 0.0136f
C1 a_n33_n130# a_n77_n42# 0.0136f
C2 a_n77_n42# a_19_n42# 0.0641f
C3 a_19_n42# a_n145_n214# 0.0677f
C4 a_n77_n42# a_n145_n214# 0.0677f
C5 a_n33_n130# a_n145_n214# 0.32f
.ends

.subckt th04 V04 Vn Vp m1_892_n998# m1_620_n488# Vin
XXM0 m1_892_n998# Vn Vin Vn sky130_fd_pr__nfet_01v8_42G4RD
XXM1 m1_620_n488# Vp Vin m1_892_n998# Vn sky130_fd_pr__pfet_01v8_DDPLQ8
XXM2 Vp m1_620_n488# Vn Vp sky130_fd_pr__nfet_01v8_VWP3K3
XXM3 Vp V04 m1_892_n998# Vp Vn sky130_fd_pr__pfet_01v8_LZD9A4
XXM4 Vn Vn m1_892_n998# V04 sky130_fd_pr__nfet_01v8_VRD6K3
C0 Vin V04 0.00141f
C1 V04 Vn 0.0639f
C2 m1_892_n998# m1_620_n488# 0.0117f
C3 Vp V04 0.0462f
C4 Vin Vn 0.0468f
C5 m1_620_n488# V04 0.00264f
C6 Vin Vp 0.14f
C7 Vp Vn 0.0386f
C8 m1_892_n998# V04 0.13f
C9 Vin m1_620_n488# 0.0346f
C10 m1_620_n488# Vn 2.16e-19
C11 m1_892_n998# Vin 0.463f
C12 m1_892_n998# Vn 0.1f
C13 m1_620_n488# Vp 0.17f
C14 m1_892_n998# Vp 0.383f
C15 m1_892_n998# 0 0.832f
C16 V04 0 0.287f
C17 Vn 0 0.259f
C18 Vp 0 2.13f
C19 m1_620_n488# 0 0.0632f
C20 Vin 0 0.679f
.ends

.subckt adc1 VGND VPWR b[0] b[1] b[2] b[3] p[0] p[10] p[11] p[12] p[13] p[14] p[1]
+ p[2] p[3] p[4] p[5] p[6] p[7] p[8] p[9] Vin
X_49_ net7 _02_ _19_ _20_ _21_ VGND VGND VPWR VPWR net17 _49_/a_208_47# _49_/a_75_199#
+ _49_/a_544_297# _49_/a_315_47# _49_/a_201_297# sky130_fd_sc_hd__a311o_1
X_48_ net11 _02_ _07_ VGND VGND VPWR VPWR _21_ _48_/a_181_47# _48_/a_109_47# _48_/a_27_47#
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ net5 _12_ _17_ VGND VGND VPWR VPWR _20_ _47_/a_384_47# _47_/a_81_21# _47_/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xth02_0 th15_0/Vin p[1] th02_0/m1_983_133# VPWR th02_0/m1_571_144# VGND th02
X_46_ _04_ VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__inv_2
X_29_ net11 net13 net12 VGND VGND VPWR VPWR _03_ _29_/a_29_53# _29_/a_183_297# _29_/a_111_297#
+ sky130_fd_sc_hd__or3_1
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28_ _00_ _01_ VGND VGND VPWR VPWR _02_ _28_/a_109_297# sky130_fd_sc_hd__nor2_1
X_45_ _02_ _09_ _12_ _13_ _18_ VGND VGND VPWR VPWR net16 _45_/a_193_297# _45_/a_465_47#
+ _45_/a_205_47# _45_/a_109_297# _45_/a_27_47# sky130_fd_sc_hd__a221o_1
X_44_ net14 _14_ _15_ _17_ net2 VGND VGND VPWR VPWR _18_ _44_/a_256_47# _44_/a_584_47#
+ _44_/a_93_21# _44_/a_250_297# _44_/a_346_47# sky130_fd_sc_hd__a32o_1
X_27_ net14 net15 net3 net2 VGND VGND VPWR VPWR _01_ _27_/a_277_297# _27_/a_205_297#
+ _27_/a_27_297# _27_/a_109_297# sky130_fd_sc_hd__or4_1
XFILLER_0_7_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_43_ _00_ _06_ _10_ _16_ VGND VGND VPWR VPWR _17_ _43_/a_369_47# _43_/a_469_47# _43_/a_297_47#
+ _43_/a_193_413# _43_/a_27_47# sky130_fd_sc_hd__and4b_1
X_26_ net5 net4 net6 VGND VGND VPWR VPWR _00_ _26_/a_29_53# _26_/a_183_297# _26_/a_111_297#
+ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_42_ net3 net15 net14 VGND VGND VPWR VPWR _16_ _42_/a_109_93# _42_/a_368_53# _42_/a_209_311#
+ _42_/a_296_53# sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_3_Left_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND VPWR VPWR b[0] output16/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_41_ _06_ _10_ VGND VGND VPWR VPWR _15_ _41_/a_145_75# _41_/a_59_75# sky130_fd_sc_hd__and2_1
Xoutput17 net17 VGND VGND VPWR VPWR b[1] output17/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_40_ net15 net3 net2 _00_ VGND VGND VPWR VPWR _14_ _40_/a_297_297# _40_/a_191_297#
+ _40_/a_109_297# sky130_fd_sc_hd__nor4_1
Xoutput18 net18 VGND VGND VPWR VPWR b[2] output18/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xth09_0 p[8] Vin VGND th09_0/m1_485_n505# VPWR th09_0/m1_962_372# th09
XPHY_EDGE_ROW_0_Left_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR b[3] output19/a_27_47# sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xth14_0 p[13] th15_0/Vin VGND th14_0/m1_641_n318# VPWR th14_0/m1_891_419# th14
Xinput1 p[0] VGND VGND VPWR VPWR net1 input1/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xth07_0 VPWR Vin p[6] th07_0/m1_808_n892# VGND th07
Xinput2 p[10] VGND VGND VPWR VPWR net2 input2/a_27_47# sky130_fd_sc_hd__buf_1
Xinput3 p[11] VGND VGND VPWR VPWR net3 input3/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xth12_0 p[11] Vin th12_0/m1_394_n856# th12_0/m1_529_n42# VPWR VGND th12
Xinput4 p[12] VGND VGND VPWR VPWR net4 input4/a_75_212# sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xth05_0 VPWR p[4] Vin th05_0/m1_752_n794# VGND th05
Xinput5 p[13] VGND VGND VPWR VPWR net5 input5/a_664_47# input5/a_841_47# input5/a_381_47#
+ input5/a_62_47# input5/a_558_47# sky130_fd_sc_hd__dlymetal6s2s_1
Xinput6 p[14] VGND VGND VPWR VPWR net6 input6/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_1_Left_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xth10_0 p[9] Vin th10_0/m1_502_n495# th10_0/m1_536_174# VGND VPWR th10
Xinput7 p[1] VGND VGND VPWR VPWR net7 input7/a_27_47# sky130_fd_sc_hd__buf_1
Xinput10 p[4] VGND VGND VPWR VPWR net10 input10/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xth03_0 p[2] Vin VPWR th03_0/m1_890_n844# th03_0/m1_638_n591# VGND th03
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 p[2] VGND VGND VPWR VPWR net8 input8/a_27_47# sky130_fd_sc_hd__buf_1
Xinput11 p[5] VGND VGND VPWR VPWR net11 input11/a_27_47# sky130_fd_sc_hd__buf_1
X_39_ net5 net6 VGND VGND VPWR VPWR _13_ _39_/a_129_47# _39_/a_47_47# _39_/a_285_47#
+ _39_/a_377_297# sky130_fd_sc_hd__xnor2_1
Xinput9 p[3] VGND VGND VPWR VPWR net9 input9/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput12 p[6] VGND VGND VPWR VPWR net12 input12/a_27_47# sky130_fd_sc_hd__buf_1
X_55_ _14_ _15_ _20_ _22_ VGND VGND VPWR VPWR net19 _55_/a_472_297# _55_/a_80_21#
+ _55_/a_300_47# _55_/a_217_297# sky130_fd_sc_hd__a211o_1
X_38_ net4 _06_ _10_ _11_ VGND VGND VPWR VPWR _12_ _38_/a_109_47# _38_/a_197_47# _38_/a_303_47#
+ _38_/a_27_47# sky130_fd_sc_hd__and4_1
X_54_ _25_ VGND VGND VPWR VPWR net18 _54_/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput13 p[7] VGND VGND VPWR VPWR net13 input13/a_27_47# sky130_fd_sc_hd__buf_1
X_37_ net14 net15 net3 net2 VGND VGND VPWR VPWR _11_ _37_/a_109_47# _37_/a_197_47#
+ _37_/a_303_47# _37_/a_27_47# sky130_fd_sc_hd__and4_1
Xth01_0 p[0] VGND th01_0/m1_991_n1219# th01_0/m1_571_n501# VPWR th15_0/Vin th01
Xinput14 p[8] VGND VGND VPWR VPWR net14 input14/a_27_47# sky130_fd_sc_hd__buf_1
X_53_ _21_ _22_ _24_ VGND VGND VPWR VPWR _25_ _53_/a_29_53# _53_/a_183_297# _53_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_36_ net11 net10 net13 net12 VGND VGND VPWR VPWR _10_ _36_/a_109_47# _36_/a_197_47#
+ _36_/a_303_47# _36_/a_27_47# sky130_fd_sc_hd__and4_1
X_52_ _02_ _06_ _23_ _12_ net5 VGND VGND VPWR VPWR _24_ _52_/a_256_47# _52_/a_584_47#
+ _52_/a_93_21# _52_/a_250_297# _52_/a_346_47# sky130_fd_sc_hd__a32o_1
Xinput15 p[9] VGND VGND VPWR VPWR net15 input15/a_27_47# sky130_fd_sc_hd__buf_1
X_35_ _04_ _05_ _07_ _08_ VGND VGND VPWR VPWR _09_ _35_/a_489_413# _35_/a_226_47#
+ _35_/a_556_47# _35_/a_226_297# _35_/a_76_199# sky130_fd_sc_hd__a2bb2o_1
X_51_ _03_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__inv_2
X_34_ net11 net12 VGND VGND VPWR VPWR _08_ _34_/a_129_47# _34_/a_47_47# _34_/a_285_47#
+ _34_/a_377_297# sky130_fd_sc_hd__xnor2_1
X_33_ net13 _06_ net10 VGND VGND VPWR VPWR _07_ _33_/a_109_93# _33_/a_368_53# _33_/a_209_311#
+ _33_/a_296_53# sky130_fd_sc_hd__and3b_1
X_50_ net5 net6 _15_ _11_ VGND VGND VPWR VPWR _22_ _50_/a_515_93# _50_/a_223_47# _50_/a_615_93#
+ _50_/a_343_93# _50_/a_429_93# _50_/a_27_47# sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpreamp_0 Vin th15_0/Vin VGND VPWR preamp
X_32_ net7 net1 net9 net8 VGND VGND VPWR VPWR _06_ _32_/a_109_47# _32_/a_197_47# _32_/a_303_47#
+ _32_/a_27_47# sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_5_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31_ net7 net8 VGND VGND VPWR VPWR _05_ _31_/a_117_297# _31_/a_285_297# _31_/a_285_47#
+ _31_/a_35_297# sky130_fd_sc_hd__xor2_1
Xth15_0 p[14] th15_0/Vin th15_0/m1_597_n912# th15_0/m1_849_n157# VPWR VGND th15
X_30_ net9 net10 _03_ net1 VGND VGND VPWR VPWR _04_ _30_/a_465_297# _30_/a_297_297#
+ _30_/a_215_297# _30_/a_392_297# _30_/a_109_53# sky130_fd_sc_hd__or4b_1
Xth08_0 VPWR Vin p[7] th08_0/m1_477_n803# VGND th08
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xth13_0 p[12] Vin th13_0/m1_831_275# VGND th13_0/m1_559_n458# VPWR th13
XFILLER_0_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xth06_0 VPWR Vin p[5] th06_0/m1_904_n796# VGND th06
XFILLER_0_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xth11_0 p[10] Vin VPWR th11_0/m1_705_187# VGND th11_0/m1_577_n654# th11
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xth04_0 p[3] VGND VPWR th04_0/m1_892_n998# th04_0/m1_620_n488# Vin th04
C0 input9/a_75_212# net13 4.4e-19
C1 _13_ _50_/a_343_93# 5.63e-20
C2 _08_ _33_/a_209_311# 0.0122f
C3 _10_ p[14] 0.00247f
C4 _18_ p[14] 2.75e-20
C5 b[1] p[2] 0.00184f
C6 th13_0/m1_559_n458# output16/a_27_47# 1.24e-20
C7 _09_ _38_/a_27_47# 0.00195f
C8 _49_/a_201_297# VGND -0.00403f
C9 _12_ input4/a_75_212# 2.09e-20
C10 net2 p[1] 7.54e-20
C11 VPWR _36_/a_303_47# -4.83e-19
C12 _26_/a_29_53# net11 1.08e-20
C13 _05_ _52_/a_93_21# 1.12e-20
C14 p[7] b[1] 0.00476f
C15 _00_ _21_ 9.26e-20
C16 net15 net8 0.2f
C17 net15 net3 0.394f
C18 b[1] _30_/a_109_53# 0.00655f
C19 net11 _48_/a_109_47# 1.74e-19
C20 b[1] th02_0/m1_983_133# 7.26e-20
C21 _11_ net12 3.82e-21
C22 th14_0/m1_641_n318# th12_0/m1_529_n42# 0.00311f
C23 net4 _39_/a_377_297# 8.88e-19
C24 net10 p[3] 0.00113f
C25 _09_ _52_/a_93_21# 0.0227f
C26 _43_/a_193_413# _22_ 0.00133f
C27 _43_/a_369_47# _14_ 0.00135f
C28 net7 input5/a_381_47# 4.91e-19
C29 p[3] _10_ 1.37e-20
C30 net3 _29_/a_29_53# 1.68e-20
C31 net8 _06_ 0.00282f
C32 net3 _06_ 0.0072f
C33 _44_/a_250_297# th15_0/Vin 7.01e-19
C34 net4 _45_/a_27_47# 0.024f
C35 input2/a_27_47# p[1] 0.012f
C36 _19_ b[1] 0.00967f
C37 net10 net13 0.375f
C38 _35_/a_226_47# _29_/a_29_53# 2.64e-19
C39 th06_0/m1_904_n796# VGND 0.0173f
C40 th14_0/m1_641_n318# VGND 0.00635f
C41 _10_ net13 0.00151f
C42 _30_/a_392_297# net12 2.19e-20
C43 _31_/a_285_297# _05_ 6.12e-19
C44 _29_/a_29_53# _07_ 1.19e-20
C45 p[0] input5/a_62_47# 1.39e-19
C46 output19/a_27_47# net6 0.00112f
C47 _35_/a_226_47# _06_ 0.00487f
C48 VGND input5/a_664_47# 0.0136f
C49 _05_ th04_0/m1_892_n998# 5.09e-21
C50 _18_ net13 1.06e-20
C51 _06_ _07_ 0.185f
C52 th15_0/Vin _42_/a_368_53# 1.2e-20
C53 th15_0/m1_849_n157# _11_ 7.84e-20
C54 _47_/a_81_21# _15_ 0.00332f
C55 _31_/a_35_297# net5 2.04e-21
C56 _24_ b[1] 2.68e-19
C57 _33_/a_368_53# net12 2.63e-19
C58 th03_0/m1_638_n591# p[1] 0.135f
C59 th11_0/m1_705_187# p[0] 1.49e-19
C60 p[5] th06_0/m1_904_n796# 0.114f
C61 Vin input13/a_27_47# 0.00534f
C62 _40_/a_109_297# th15_0/Vin 7.23e-19
C63 _35_/a_76_199# net5 3.38e-19
C64 _44_/a_584_47# net14 7.2e-19
C65 _05_ input8/a_27_47# 1.58e-19
C66 VPWR _37_/a_109_47# -4.38e-19
C67 input10/a_27_47# input12/a_27_47# 0.0154f
C68 th01_0/m1_571_n501# VGND 8.66e-21
C69 _15_ _22_ 0.0236f
C70 input14/a_27_47# b[3] 0.00268f
C71 _35_/a_489_413# _09_ 0.0296f
C72 _35_/a_556_47# _08_ 7.71e-19
C73 net2 net7 0.00234f
C74 _20_ _36_/a_27_47# 0.00148f
C75 input15/a_27_47# net6 0.146f
C76 input14/a_27_47# th12_0/m1_529_n42# 7.48e-19
C77 net10 _34_/a_377_297# 1.62e-19
C78 _39_/a_129_47# b[0] 2.6e-20
C79 _52_/a_250_297# _23_ 3.17e-19
C80 _13_ _22_ 0.00309f
C81 VGND net18 0.255f
C82 _53_/a_29_53# _25_ 0.00146f
C83 th05_0/m1_752_n794# p[4] 0.00599f
C84 _44_/a_93_21# _44_/a_250_297# -6.97e-22
C85 _03_ net17 5.1e-19
C86 p[10] th15_0/Vin 0.185f
C87 input14/a_27_47# VGND 0.0389f
C88 input2/a_27_47# net7 0.00213f
C89 b[1] _34_/a_129_47# 3.51e-19
C90 p[5] net18 1.98e-19
C91 net2 net6 0.00139f
C92 _04_ _36_/a_109_47# 2.39e-19
C93 input10/a_27_47# VGND 0.00285f
C94 net1 output17/a_27_47# 8.12e-19
C95 th13_0/m1_831_275# th15_0/m1_849_n157# 5.99e-19
C96 _20_ net15 0.0021f
C97 _02_ _52_/a_256_47# 0.00344f
C98 _04_ _52_/a_584_47# 2.5e-19
C99 _03_ _49_/a_75_199# 0.0849f
C100 net17 _14_ 2.4e-20
C101 Vin th09_0/m1_485_n505# 0.134f
C102 _26_/a_29_53# net6 0.0032f
C103 _04_ _27_/a_277_297# 0.00113f
C104 th03_0/m1_638_n591# net7 3.67e-20
C105 _00_ net7 8.12e-21
C106 p[3] _33_/a_209_311# 9.2e-21
C107 net4 _24_ 8.65e-20
C108 _45_/a_193_297# _35_/a_226_47# 8.15e-21
C109 VPWR _54_/a_75_212# 0.0475f
C110 _29_/a_111_297# _09_ 5.79e-20
C111 _20_ _29_/a_29_53# 0.0111f
C112 p[5] input10/a_27_47# 0.0193f
C113 p[6] input13/a_27_47# 1.07e-19
C114 _14_ _49_/a_75_199# 6.79e-20
C115 _20_ _06_ 0.133f
C116 net1 input5/a_841_47# 1.33e-19
C117 output19/a_27_47# _10_ 2.79e-20
C118 _01_ p[2] 0.00164f
C119 Vin net19 1.54e-19
C120 _31_/a_35_297# VGND -0.00828f
C121 _33_/a_209_311# net13 0.0227f
C122 _45_/a_27_47# _21_ 1.18e-20
C123 _45_/a_205_47# net5 8.28e-20
C124 _17_ _39_/a_47_47# 1.47e-20
C125 Vin input1/a_75_212# 0.01f
C126 _21_ _23_ 0.0217f
C127 _17_ _40_/a_191_297# 4.35e-19
C128 _35_/a_76_199# VGND -0.0034f
C129 _19_ _27_/a_27_297# 0.082f
C130 _53_/a_29_53# _06_ 0.0709f
C131 VPWR _30_/a_465_297# -4.57e-19
C132 _00_ net6 0.00178f
C133 input3/a_27_47# input5/a_62_47# 0.00179f
C134 _12_ th15_0/Vin 0.00101f
C135 input15/a_27_47# _10_ 4.5e-19
C136 _12_ _52_/a_346_47# 3.8e-19
C137 _24_ _52_/a_250_297# 3.03e-19
C138 input15/a_27_47# _18_ 8.27e-21
C139 net5 _41_/a_59_75# 2.41e-19
C140 _44_/a_250_297# _04_ 5.57e-21
C141 p[13] th15_0/Vin 0.0887f
C142 VGND net5 1.2f
C143 net11 _45_/a_27_47# 3.64e-20
C144 _37_/a_27_47# input5/a_841_47# 4.64e-20
C145 _06_ _50_/a_343_93# 0.0376f
C146 net6 output16/a_27_47# 1.5e-19
C147 _19_ _01_ 0.031f
C148 net11 _23_ 0.0461f
C149 _26_/a_183_297# _22_ 0.00184f
C150 _02_ _42_/a_209_311# 9.92e-19
C151 Vin b[1] 0.376f
C152 _21_ _30_/a_109_53# 3.31e-20
C153 net10 net2 2.05e-20
C154 _00_ _55_/a_80_21# 5.5e-19
C155 _03_ net9 0.149f
C156 net2 _10_ 3.15e-19
C157 p[14] _42_/a_209_311# 5.85e-22
C158 _17_ _02_ 0.00482f
C159 net5 _50_/a_223_47# 0.00202f
C160 _18_ net2 0.00181f
C161 _26_/a_29_53# net10 3.48e-22
C162 _00_ _47_/a_384_47# 5.15e-20
C163 _26_/a_29_53# _10_ 0.0265f
C164 _25_ _22_ 5.39e-19
C165 _17_ p[14] 1.07e-19
C166 _05_ input13/a_27_47# 3.93e-19
C167 _26_/a_29_53# _18_ 5.26e-20
C168 _43_/a_469_47# net15 7.41e-19
C169 _43_/a_193_413# net14 1.11e-19
C170 _43_/a_27_47# _01_ 9.77e-20
C171 net3 input6/a_27_47# 2.52e-19
C172 _13_ _38_/a_27_47# 4.58e-19
C173 output18/a_27_47# output16/a_27_47# 7.85e-19
C174 VPWR _08_ -0.0171f
C175 p[2] p[1] 0.0489f
C176 _36_/a_27_47# _22_ 2.82e-20
C177 p[7] net11 4.23e-20
C178 VGND input12/a_27_47# 0.0407f
C179 net10 input2/a_27_47# 1.17e-20
C180 _19_ _42_/a_109_93# 1.14e-21
C181 _09_ input13/a_27_47# 1.27e-21
C182 VPWR _44_/a_256_47# -7.56e-19
C183 _24_ _21_ 0.0388f
C184 VGND b[3] 0.148f
C185 _45_/a_205_47# VGND -2.47e-19
C186 _37_/a_27_47# _11_ 0.0018f
C187 _04_ p[10] 8.48e-21
C188 _13_ _52_/a_93_21# 1.31e-19
C189 p[5] input12/a_27_47# 0.00359f
C190 th02_0/m1_983_133# p[1] 0.122f
C191 VGND th12_0/m1_529_n42# 0.00796f
C192 net15 _47_/a_81_21# 0.00106f
C193 _03_ net8 0.0287f
C194 _03_ net3 4.27e-20
C195 _31_/a_117_297# _03_ 5.32e-19
C196 VPWR input7/a_27_47# 0.0772f
C197 _00_ _10_ 0.301f
C198 _00_ _18_ 0.157f
C199 b[1] p[6] 0.00562f
C200 _04_ _49_/a_544_297# 0.00204f
C201 _19_ net11 6.27e-21
C202 Vin p[8] 0.564f
C203 VPWR _39_/a_47_47# 0.0668f
C204 net14 p[9] 1.05e-19
C205 input3/a_27_47# net3 0.03f
C206 net4 Vin 4.16e-19
C207 net3 _14_ 0.0295f
C208 net14 _15_ 0.225f
C209 _35_/a_226_47# _03_ 0.028f
C210 net8 _14_ 4.23e-19
C211 net15 _22_ 2.74e-19
C212 VGND _41_/a_59_75# 0.0205f
C213 VPWR _40_/a_191_297# -6.82e-19
C214 _47_/a_81_21# _06_ 0.0388f
C215 _03_ _07_ 0.0113f
C216 _13_ b[0] 0.00299f
C217 net16 output16/a_27_47# 0.0101f
C218 _02_ _30_/a_215_297# 3.58e-21
C219 _53_/a_111_297# _22_ 4.7e-20
C220 Vin _33_/a_109_93# 1.63e-19
C221 _19_ p[1] 3.92e-20
C222 p[6] _48_/a_27_47# 8.49e-19
C223 th14_0/m1_891_419# p[11] 0.0117f
C224 _39_/a_377_297# net6 0.00143f
C225 _22_ _29_/a_29_53# 2.24e-21
C226 _02_ _38_/a_109_47# 1.63e-19
C227 _22_ _06_ 0.124f
C228 VPWR _49_/a_208_47# -5.93e-19
C229 _40_/a_297_297# net6 7.47e-22
C230 _12_ net12 7.94e-21
C231 p[5] VGND 0.283f
C232 _43_/a_193_413# _16_ 0.0261f
C233 p[2] net7 0.00157f
C234 _39_/a_47_47# p[12] 0.00138f
C235 VGND _50_/a_223_47# 0.0159f
C236 VPWR th11_0/m1_577_n654# -4.9e-19
C237 _45_/a_27_47# net6 0.021f
C238 _23_ net6 2.13e-19
C239 th11_0/m1_705_187# th01_0/m1_571_n501# 0.00336f
C240 VGND _53_/a_183_297# -4.34e-19
C241 Vin _27_/a_27_297# 2.8e-19
C242 net2 p[11] 0.00681f
C243 _04_ _12_ 1.42e-19
C244 _31_/a_35_297# net17 0.0514f
C245 net9 input5/a_664_47# 5.29e-19
C246 p[3] _30_/a_215_297# 5.18e-19
C247 VPWR _02_ 0.332f
C248 th15_0/Vin _37_/a_109_47# 5.47e-20
C249 _50_/a_27_47# _50_/a_343_93# -7.11e-33
C250 _49_/a_201_297# net8 7.3e-19
C251 _12_ th15_0/m1_849_n157# 2.47e-21
C252 p[13] _04_ 0.00111f
C253 net11 _34_/a_129_47# 0.00242f
C254 VPWR p[14] 0.0553f
C255 _31_/a_35_297# _49_/a_75_199# 6.24e-19
C256 _30_/a_215_297# net13 0.0246f
C257 _12_ _38_/a_197_47# 0.00173f
C258 Vin th13_0/m1_559_n458# 2.77e-19
C259 _15_ _16_ 0.0607f
C260 _19_ net7 0.0458f
C261 _34_/a_47_47# net12 0.0385f
C262 _35_/a_226_47# _49_/a_201_297# 1.66e-20
C263 Vin _01_ 5.85e-20
C264 _31_/a_285_47# Vin 2.61e-20
C265 VPWR _32_/a_109_47# 0.00124f
C266 _27_/a_109_297# net2 7.24e-20
C267 _05_ b[1] 0.0316f
C268 _44_/a_346_47# _10_ 9.13e-21
C269 _39_/a_47_47# input4/a_75_212# 3.1e-19
C270 _02_ p[12] 8.05e-19
C271 _43_/a_369_47# VGND -8.43e-19
C272 _25_ _38_/a_27_47# 5.76e-19
C273 _03_ _20_ 0.0794f
C274 net17 net5 4.21e-21
C275 _09_ b[1] 0.00408f
C276 _02_ b[2] 2.81e-19
C277 p[12] p[14] 2.26e-19
C278 p[2] input9/a_75_212# 5.13e-20
C279 th14_0/m1_641_n318# net3 3.58e-19
C280 net8 input5/a_664_47# 0.0116f
C281 _48_/a_181_47# p[6] 8.16e-20
C282 _04_ _34_/a_47_47# 1.17e-20
C283 VPWR p[3] 0.114f
C284 _17_ output19/a_27_47# 0.00122f
C285 _45_/a_193_297# _22_ 0.0234f
C286 input5/a_381_47# _42_/a_209_311# 3.88e-19
C287 net3 input5/a_664_47# 0.00215f
C288 _20_ _14_ 0.144f
C289 _43_/a_27_47# net7 6.31e-19
C290 input5/a_558_47# net5 0.0597f
C291 _10_ _39_/a_377_297# 7.42e-19
C292 _02_ _55_/a_217_297# 6.01e-19
C293 _36_/a_303_47# net12 1.37e-19
C294 p[7] input9/a_75_212# 0.00102f
C295 _31_/a_35_297# th11_0/m1_705_187# 9e-21
C296 _09_ _48_/a_27_47# 0.00541f
C297 net16 _45_/a_27_47# 8.68e-19
C298 VPWR net13 0.599f
C299 th14_0/m1_891_419# _42_/a_209_311# 6.86e-21
C300 _45_/a_27_47# _10_ 0.0143f
C301 _24_ net6 0.00121f
C302 net10 _23_ 0.00216f
C303 _45_/a_27_47# _18_ 0.00347f
C304 _17_ input15/a_27_47# 6.14e-19
C305 _10_ _23_ 0.00192f
C306 p[10] net1 0.00387f
C307 p[10] output17/a_27_47# 0.12f
C308 _43_/a_27_47# net6 9.07e-20
C309 input5/a_62_47# net5 0.00329f
C310 _17_ _37_/a_197_47# 9.19e-21
C311 net11 Vin 0.00253f
C312 _49_/a_544_297# net1 0.00175f
C313 net2 _42_/a_209_311# 5.1e-19
C314 _03_ th03_0/m1_890_n844# 3.64e-21
C315 _38_/a_27_47# _06_ 0.0172f
C316 _22_ _50_/a_27_47# 0.0276f
C317 _14_ _50_/a_343_93# 9.76e-19
C318 _15_ _50_/a_429_93# 6.82e-19
C319 b[1] input11/a_27_47# 0.00688f
C320 net3 input14/a_27_47# 9.36e-19
C321 _05_ _33_/a_109_93# 0.0206f
C322 VPWR _34_/a_377_297# -0.00192f
C323 Vin p[1] 0.18f
C324 _20_ _49_/a_201_297# 5.24e-21
C325 _17_ net2 0.181f
C326 VPWR th10_0/m1_536_174# 0.0406f
C327 net4 _09_ 0.00262f
C328 p[7] net10 6e-19
C329 net10 _30_/a_109_53# 5.6e-20
C330 _09_ _33_/a_109_93# 7.36e-20
C331 _40_/a_109_297# _11_ 0.00522f
C332 p[6] _21_ 0.00219f
C333 _43_/a_27_47# _55_/a_80_21# 1.56e-19
C334 _52_/a_93_21# _06_ 0.0584f
C335 net17 VGND 0.212f
C336 input2/a_27_47# _42_/a_209_311# 1e-22
C337 net9 net5 0.0368f
C338 _05_ _52_/a_250_297# 8.86e-22
C339 VGND _49_/a_75_199# 5.87e-20
C340 net15 net14 1.07f
C341 b[1] _30_/a_297_297# 3.14e-19
C342 _31_/a_35_297# net8 0.0408f
C343 VGND input5/a_558_47# -0.00104f
C344 _09_ _52_/a_250_297# 1.97e-20
C345 input10/a_27_47# p[4] 0.0217f
C346 net16 _24_ 6.93e-19
C347 _43_/a_193_413# net19 3.31e-19
C348 _43_/a_469_47# _14_ 0.00259f
C349 p[13] output17/a_27_47# 0.00118f
C350 p[13] net1 2.13e-19
C351 net14 _29_/a_29_53# 1.61e-20
C352 VPWR output19/a_27_47# 0.0245f
C353 net11 p[6] 0.0135f
C354 net14 _06_ 1.94e-19
C355 _17_ _00_ 0.0851f
C356 _32_/a_27_47# b[1] 6.39e-19
C357 _24_ _10_ 0.00484f
C358 _31_/a_285_297# _06_ 1.01e-20
C359 _44_/a_256_47# th15_0/Vin 1.36e-19
C360 net4 _45_/a_109_297# 6.43e-20
C361 VPWR input5/a_381_47# 8.33e-19
C362 Vin net7 0.00646f
C363 th09_0/m1_485_n505# p[9] 0.0164f
C364 _35_/a_76_199# _35_/a_226_47# -2.84e-32
C365 _05_ _01_ 5.03e-19
C366 _35_/a_76_199# _07_ 0.00226f
C367 _35_/a_489_413# _06_ 9.22e-19
C368 VGND input5/a_62_47# 0.0499f
C369 p[13] input5/a_841_47# 7.34e-19
C370 _31_/a_285_47# _05_ 5.61e-19
C371 _43_/a_27_47# _10_ 0.0279f
C372 th15_0/Vin input7/a_27_47# 2.79e-19
C373 net8 net5 0.48f
C374 net3 net5 0.0365f
C375 _43_/a_27_47# _18_ 0.0201f
C376 _47_/a_81_21# _14_ 6.24e-20
C377 _47_/a_299_297# _15_ 0.0103f
C378 _03_ _22_ 2.55e-20
C379 _09_ _01_ 4.69e-21
C380 VPWR input15/a_27_47# 0.0113f
C381 VPWR th14_0/m1_891_419# 0.049f
C382 th11_0/m1_705_187# VGND 0.01f
C383 _39_/a_47_47# th15_0/Vin 8.52e-22
C384 _40_/a_191_297# th15_0/Vin 3.41e-19
C385 input3/a_27_47# _22_ 5.13e-20
C386 net19 p[9] 0.0767f
C387 _15_ net19 0.166f
C388 _14_ _22_ 0.00449f
C389 VPWR _37_/a_197_47# -3.27e-19
C390 _49_/a_315_47# b[1] 5.66e-19
C391 _35_/a_226_297# _09_ 4.98e-19
C392 input2/a_27_47# _30_/a_215_297# 3.51e-20
C393 Vin net6 6.97e-19
C394 _45_/a_193_297# _52_/a_93_21# 6.01e-19
C395 _30_/a_465_297# net12 8.01e-20
C396 _05_ _21_ 0.0104f
C397 th15_0/m1_597_n912# p[14] 4.12e-21
C398 net10 _34_/a_129_47# 0.003f
C399 _39_/a_285_47# b[0] 1.88e-19
C400 net15 _16_ 0.214f
C401 _52_/a_256_47# _23_ 6.66e-19
C402 p[7] _33_/a_209_311# 7.23e-19
C403 input15/a_27_47# p[12] 3.73e-19
C404 VPWR net2 0.958f
C405 _53_/a_29_53# net18 0.0118f
C406 _09_ _21_ 0.263f
C407 VGND net9 0.372f
C408 _12_ _11_ 0.195f
C409 _44_/a_93_21# _44_/a_256_47# -6.6e-20
C410 th15_0/Vin th11_0/m1_577_n654# 0.00967f
C411 _29_/a_111_297# _06_ 6.74e-20
C412 _26_/a_29_53# VPWR 0.0356f
C413 _16_ _06_ 0.00162f
C414 b[1] _34_/a_285_47# 0.00368f
C415 th12_0/m1_394_n856# th09_0/m1_485_n505# 4.53e-19
C416 _38_/a_27_47# _50_/a_27_47# 2.37e-20
C417 Vin input9/a_75_212# 0.00188f
C418 net3 b[3] 2.43e-20
C419 _02_ _52_/a_346_47# 0.00526f
C420 net11 _05_ 2.76e-19
C421 _31_/a_35_297# _20_ 1.69e-19
C422 _02_ th15_0/Vin 7.82e-21
C423 net9 _50_/a_223_47# 2e-19
C424 net3 th12_0/m1_529_n42# 3.65e-21
C425 b[1] _15_ 1.19e-19
C426 _26_/a_111_297# net6 1.12e-19
C427 VPWR input2/a_27_47# 0.00832f
C428 _44_/a_346_47# _17_ 7.2e-19
C429 _34_/a_285_47# _48_/a_27_47# 6.66e-20
C430 th15_0/Vin p[14] 0.356f
C431 _49_/a_201_297# _22_ 2.45e-20
C432 net11 _09_ 0.0262f
C433 _29_/a_183_297# _03_ 7.36e-19
C434 _35_/a_76_199# _20_ 3.21e-20
C435 input12/a_27_47# p[4] 9.06e-19
C436 th08_0/m1_477_n803# input12/a_27_47# 1.64e-20
C437 th03_0/m1_638_n591# th01_0/m1_991_n1219# 2.42e-20
C438 VPWR th03_0/m1_638_n591# 0.0124f
C439 net8 VGND 0.405f
C440 net3 VGND 0.323f
C441 VPWR _00_ 0.416f
C442 _08_ net12 0.0269f
C443 input15/a_27_47# input4/a_75_212# 1.1e-21
C444 _31_/a_117_297# VGND -0.00177f
C445 _33_/a_296_53# net13 3.71e-20
C446 _20_ net5 0.0651f
C447 _35_/a_226_47# VGND -0.0111f
C448 _19_ _27_/a_109_297# 7.54e-21
C449 net16 Vin 3.38e-19
C450 VGND _07_ 0.195f
C451 net10 Vin 0.00328f
C452 _04_ _08_ 5.99e-19
C453 VPWR output16/a_27_47# 0.123f
C454 _17_ _45_/a_27_47# 1.16e-20
C455 Vin _10_ 0.00189f
C456 p[7] _35_/a_556_47# 4.37e-20
C457 Vin _18_ 3.79e-21
C458 _32_/a_27_47# _01_ 0.0266f
C459 net17 _49_/a_75_199# 0.00127f
C460 VGND p[4] 0.35f
C461 _31_/a_35_297# th03_0/m1_890_n844# 4.56e-19
C462 net11 _45_/a_109_297# 7.46e-20
C463 th08_0/m1_477_n803# VGND 0.00633f
C464 p[8] p[9] 0.11f
C465 _06_ _50_/a_429_93# 0.00169f
C466 net17 input5/a_558_47# 2.88e-21
C467 _44_/a_93_21# p[14] 2.07e-19
C468 net4 _15_ 0.00427f
C469 net11 input11/a_27_47# 0.00318f
C470 _05_ net7 0.0129f
C471 p[5] th08_0/m1_477_n803# 2.39e-19
C472 p[5] p[4] 0.254f
C473 input13/a_27_47# _06_ 4.89e-19
C474 net4 _13_ 0.212f
C475 net5 _50_/a_343_93# 0.00124f
C476 _09_ net7 0.00258f
C477 _32_/a_27_47# _21_ 8.95e-19
C478 _26_/a_111_297# _10_ 7.13e-20
C479 _03_ _52_/a_93_21# 0.00985f
C480 net18 _22_ 1.68e-19
C481 _43_/a_193_413# _01_ 8.16e-19
C482 _43_/a_297_47# net14 1.09e-21
C483 _49_/a_315_47# _01_ 1.82e-19
C484 net14 input6/a_27_47# 7.05e-19
C485 Vin th02_0/m1_571_144# 8.17e-20
C486 th11_0/m1_705_187# net17 1.25e-19
C487 th15_0/Vin th10_0/m1_536_174# 0.0771f
C488 net10 p[6] 0.0081f
C489 _02_ net12 2.28e-19
C490 VPWR _44_/a_346_47# -8.74e-19
C491 _27_/a_27_297# _15_ 9.85e-20
C492 _04_ th11_0/m1_577_n654# 4.01e-19
C493 _20_ _41_/a_59_75# 1.78e-20
C494 p[13] _44_/a_250_297# 4.09e-20
C495 _45_/a_465_47# VGND -8.14e-19
C496 _09_ net6 5.43e-20
C497 _17_ _19_ 8.82e-21
C498 _32_/a_197_47# _02_ 3.78e-19
C499 _20_ VGND 0.471f
C500 _13_ _52_/a_250_297# 5.43e-19
C501 th12_0/m1_394_n856# p[8] 0.00768f
C502 net15 _47_/a_299_297# 1.44e-20
C503 _03_ net14 1.5e-19
C504 _31_/a_285_297# _03_ 0.00677f
C505 _04_ _02_ 0.0541f
C506 input3/a_27_47# net14 3.47e-19
C507 b[1] _25_ 0.0015f
C508 _05_ input9/a_75_212# 1.24e-21
C509 net17 net9 1.26e-20
C510 _35_/a_489_413# _03_ 0.0205f
C511 _47_/a_299_297# _06_ 0.0174f
C512 net15 net19 0.0501f
C513 _01_ _15_ 0.007f
C514 net14 _14_ 0.184f
C515 VGND _41_/a_145_75# 4.11e-19
C516 VPWR _40_/a_297_297# -5.42e-19
C517 Vin _33_/a_209_311# 2.54e-19
C518 _20_ _50_/a_223_47# 1.71e-19
C519 VGND _53_/a_29_53# -0.0168f
C520 _43_/a_27_47# _17_ 0.00131f
C521 b[1] _36_/a_27_47# 7.95e-19
C522 output19/a_27_47# th15_0/Vin 0.0163f
C523 Vin p[11] 0.00572f
C524 VPWR _45_/a_27_47# -0.00418f
C525 net9 _49_/a_75_199# 0.00382f
C526 th15_0/m1_849_n157# p[14] 0.0846f
C527 p[3] net12 0.00564f
C528 _39_/a_129_47# net6 6.91e-19
C529 _35_/a_76_199# _22_ 6.58e-21
C530 net9 input5/a_558_47# 4.42e-19
C531 net19 _06_ 0.00522f
C532 VPWR _23_ -0.00374f
C533 _47_/a_81_21# net5 4.59e-19
C534 th15_0/Vin input5/a_381_47# 3.39e-19
C535 _21_ _34_/a_285_47# 6.94e-20
C536 _50_/a_343_93# _41_/a_59_75# 6.13e-22
C537 _39_/a_377_297# p[12] 4.68e-19
C538 _45_/a_109_297# net6 7.82e-19
C539 VGND _50_/a_343_93# -3.89e-19
C540 net13 net12 0.363f
C541 _21_ _15_ 1.13e-21
C542 _11_ _54_/a_75_212# 3.22e-20
C543 _22_ net5 0.405f
C544 _04_ p[3] 0.00437f
C545 input15/a_27_47# th15_0/Vin 0.00696f
C546 th14_0/m1_891_419# th15_0/Vin 0.0726f
C547 _15_ _42_/a_109_93# 0.00367f
C548 p[13] p[10] 0.00616f
C549 th03_0/m1_890_n844# VGND 0.0241f
C550 VPWR p[2] 0.248f
C551 Vin _27_/a_109_297# 5.3e-20
C552 _45_/a_27_47# p[12] 2.9e-19
C553 net17 net8 0.18f
C554 net3 net17 3.72e-19
C555 net15 b[1] 0.00314f
C556 _31_/a_117_297# net17 0.00149f
C557 net9 input5/a_62_47# 3.12e-19
C558 _13_ _21_ 1.69e-19
C559 th15_0/Vin _37_/a_197_47# 1.87e-19
C560 _05_ net10 0.457f
C561 _05_ _10_ 9.25e-21
C562 _29_/a_111_297# _03_ 7.48e-19
C563 net14 _49_/a_201_297# 1.52e-19
C564 VPWR p[7] 0.0867f
C565 _04_ net13 0.569f
C566 net16 _09_ 0.00707f
C567 net8 _49_/a_75_199# 0.00214f
C568 VPWR _30_/a_109_53# 9.49e-19
C569 b[1] _29_/a_29_53# 0.0026f
C570 net3 _49_/a_75_199# 2.01e-19
C571 _23_ b[2] 2.87e-20
C572 _32_/a_27_47# net7 0.00559f
C573 th01_0/m1_991_n1219# th02_0/m1_983_133# 4.16e-19
C574 VPWR th02_0/m1_983_133# 0.0376f
C575 _09_ net10 0.037f
C576 net8 input5/a_558_47# 0.00357f
C577 net3 input5/a_558_47# 0.0137f
C578 b[1] _06_ 0.0885f
C579 _44_/a_93_21# output19/a_27_47# 7.25e-20
C580 _09_ _10_ 0.0222f
C581 _12_ _38_/a_303_47# 0.00153f
C582 _14_ _16_ 0.0584f
C583 net2 th15_0/Vin 0.0484f
C584 _34_/a_377_297# net12 0.00251f
C585 _09_ _18_ 7.01e-21
C586 _35_/a_226_47# _49_/a_75_199# 8.73e-20
C587 net1 input7/a_27_47# 0.0383f
C588 net4 _36_/a_27_47# 0.0103f
C589 _44_/a_584_47# _10_ 1.14e-20
C590 _49_/a_75_199# _07_ 4.05e-21
C591 _49_/a_201_297# input8/a_27_47# 2.46e-21
C592 _48_/a_27_47# _06_ 0.0251f
C593 net18 _38_/a_27_47# 0.00997f
C594 _13_ net11 2.34e-19
C595 b[1] th05_0/m1_752_n794# 0.0202f
C596 VPWR _19_ 0.0335f
C597 th14_0/m1_641_n318# net14 0.00168f
C598 _45_/a_27_47# input4/a_75_212# 2.18e-20
C599 net8 input5/a_62_47# 2.05e-19
C600 net14 input5/a_664_47# 0.0179f
C601 net3 input5/a_62_47# 0.00164f
C602 _04_ _34_/a_377_297# 1.7e-20
C603 _49_/a_315_47# net7 0.00706f
C604 _43_/a_193_413# net7 3.49e-19
C605 VPWR _24_ 0.0129f
C606 _47_/a_81_21# _41_/a_59_75# 1.5e-19
C607 _10_ _39_/a_129_47# 2.51e-19
C608 _02_ _55_/a_472_297# 1.25e-19
C609 th11_0/m1_705_187# net8 0.00167f
C610 _52_/a_93_21# net18 8.21e-21
C611 _47_/a_81_21# VGND -0.0112f
C612 net16 _45_/a_109_297# 5.1e-20
C613 p[8] net15 1.73e-20
C614 net4 net15 8.68e-19
C615 _43_/a_27_47# VPWR 0.0186f
C616 th03_0/m1_638_n591# th15_0/Vin 2.04e-19
C617 _45_/a_109_297# _10_ 0.00202f
C618 _00_ th15_0/Vin 1.03e-19
C619 net4 _53_/a_111_297# 2.09e-19
C620 _22_ _41_/a_59_75# 6.24e-22
C621 _17_ Vin 3.65e-19
C622 VGND _22_ 0.0404f
C623 p[2] th04_0/m1_620_n488# 6.98e-20
C624 _44_/a_93_21# net2 0.0273f
C625 input1/a_75_212# p[0] 0.0197f
C626 net4 _06_ 0.281f
C627 _43_/a_193_413# net6 2.41e-20
C628 _17_ _37_/a_303_47# 1.23e-20
C629 _33_/a_109_93# _06_ 6.96e-19
C630 _02_ net1 0.00251f
C631 net8 net9 0.0605f
C632 net3 net9 5.09e-20
C633 p[7] th04_0/m1_620_n488# 1.62e-21
C634 _24_ b[2] 1.85e-19
C635 _20_ net17 4e-20
C636 _15_ net7 8.4e-20
C637 th04_0/m1_620_n488# th02_0/m1_983_133# 2.13e-21
C638 _22_ _50_/a_223_47# 0.031f
C639 _15_ _50_/a_515_93# 0.00147f
C640 VPWR _34_/a_129_47# -9.47e-19
C641 net14 input14/a_27_47# 0.0232f
C642 _05_ _33_/a_209_311# 0.0311f
C643 _35_/a_226_47# net9 1.22e-20
C644 net9 _07_ 1.39e-20
C645 _53_/a_183_297# _22_ 3.71e-20
C646 _02_ input5/a_841_47# 0.00591f
C647 _20_ _49_/a_75_199# 0.0233f
C648 _27_/a_27_297# net15 0.00888f
C649 VPWR th07_0/m1_808_n892# 0.0188f
C650 _39_/a_47_47# _11_ 3.9e-19
C651 th14_0/m1_641_n318# _16_ 2.77e-20
C652 net10 _30_/a_297_297# 1.68e-19
C653 _08_ _33_/a_368_53# 5.04e-19
C654 _09_ _33_/a_209_311# 3.79e-20
C655 _48_/a_181_47# _06_ 6.4e-19
C656 _10_ _30_/a_297_297# 1.25e-20
C657 _40_/a_191_297# _11_ 0.00207f
C658 _38_/a_27_47# net5 1.76e-19
C659 _43_/a_193_413# _55_/a_80_21# 2.54e-19
C660 _43_/a_27_47# _55_/a_217_297# 2.18e-19
C661 _35_/a_76_199# _52_/a_93_21# 6.83e-21
C662 b[1] p[0] 0.00454f
C663 _52_/a_250_297# _06_ 0.0058f
C664 _21_ _25_ 0.00164f
C665 p[9] net6 0.139f
C666 _44_/a_93_21# _00_ 4.54e-20
C667 _15_ net6 0.17f
C668 net10 _32_/a_27_47# 2.76e-20
C669 _32_/a_27_47# _10_ 0.00217f
C670 _21_ _36_/a_27_47# 0.0276f
C671 p[3] net1 6.54e-19
C672 Vin _30_/a_215_297# 1.01e-19
C673 net3 net8 9.23e-19
C674 _32_/a_27_47# _18_ 1.18e-20
C675 net15 _01_ 0.0314f
C676 _31_/a_117_297# net8 5.91e-19
C677 _36_/a_197_47# net13 1.06e-19
C678 _52_/a_93_21# net5 0.0124f
C679 _13_ net6 0.0106f
C680 net4 _39_/a_285_47# 9.71e-19
C681 _26_/a_29_53# net12 6.55e-19
C682 p[14] _37_/a_27_47# 3.97e-19
C683 _29_/a_183_297# VGND 4.41e-19
C684 net19 input6/a_27_47# 0.00574f
C685 _01_ _29_/a_29_53# 8.33e-20
C686 net1 net13 3.51e-19
C687 _01_ _06_ 0.00157f
C688 VPWR th09_0/m1_962_372# 0.00391f
C689 _04_ net2 0.158f
C690 _44_/a_346_47# th15_0/Vin 1.88e-19
C691 net11 _25_ 0.0262f
C692 net4 _45_/a_193_297# 7.41e-19
C693 net5 b[0] 3.39e-19
C694 _31_/a_35_297# input8/a_27_47# 0.00955f
C695 _02_ _11_ 0.0621f
C696 _55_/a_80_21# _15_ 0.107f
C697 net11 _36_/a_27_47# 0.0717f
C698 _35_/a_226_47# _07_ 8.96e-19
C699 _35_/a_226_297# _06_ 1.28e-19
C700 _26_/a_29_53# _04_ 2.3e-21
C701 th03_0/m1_890_n844# _49_/a_75_199# 1.69e-21
C702 _43_/a_193_413# _10_ 0.0174f
C703 _43_/a_193_413# _18_ 0.0413f
C704 net14 net5 0.0263f
C705 p[14] _11_ 4.99e-20
C706 _53_/a_111_297# _21_ 4.38e-19
C707 _47_/a_384_47# _15_ 0.00112f
C708 net15 _42_/a_109_93# 4.62e-19
C709 Vin th01_0/m1_991_n1219# 0.0178f
C710 VPWR Vin 2.7f
C711 _21_ _29_/a_29_53# 0.0775f
C712 _04_ input2/a_27_47# 4.5e-21
C713 _21_ _06_ 0.143f
C714 _40_/a_297_297# th15_0/Vin 1.26e-19
C715 _20_ net9 0.328f
C716 input3/a_27_47# net19 0.00105f
C717 VPWR _37_/a_303_47# -3.13e-19
C718 _14_ net19 0.00714f
C719 _42_/a_109_93# _06_ 5.53e-20
C720 _35_/a_556_47# _09_ 0.00122f
C721 net10 _34_/a_285_47# 0.0454f
C722 VGND _38_/a_27_47# 0.00767f
C723 _04_ _00_ 1.98e-20
C724 Vin p[12] 0.0619f
C725 _10_ p[9] 0.00225f
C726 net4 _50_/a_27_47# 0.0239f
C727 _44_/a_93_21# _44_/a_346_47# -5.12e-20
C728 _10_ _15_ 0.479f
C729 net15 p[1] 1.8e-19
C730 net11 _29_/a_29_53# 0.00514f
C731 _18_ _15_ 0.042f
C732 _13_ net16 0.0198f
C733 net11 _06_ 0.546f
C734 _03_ b[1] 0.0738f
C735 _26_/a_111_297# VPWR -5.92e-20
C736 _13_ net10 4.52e-21
C737 _52_/a_93_21# VGND -0.0175f
C738 p[2] th15_0/Vin 1.51e-21
C739 _13_ _10_ 0.0621f
C740 net14 b[3] 8.65e-19
C741 input3/a_27_47# b[1] 2.97e-19
C742 _13_ _18_ 0.019f
C743 _20_ net8 5.07e-19
C744 th13_0/m1_831_275# p[14] 4.94e-20
C745 _20_ net3 4.07e-19
C746 _02_ _52_/a_584_47# 0.00389f
C747 b[1] _14_ 1.1e-19
C748 net9 _50_/a_343_93# 6.64e-19
C749 net14 th12_0/m1_529_n42# 3.01e-19
C750 VPWR p[6] 0.136f
C751 net11 th05_0/m1_752_n794# 1.09e-19
C752 net5 _16_ 1.99e-20
C753 th15_0/Vin th02_0/m1_983_133# 0.0143f
C754 VGND b[0] 0.181f
C755 _35_/a_226_47# _20_ 5.19e-20
C756 _20_ _07_ 1.28e-21
C757 _22_ _49_/a_75_199# 9.85e-21
C758 _30_/a_392_297# net13 6.64e-20
C759 net1 input5/a_381_47# 1.27e-19
C760 input5/a_381_47# output17/a_27_47# 6.6e-20
C761 net14 VGND 0.441f
C762 _31_/a_285_297# VGND -0.00136f
C763 th04_0/m1_892_n998# VGND 0.0189f
C764 _33_/a_368_53# net13 2.1e-20
C765 Vin th04_0/m1_620_n488# 0.00167f
C766 _17_ _39_/a_129_47# 1.38e-20
C767 _43_/a_193_413# p[11] 8.34e-20
C768 _35_/a_489_413# VGND -8.78e-19
C769 _36_/a_27_47# net6 5.1e-19
C770 net15 net7 2.91e-19
C771 _05_ _30_/a_215_297# 0.0453f
C772 net8 _50_/a_343_93# 7.25e-19
C773 net14 _50_/a_223_47# 5.89e-21
C774 th14_0/m1_641_n318# net19 1.17e-19
C775 _17_ _45_/a_109_297# 4.29e-22
C776 input8/a_27_47# VGND 0.0574f
C777 net19 input5/a_664_47# 1.38e-21
C778 th14_0/m1_891_419# input5/a_841_47# 3.61e-21
C779 _36_/a_109_47# net13 0.00126f
C780 _49_/a_201_297# b[1] 0.0025f
C781 net7 _29_/a_29_53# 6.01e-19
C782 p[10] input7/a_27_47# 1.82e-19
C783 net8 th03_0/m1_890_n844# 3.83e-19
C784 _03_ _33_/a_109_93# 2.78e-19
C785 net7 _06_ 0.00447f
C786 input3/a_27_47# p[8] 6.2e-19
C787 net1 net2 1.64e-19
C788 _43_/a_27_47# th15_0/Vin 1.9e-19
C789 _06_ _50_/a_515_93# 0.00244f
C790 net2 output17/a_27_47# 0.0285f
C791 output18/a_27_47# _25_ 0.072f
C792 _44_/a_250_297# p[14] 7.34e-21
C793 net4 _14_ 1.54e-20
C794 net15 net6 0.0664f
C795 _28_/a_109_297# _15_ 0.00346f
C796 _47_/a_81_21# net9 3.49e-19
C797 p[9] p[11] 0.00354f
C798 input15/a_27_47# _37_/a_27_47# 3.27e-19
C799 _21_ _50_/a_27_47# 3.38e-21
C800 _23_ net12 2.28e-21
C801 _15_ p[11] 0.00591f
C802 VPWR _05_ 0.118f
C803 _29_/a_29_53# net6 1.4e-20
C804 _26_/a_183_297# _10_ 5.74e-19
C805 th06_0/m1_904_n796# b[1] 4.33e-20
C806 VGND _16_ -0.00582f
C807 _29_/a_111_297# VGND -1.9e-19
C808 net6 _06_ 0.308f
C809 input2/a_27_47# output17/a_27_47# 0.107f
C810 net9 _22_ 0.0023f
C811 net1 input2/a_27_47# 4.81e-19
C812 b[1] input5/a_664_47# 0.00195f
C813 _43_/a_369_47# net14 6.79e-21
C814 _03_ _27_/a_27_297# 2.68e-19
C815 th08_0/m1_477_n803# th03_0/m1_890_n844# 2.96e-20
C816 p[10] th11_0/m1_577_n654# 4.13e-19
C817 VPWR _09_ 0.297f
C818 p[0] p[1] 0.0399f
C819 input14/a_27_47# net19 3.63e-19
C820 net16 _25_ 1.16e-19
C821 input15/a_27_47# _11_ 4.4e-19
C822 net2 _37_/a_27_47# 0.0692f
C823 VPWR _44_/a_584_47# -2.28e-19
C824 _00_ net1 9.43e-19
C825 net15 _55_/a_80_21# 0.00759f
C826 _27_/a_27_297# _14_ 1.66e-21
C827 net10 _25_ 2.66e-19
C828 net11 _50_/a_27_47# 6.05e-21
C829 _10_ _25_ 0.0109f
C830 p[7] net12 0.0406f
C831 _30_/a_109_53# net12 4.25e-20
C832 input9/a_75_212# _29_/a_29_53# 9.7e-21
C833 _47_/a_81_21# net8 2.08e-21
C834 net3 _47_/a_81_21# 6.66e-19
C835 net10 _36_/a_27_47# 0.0366f
C836 _03_ _01_ 2.85e-19
C837 _31_/a_285_47# _03_ 8.54e-19
C838 _10_ _36_/a_27_47# 0.00109f
C839 _04_ p[2] 2.84e-20
C840 output18/a_27_47# _06_ 0.0114f
C841 _55_/a_80_21# _06_ 5.15e-19
C842 _18_ _36_/a_27_47# 5.46e-20
C843 _12_ _39_/a_47_47# 0.0317f
C844 Vin th15_0/m1_597_n912# 7.85e-19
C845 VPWR _39_/a_129_47# -9.47e-19
C846 b[1] net18 0.00134f
C847 net2 _11_ 0.234f
C848 th12_0/m1_394_n856# p[11] 9.12e-21
C849 _35_/a_226_297# _03_ 0.00101f
C850 net8 _22_ 3.3e-20
C851 _01_ _14_ 0.0193f
C852 net3 _22_ 9.39e-20
C853 _09_ b[2] 4.28e-20
C854 _04_ _30_/a_109_53# 9.19e-21
C855 _20_ _50_/a_343_93# 0.00826f
C856 _08_ _34_/a_47_47# 0.00123f
C857 _43_/a_193_413# _17_ 0.0503f
C858 _26_/a_29_53# _11_ 1.09e-19
C859 VPWR _45_/a_109_297# -0.011f
C860 _39_/a_285_47# net6 1.53e-19
C861 _30_/a_215_297# _30_/a_297_297# -8.88e-34
C862 _35_/a_226_47# _22_ 1.39e-20
C863 _20_ th03_0/m1_890_n844# 3.1e-19
C864 _22_ _07_ 1.19e-20
C865 _03_ _21_ 0.0818f
C866 b[1] input10/a_27_47# 0.00691f
C867 _00_ _37_/a_27_47# 6.15e-20
C868 VPWR input11/a_27_47# 0.0378f
C869 _47_/a_299_297# net5 0.00198f
C870 net15 _10_ 0.0101f
C871 _29_/a_183_297# net9 3.51e-19
C872 p[0] net7 1.36e-19
C873 _39_/a_129_47# p[12] 2.4e-20
C874 _53_/a_111_297# _10_ 2.06e-19
C875 _18_ net15 0.0382f
C876 _45_/a_193_297# net6 9.84e-20
C877 VGND _50_/a_429_93# 4.71e-19
C878 _19_ _04_ 0.356f
C879 net16 _06_ 0.0511f
C880 net10 _29_/a_29_53# 1.77e-19
C881 p[13] th11_0/m1_577_n654# 0.029f
C882 input3/a_27_47# _42_/a_109_93# 0.00249f
C883 p[9] _42_/a_209_311# 5.51e-21
C884 net10 _06_ 0.184f
C885 _10_ _29_/a_29_53# 5.17e-19
C886 Vin th15_0/Vin 0.999f
C887 net19 net5 0.00124f
C888 _10_ _06_ 1.14f
C889 _15_ _42_/a_209_311# 0.0521f
C890 _14_ _42_/a_109_93# 0.00141f
C891 Vin _27_/a_205_297# 2.93e-20
C892 _45_/a_109_297# p[12] 5.61e-21
C893 _12_ _02_ 0.265f
C894 _18_ _06_ 0.54f
C895 net14 net17 5.43e-19
C896 _31_/a_35_297# b[1] 0.0176f
C897 _00_ _11_ 0.238f
C898 VGND input13/a_27_47# 0.0473f
C899 th15_0/Vin _37_/a_303_47# 1.45e-19
C900 _17_ p[9] 1.03e-20
C901 p[13] _02_ 2.99e-19
C902 _17_ _15_ 0.0752f
C903 net11 _03_ 0.0952f
C904 _49_/a_544_297# net13 3.43e-19
C905 _01_ _49_/a_201_297# 0.0105f
C906 net10 th05_0/m1_752_n794# 6.61e-20
C907 net14 _49_/a_75_199# 3.67e-19
C908 VPWR _30_/a_297_297# -5.22e-19
C909 _35_/a_76_199# b[1] 0.00458f
C910 net14 input5/a_558_47# 0.0325f
C911 p[5] input13/a_27_47# 3.09e-19
C912 _27_/a_27_297# input5/a_664_47# 0.0116f
C913 _44_/a_250_297# output19/a_27_47# 6.42e-20
C914 _29_/a_183_297# net3 7.38e-21
C915 th09_0/m1_485_n505# b[3] 2.57e-19
C916 p[8] input14/a_27_47# 0.0132f
C917 VPWR _32_/a_27_47# 0.0395f
C918 th09_0/m1_485_n505# th12_0/m1_529_n42# 0.0107f
C919 _26_/a_29_53# _52_/a_584_47# 7.45e-20
C920 _20_ _47_/a_81_21# 0.0457f
C921 net6 _50_/a_27_47# 0.0428f
C922 b[1] net5 0.00349f
C923 input8/a_27_47# _49_/a_75_199# 1.99e-20
C924 _02_ _34_/a_47_47# 1.09e-19
C925 net16 _39_/a_285_47# 1.29e-19
C926 net14 input5/a_62_47# 5.28e-20
C927 net19 b[3] 0.0546f
C928 _44_/a_93_21# Vin 2.93e-21
C929 _20_ _22_ 0.183f
C930 net19 th12_0/m1_529_n42# 4.2e-21
C931 _47_/a_299_297# _41_/a_59_75# 0.00146f
C932 th09_0/m1_485_n505# VGND 0.00241f
C933 _10_ _39_/a_285_47# 0.00289f
C934 _02_ _55_/a_300_47# 0.00371f
C935 _12_ net13 0.00632f
C936 _47_/a_299_297# VGND -3.63e-19
C937 net16 _45_/a_193_297# 0.00187f
C938 _43_/a_193_413# VPWR 0.0063f
C939 VPWR _49_/a_315_47# 3.4e-19
C940 net19 _41_/a_59_75# 1.97e-20
C941 _45_/a_193_297# _10_ 0.0047f
C942 VGND net19 0.151f
C943 _53_/a_29_53# _22_ 0.00749f
C944 net11 _49_/a_201_297# 1.42e-19
C945 _44_/a_250_297# net2 0.0188f
C946 _21_ input5/a_664_47# 9.42e-22
C947 net15 p[11] 1.71e-19
C948 _03_ net7 0.078f
C949 b[1] input12/a_27_47# 0.00658f
C950 th13_0/m1_831_275# output16/a_27_47# 7.67e-22
C951 _47_/a_81_21# _50_/a_343_93# 0.00282f
C952 _47_/a_299_297# _50_/a_223_47# 2.74e-20
C953 input1/a_75_212# VGND 0.0586f
C954 net1 p[2] 0.0277f
C955 _43_/a_297_47# net6 8.23e-22
C956 th14_0/m1_641_n318# _42_/a_109_93# 1.75e-19
C957 _35_/a_76_199# _33_/a_109_93# 3.08e-19
C958 net6 input6/a_27_47# 0.00208f
C959 _33_/a_209_311# _06_ 0.0187f
C960 net14 net9 7.12e-20
C961 th04_0/m1_892_n998# net9 5.18e-21
C962 p[7] net1 7.5e-20
C963 _14_ net7 0.00251f
C964 _22_ _50_/a_343_93# 0.0597f
C965 _15_ _50_/a_615_93# 0.00183f
C966 net1 _30_/a_109_53# 0.0297f
C967 VPWR _34_/a_285_47# -0.00233f
C968 _05_ _33_/a_296_53# 4.53e-19
C969 net1 th02_0/m1_983_133# 4.09e-19
C970 th02_0/m1_983_133# output17/a_27_47# 0.00138f
C971 Vin net12 0.00543f
C972 net4 net5 0.0447f
C973 _34_/a_47_47# net13 1.68e-19
C974 VPWR p[9] 0.429f
C975 _40_/a_109_297# net2 0.0011f
C976 VPWR _15_ 0.912f
C977 net16 _50_/a_27_47# 2.35e-20
C978 _03_ net6 2.9e-20
C979 _39_/a_377_297# _11_ 2.57e-20
C980 p[10] th14_0/m1_891_419# 5.19e-20
C981 input8/a_27_47# net9 3.71e-20
C982 _40_/a_297_297# _11_ 9.94e-19
C983 net10 _50_/a_27_47# 3.78e-21
C984 _35_/a_226_47# _52_/a_93_21# 4.89e-20
C985 _35_/a_76_199# _52_/a_250_297# 3.4e-21
C986 b[1] VGND 0.56f
C987 _10_ _50_/a_27_47# 0.0154f
C988 _21_ net18 0.00215f
C989 _52_/a_256_47# _06_ 0.00207f
C990 _19_ output17/a_27_47# 7.69e-19
C991 input5/a_664_47# p[1] 1.21e-20
C992 VPWR _13_ 0.0804f
C993 _04_ Vin 0.00428f
C994 _18_ _50_/a_27_47# 0.0665f
C995 _44_/a_250_297# _00_ 6.39e-20
C996 _19_ net1 2.86e-19
C997 _45_/a_27_47# _11_ 0.0703f
C998 _14_ net6 2.11e-19
C999 _23_ _11_ 2e-20
C1000 Vin th15_0/m1_849_n157# 0.0502f
C1001 net3 net14 0.689f
C1002 net14 net8 0.0516f
C1003 p[5] b[1] 0.00883f
C1004 _31_/a_285_297# net8 0.0215f
C1005 p[12] p[9] 1.02e-19
C1006 VGND _48_/a_27_47# 0.0548f
C1007 _36_/a_303_47# net13 5.5e-20
C1008 _31_/a_35_297# _01_ 4.27e-19
C1009 p[12] _15_ 0.00116f
C1010 _52_/a_250_297# net5 0.018f
C1011 p[10] net2 0.0373f
C1012 _03_ input9/a_75_212# 9.32e-20
C1013 _27_/a_27_297# net5 3.48e-19
C1014 p[0] th02_0/m1_571_144# 0.0179f
C1015 _49_/a_201_297# net7 0.00419f
C1016 _35_/a_76_199# _01_ 3.08e-21
C1017 _13_ p[12] 8.72e-19
C1018 net11 net18 0.00221f
C1019 _44_/a_584_47# th15_0/Vin 2.71e-19
C1020 p[8] b[3] 0.0392f
C1021 _29_/a_111_297# net9 8.06e-21
C1022 net8 input8/a_27_47# 0.0181f
C1023 p[8] th12_0/m1_529_n42# 0.00973f
C1024 _55_/a_80_21# _14_ 0.0175f
C1025 _55_/a_217_297# _15_ 0.0474f
C1026 p[6] net12 0.0309f
C1027 VPWR th12_0/m1_394_n856# 0.00333f
C1028 p[13] input5/a_381_47# 0.00464f
C1029 _35_/a_489_413# _07_ 0.00429f
C1030 _43_/a_297_47# _10_ 0.00118f
C1031 p[10] input2/a_27_47# 0.0095f
C1032 _10_ input6/a_27_47# 4.57e-20
C1033 _01_ net5 0.0779f
C1034 _47_/a_81_21# _22_ 7.25e-19
C1035 net15 _42_/a_209_311# 0.0157f
C1036 net11 input10/a_27_47# 0.112f
C1037 th08_0/m1_477_n803# th04_0/m1_892_n998# 0.00566f
C1038 net4 _41_/a_59_75# 1.76e-19
C1039 _35_/a_76_199# _21_ 0.0175f
C1040 p[13] th14_0/m1_891_419# 0.0575f
C1041 p[8] VGND 0.129f
C1042 net4 VGND 0.564f
C1043 net7 input5/a_664_47# 0.00199f
C1044 _17_ net15 0.195f
C1045 _02_ _54_/a_75_212# 6.6e-20
C1046 _42_/a_209_311# _06_ 1.66e-19
C1047 _33_/a_109_93# VGND -0.0132f
C1048 net10 _03_ 0.321f
C1049 _23_ _36_/a_109_47# 3.44e-19
C1050 _03_ _10_ 0.00244f
C1051 _03_ _18_ 7.25e-23
C1052 _53_/a_29_53# _38_/a_27_47# 1.29e-19
C1053 net8 _16_ 0.00624f
C1054 net3 _16_ 1.77e-19
C1055 _17_ _06_ 0.0341f
C1056 _12_ net2 1.02e-20
C1057 _21_ net5 0.00784f
C1058 net4 _50_/a_223_47# 0.0107f
C1059 _36_/a_27_47# _30_/a_215_297# 7.13e-20
C1060 _24_ _11_ 7.29e-20
C1061 _10_ _14_ 0.0571f
C1062 net5 _42_/a_109_93# 0.00109f
C1063 p[13] net2 0.0301f
C1064 _26_/a_29_53# _12_ 0.00243f
C1065 _18_ _14_ 0.243f
C1066 net11 _35_/a_76_199# 4e-19
C1067 _48_/a_181_47# VGND 3.03e-19
C1068 _26_/a_183_297# VPWR -3.03e-19
C1069 _52_/a_93_21# _53_/a_29_53# 0.00116f
C1070 _52_/a_250_297# VGND -0.00314f
C1071 _43_/a_27_47# _11_ 4.27e-19
C1072 _27_/a_27_297# VGND -0.0157f
C1073 _20_ net14 8.01e-20
C1074 net17 net19 8.84e-23
C1075 net11 net5 0.0129f
C1076 _05_ net12 0.0414f
C1077 VPWR _25_ 0.0829f
C1078 _21_ input12/a_27_47# 2.32e-19
C1079 input13/a_27_47# net9 2.42e-19
C1080 _00_ _12_ 0.00396f
C1081 net19 input5/a_558_47# 2.24e-20
C1082 VGND th13_0/m1_559_n458# 0.0449f
C1083 VPWR _36_/a_27_47# -0.00832f
C1084 _09_ net12 0.0374f
C1085 _01_ VGND 0.0939f
C1086 _30_/a_215_297# _29_/a_29_53# 1.72e-19
C1087 _30_/a_215_297# _06_ 2.03e-20
C1088 Vin output17/a_27_47# 0.00661f
C1089 Vin net1 0.0121f
C1090 _17_ _39_/a_285_47# 7.36e-21
C1091 _04_ _05_ 0.0352f
C1092 _35_/a_226_297# VGND -4.55e-19
C1093 net17 b[1] 0.0287f
C1094 _31_/a_35_297# net7 0.0384f
C1095 _08_ _02_ 2.26e-20
C1096 _30_/a_465_297# net13 6.36e-20
C1097 net14 _50_/a_343_93# 1.07e-20
C1098 _04_ _09_ 0.0904f
C1099 net11 input12/a_27_47# 0.00246f
C1100 _25_ b[2] 0.0015f
C1101 _21_ VGND 0.295f
C1102 VPWR net15 0.61f
C1103 _03_ _33_/a_209_311# 8.38e-19
C1104 _35_/a_76_199# net7 1.79e-20
C1105 b[1] _49_/a_75_199# 0.00805f
C1106 _31_/a_285_297# th03_0/m1_890_n844# 3.4e-20
C1107 th04_0/m1_892_n998# th03_0/m1_890_n844# 0.00159f
C1108 VPWR _53_/a_111_297# 1.11e-34
C1109 VGND _42_/a_109_93# -0.0045f
C1110 b[1] input5/a_558_47# 0.00214f
C1111 _43_/a_193_413# th15_0/Vin 5.52e-19
C1112 _06_ _50_/a_615_93# 0.00264f
C1113 output18/a_27_47# net18 0.0106f
C1114 _44_/a_256_47# p[14] 6.02e-21
C1115 _20_ _16_ 0.00271f
C1116 th11_0/m1_705_187# input1/a_75_212# 5.25e-20
C1117 VPWR _29_/a_29_53# 0.0299f
C1118 VPWR _06_ 1.4f
C1119 _28_/a_109_297# _14_ 5.66e-19
C1120 _18_ input5/a_664_47# 1.09e-20
C1121 Vin _37_/a_27_47# 2.88e-19
C1122 input3/a_27_47# p[11] 0.0153f
C1123 _35_/a_226_47# input13/a_27_47# 3.94e-20
C1124 _21_ _50_/a_223_47# 2.91e-21
C1125 _02_ _39_/a_47_47# 0.0127f
C1126 net7 net5 0.195f
C1127 _14_ p[11] 1.27e-19
C1128 th03_0/m1_890_n844# input8/a_27_47# 0.00179f
C1129 _22_ _38_/a_27_47# 2.86e-19
C1130 Vin th10_0/m1_502_n495# 9.53e-19
C1131 net15 p[12] 1.84e-19
C1132 net11 VGND 0.475f
C1133 _35_/a_76_199# net6 4.6e-21
C1134 b[1] input5/a_62_47# 0.0024f
C1135 net1 p[6] 3.12e-20
C1136 _43_/a_469_47# net14 1.44e-20
C1137 VPWR th05_0/m1_752_n794# 0.0162f
C1138 _03_ _27_/a_109_297# 1.97e-20
C1139 _17_ _50_/a_27_47# 3.93e-20
C1140 _49_/a_208_47# _02_ 0.00193f
C1141 VGND p[1] 0.197f
C1142 input13/a_27_47# p[4] 7.37e-20
C1143 th15_0/Vin p[9] 0.228f
C1144 th11_0/m1_705_187# b[1] 0.00504f
C1145 p[12] _06_ 0.0132f
C1146 Vin _11_ 1.06e-19
C1147 net16 net18 0.00585f
C1148 _52_/a_93_21# _22_ 0.0347f
C1149 p[5] net11 0.0625f
C1150 _08_ net13 1.82e-19
C1151 th15_0/Vin _15_ 0.00389f
C1152 net15 _55_/a_217_297# 7.79e-19
C1153 _27_/a_205_297# _15_ 5.5e-20
C1154 net10 net18 3.35e-20
C1155 _31_/a_35_297# _55_/a_80_21# 5.9e-21
C1156 net5 net6 0.727f
C1157 b[2] _06_ 0.0116f
C1158 _43_/a_193_413# _44_/a_93_21# 0.0161f
C1159 _30_/a_297_297# net12 7.14e-21
C1160 net3 _47_/a_299_297# 2.55e-19
C1161 _55_/a_217_297# _06_ 3.46e-19
C1162 _32_/a_303_47# net5 7.18e-21
C1163 p[10] th02_0/m1_983_133# 1.21e-20
C1164 _12_ _39_/a_377_297# 6.77e-19
C1165 net10 input10/a_27_47# 0.00321f
C1166 VPWR _39_/a_285_47# -9.53e-19
C1167 _32_/a_27_47# net12 1.52e-19
C1168 b[1] net9 0.0765f
C1169 net8 net19 1.15e-19
C1170 net3 net19 0.611f
C1171 net14 _22_ 2.23e-19
C1172 _45_/a_27_47# _12_ 0.0867f
C1173 _43_/a_297_47# _17_ 5.72e-20
C1174 _55_/a_80_21# net5 2.78e-19
C1175 _17_ input6/a_27_47# 7.13e-22
C1176 VPWR _45_/a_193_297# -0.00859f
C1177 _12_ _23_ 0.00743f
C1178 _19_ p[10] 9.65e-20
C1179 _06_ input4/a_75_212# 0.00205f
C1180 _32_/a_109_47# _02_ 3.98e-19
C1181 _27_/a_27_297# net17 0.00181f
C1182 p[8] input5/a_62_47# 1.22e-19
C1183 _31_/a_35_297# net10 3.95e-20
C1184 _47_/a_384_47# net5 0.00129f
C1185 _04_ _32_/a_27_47# 1.43e-19
C1186 th12_0/m1_394_n856# th15_0/Vin 0.0254f
C1187 _44_/a_93_21# _15_ 0.0168f
C1188 VGND net7 0.421f
C1189 Vin th13_0/m1_831_275# 0.0354f
C1190 _39_/a_285_47# p[12] 3.03e-19
C1191 VGND _50_/a_515_93# -4.75e-19
C1192 b[3] net6 8.06e-19
C1193 _45_/a_205_47# net6 2.59e-20
C1194 _27_/a_27_297# _49_/a_75_199# 0.011f
C1195 th14_0/m1_641_n318# p[11] 0.114f
C1196 _35_/a_76_199# net10 0.0226f
C1197 _27_/a_27_297# input5/a_558_47# 1.57e-19
C1198 _05_ output17/a_27_47# 1.12e-19
C1199 input3/a_27_47# _42_/a_209_311# 1.56e-19
C1200 _35_/a_76_199# _10_ 7.19e-20
C1201 _05_ net1 0.151f
C1202 _14_ _42_/a_209_311# 0.00142f
C1203 _15_ _42_/a_296_53# 1.28e-19
C1204 th01_0/m1_991_n1219# p[0] 0.172f
C1205 VPWR p[0] 0.27f
C1206 _35_/a_76_199# _18_ 6.82e-21
C1207 Vin _27_/a_277_297# 1.98e-20
C1208 _45_/a_193_297# p[12] 5.2e-20
C1209 b[1] net8 0.0729f
C1210 _01_ net17 0.0988f
C1211 net3 b[1] 0.00334f
C1212 _31_/a_117_297# b[1] 0.00281f
C1213 _31_/a_285_47# net17 0.00134f
C1214 _09_ net1 5.26e-20
C1215 net16 net5 0.00476f
C1216 net6 _41_/a_59_75# 0.0373f
C1217 _17_ _14_ 0.489f
C1218 _02_ net13 0.00154f
C1219 net10 net5 0.0316f
C1220 VGND net6 0.512f
C1221 _43_/a_193_413# _04_ 5.67e-21
C1222 _04_ _49_/a_315_47# 7.71e-19
C1223 _01_ _49_/a_75_199# 0.009f
C1224 _35_/a_226_47# b[1] 0.00334f
C1225 _10_ net5 0.199f
C1226 b[1] _07_ 0.0417f
C1227 _01_ input5/a_558_47# 3.97e-20
C1228 VPWR _50_/a_27_47# -0.00335f
C1229 _18_ net5 0.0426f
C1230 net4 net9 1.99e-22
C1231 _22_ _16_ 3.8e-19
C1232 _34_/a_285_47# net12 8.07e-20
C1233 _33_/a_109_93# net9 0.00211f
C1234 _32_/a_303_47# VGND -4.83e-19
C1235 _20_ _47_/a_299_297# 0.002f
C1236 _48_/a_27_47# _07_ 0.0524f
C1237 th08_0/m1_477_n803# b[1] 6.6e-21
C1238 net6 _50_/a_223_47# 0.0194f
C1239 b[1] p[4] 0.0136f
C1240 net17 _42_/a_109_93# 3.1e-21
C1241 p[13] _19_ 0.00101f
C1242 input14/a_27_47# p[11] 3.98e-20
C1243 _21_ _49_/a_75_199# 6.64e-19
C1244 input9/a_75_212# VGND 0.0631f
C1245 _12_ _24_ 1.67e-19
C1246 p[12] _50_/a_27_47# 1.55e-19
C1247 VGND _55_/a_80_21# 0.00281f
C1248 output18/a_27_47# VGND 0.0581f
C1249 _20_ net19 1.29e-19
C1250 _03_ _30_/a_215_297# 0.0393f
C1251 p[7] _34_/a_47_47# 2.81e-19
C1252 p[3] net13 0.00398f
C1253 _04_ _15_ 3.61e-20
C1254 input5/a_558_47# _42_/a_109_93# 1.75e-19
C1255 net10 input12/a_27_47# 0.00182f
C1256 _47_/a_384_47# VGND -2.05e-19
C1257 _43_/a_27_47# _12_ 2.33e-21
C1258 p[14] th10_0/m1_536_174# 3.8e-19
C1259 p[8] net3 1.87e-19
C1260 net4 net3 9.28e-21
C1261 th15_0/m1_849_n157# _15_ 2.53e-19
C1262 _43_/a_297_47# VPWR -2.11e-19
C1263 net11 net17 3.19e-20
C1264 _10_ b[3] 6.63e-21
C1265 VPWR input6/a_27_47# 0.00129f
C1266 _45_/a_205_47# _10_ 6.19e-20
C1267 _13_ _04_ 1.17e-21
C1268 net17 p[1] 8.41e-20
C1269 _09_ _11_ 0.0665f
C1270 _18_ th12_0/m1_529_n42# 1.01e-20
C1271 net11 _49_/a_75_199# 4.49e-19
C1272 _43_/a_369_47# net6 3.62e-21
C1273 th14_0/m1_641_n318# _42_/a_209_311# 1.87e-19
C1274 input5/a_664_47# _42_/a_209_311# 0.0124f
C1275 _35_/a_76_199# _33_/a_209_311# 9.95e-21
C1276 _35_/a_226_47# _33_/a_109_93# 4.9e-19
C1277 _33_/a_296_53# _06_ 1.11e-20
C1278 _33_/a_109_93# _07_ 3.2e-19
C1279 net16 VGND 0.144f
C1280 _01_ net9 0.157f
C1281 _10_ _41_/a_59_75# 0.0235f
C1282 net2 input7/a_27_47# 3.24e-19
C1283 input5/a_558_47# p[1] 1.61e-21
C1284 net10 VGND 0.446f
C1285 VPWR _03_ 0.835f
C1286 _20_ b[1] 0.00465f
C1287 _24_ _34_/a_47_47# 6.84e-21
C1288 _10_ VGND 1.15f
C1289 net1 _30_/a_297_297# 7.34e-20
C1290 _05_ _33_/a_368_53# 9.2e-19
C1291 _18_ VGND 0.0166f
C1292 net15 th15_0/Vin 0.00757f
C1293 th14_0/m1_891_419# th11_0/m1_577_n654# 0.0383f
C1294 output19/a_27_47# p[14] 0.0459f
C1295 VPWR input3/a_27_47# 0.0688f
C1296 _40_/a_191_297# net2 0.00143f
C1297 _27_/a_27_297# net8 0.0108f
C1298 _27_/a_27_297# net3 0.0166f
C1299 VPWR _14_ 0.186f
C1300 p[5] net10 0.00544f
C1301 p[10] Vin 0.0929f
C1302 net16 _50_/a_223_47# 4.77e-21
C1303 _48_/a_181_47# _07_ 5.93e-19
C1304 _32_/a_27_47# net1 0.0211f
C1305 _35_/a_226_47# _52_/a_250_297# 2.63e-20
C1306 b[1] _53_/a_29_53# 4.99e-19
C1307 _10_ _50_/a_223_47# 0.0295f
C1308 _52_/a_346_47# _06_ 0.0031f
C1309 th15_0/Vin _06_ 0.00739f
C1310 _21_ net9 0.0282f
C1311 input2/a_27_47# input7/a_27_47# 1.62e-19
C1312 _18_ _50_/a_223_47# 0.0367f
C1313 _45_/a_109_297# _11_ 0.00168f
C1314 _10_ _53_/a_183_297# 2.86e-19
C1315 input15/a_27_47# p[14] 0.00367f
C1316 net2 th11_0/m1_577_n654# 0.0079f
C1317 _01_ net8 0.0802f
C1318 net3 _01_ 1.16e-19
C1319 _31_/a_285_47# net8 0.00129f
C1320 _53_/a_29_53# _48_/a_27_47# 3.14e-21
C1321 net17 net7 0.2f
C1322 p[14] _37_/a_197_47# 1.52e-19
C1323 VGND th02_0/m1_571_144# 0.00939f
C1324 _00_ _39_/a_47_47# 1.85e-20
C1325 net7 _49_/a_75_199# 0.09f
C1326 b[1] th03_0/m1_890_n844# 3.03e-20
C1327 net11 net9 0.136f
C1328 net7 input5/a_558_47# 0.00358f
C1329 _44_/a_93_21# net15 0.00573f
C1330 net4 _20_ 3.01e-20
C1331 _31_/a_285_297# input8/a_27_47# 1.04e-19
C1332 _55_/a_217_297# _14_ 0.0116f
C1333 _55_/a_472_297# _15_ 0.00626f
C1334 VPWR _49_/a_201_297# 0.0175f
C1335 net2 p[14] 5.39e-19
C1336 _26_/a_29_53# _02_ 0.0466f
C1337 _25_ net12 4.46e-20
C1338 net8 _21_ 0.00656f
C1339 _43_/a_369_47# _10_ 0.00199f
C1340 _12_ Vin 2.56e-21
C1341 _43_/a_369_47# _18_ 1.49e-19
C1342 net3 _42_/a_109_93# 0.0435f
C1343 p[11] th12_0/m1_529_n42# 0.0172f
C1344 _36_/a_27_47# net12 0.0185f
C1345 _35_/a_226_47# _21_ 9.87e-19
C1346 p[13] Vin 0.242f
C1347 _21_ _07_ 0.133f
C1348 net4 _53_/a_29_53# 3.26e-19
C1349 net7 input5/a_62_47# 2.04e-19
C1350 _32_/a_27_47# _11_ 1.65e-20
C1351 _22_ net19 2.17e-19
C1352 _33_/a_209_311# VGND -0.00749f
C1353 _28_/a_109_297# VGND -9.87e-19
C1354 th11_0/m1_705_187# net7 1.13e-19
C1355 _43_/a_193_413# _37_/a_27_47# 0.0102f
C1356 th14_0/m1_641_n318# VPWR 0.00238f
C1357 th06_0/m1_904_n796# VPWR 0.00203f
C1358 VGND p[11] 0.224f
C1359 _00_ _02_ 0.0269f
C1360 _04_ _36_/a_27_47# 0.00169f
C1361 VPWR input5/a_664_47# 0.00488f
C1362 net14 _16_ 0.00266f
C1363 net11 net8 1.5e-19
C1364 _20_ _27_/a_27_297# 3.14e-20
C1365 net4 _50_/a_343_93# 0.00124f
C1366 net5 _42_/a_209_311# 3.27e-21
C1367 net3 p[1] 1.67e-20
C1368 net11 _35_/a_226_47# 3.21e-19
C1369 net11 _07_ 0.0206f
C1370 Vin _34_/a_47_47# 5.61e-19
C1371 VPWR th01_0/m1_571_n501# 0.0263f
C1372 _17_ net5 0.00408f
C1373 _52_/a_256_47# VGND -0.00161f
C1374 th15_0/Vin p[0] 0.336f
C1375 _43_/a_193_413# _11_ 5.45e-19
C1376 _26_/a_29_53# net13 2.23e-20
C1377 _29_/a_29_53# net12 0.0132f
C1378 _27_/a_109_297# VGND -6.15e-19
C1379 net12 _06_ 0.284f
C1380 net9 net7 0.00233f
C1381 _20_ _01_ 0.161f
C1382 b[1] _22_ 9.74e-20
C1383 _04_ net15 0.0569f
C1384 _37_/a_27_47# p[9] 0.0117f
C1385 net11 p[4] 0.0557f
C1386 th08_0/m1_477_n803# net11 1.78e-19
C1387 _37_/a_27_47# _15_ 1.11e-19
C1388 VPWR net18 0.104f
C1389 th15_0/Vin _50_/a_27_47# 2.06e-19
C1390 _31_/a_35_297# _30_/a_215_297# 6.37e-19
C1391 th10_0/m1_502_n495# p[9] 0.0156f
C1392 _08_ _23_ 1.81e-19
C1393 _04_ _29_/a_29_53# 0.0408f
C1394 th05_0/m1_752_n794# net12 5e-20
C1395 _05_ p[10] 6.39e-20
C1396 net10 net17 8.67e-21
C1397 _04_ _06_ 0.0132f
C1398 VPWR input14/a_27_47# 0.0739f
C1399 th15_0/m1_849_n157# _06_ 2.65e-19
C1400 _20_ _21_ 0.191f
C1401 VPWR input10/a_27_47# 0.0102f
C1402 _11_ p[9] 1.01e-19
C1403 _11_ _15_ 0.113f
C1404 _35_/a_556_47# VGND 1.95e-19
C1405 net3 net7 7.45e-20
C1406 _38_/a_197_47# _06_ 4.32e-19
C1407 net8 net7 0.295f
C1408 _31_/a_117_297# net7 0.00472f
C1409 _45_/a_27_47# _39_/a_47_47# 1.31e-19
C1410 _09_ _49_/a_544_297# 2.56e-20
C1411 _01_ _50_/a_343_93# 0.0131f
C1412 net14 _50_/a_429_93# 6.04e-21
C1413 _32_/a_303_47# net9 0.00218f
C1414 _17_ b[3] 5.76e-20
C1415 p[6] _34_/a_47_47# 0.00141f
C1416 _39_/a_47_47# _23_ 5.24e-21
C1417 _30_/a_215_297# net5 8.27e-21
C1418 _13_ _11_ 0.164f
C1419 net18 b[2] 0.0131f
C1420 th14_0/m1_891_419# input5/a_381_47# 4.77e-20
C1421 p[7] _08_ 0.00276f
C1422 _17_ th12_0/m1_529_n42# 1.35e-20
C1423 _21_ _53_/a_29_53# 0.00959f
C1424 _35_/a_226_47# net7 2.93e-20
C1425 VPWR _31_/a_35_297# 0.0284f
C1426 input9/a_75_212# net9 0.0245f
C1427 _43_/a_297_47# th15_0/Vin 2.63e-20
C1428 VGND _42_/a_209_311# -0.008f
C1429 p[2] input7/a_27_47# 0.0023f
C1430 net11 _20_ 0.00128f
C1431 th15_0/Vin input6/a_27_47# 0.00615f
C1432 output19/a_27_47# net2 0.00168f
C1433 net4 _22_ 0.0866f
C1434 _17_ _41_/a_59_75# 0.00149f
C1435 VPWR _35_/a_76_199# -0.00947f
C1436 _33_/a_109_93# _22_ 1.34e-22
C1437 net3 net6 0.00152f
C1438 _17_ VGND 0.313f
C1439 _12_ _05_ 2.52e-19
C1440 net2 input5/a_381_47# 0.0138f
C1441 _36_/a_197_47# _25_ 2.37e-21
C1442 net11 _53_/a_29_53# 8.31e-19
C1443 _32_/a_303_47# net8 2.22e-34
C1444 _49_/a_208_47# p[2] 4.19e-20
C1445 _45_/a_27_47# _02_ 0.00449f
C1446 _12_ _09_ 0.00526f
C1447 VPWR net5 0.613f
C1448 _03_ _27_/a_205_297# 1.46e-20
C1449 input15/a_27_47# net2 0.00296f
C1450 th14_0/m1_891_419# net2 0.011f
C1451 _17_ _50_/a_223_47# 5.24e-20
C1452 _02_ _23_ 0.0648f
C1453 input3/a_27_47# th15_0/Vin 0.00105f
C1454 _19_ input7/a_27_47# 3.12e-21
C1455 _52_/a_250_297# _22_ 0.0996f
C1456 th15_0/Vin _14_ 0.00355f
C1457 net2 _37_/a_197_47# 4.74e-20
C1458 net8 _55_/a_80_21# 1.84e-21
C1459 net1 _36_/a_27_47# 6.99e-20
C1460 _13_ th13_0/m1_831_275# 6e-20
C1461 net3 _55_/a_80_21# 2.35e-19
C1462 net10 net9 0.111f
C1463 _10_ net9 0.0438f
C1464 net17 _33_/a_209_311# 7.03e-21
C1465 _18_ net9 1.51e-19
C1466 _44_/a_93_21# input6/a_27_47# 8.53e-19
C1467 _01_ _47_/a_81_21# 6.05e-21
C1468 net12 _50_/a_27_47# 7.99e-21
C1469 _02_ p[2] 8.49e-19
C1470 p[12] net5 0.00392f
C1471 _05_ _34_/a_47_47# 1.26e-20
C1472 _12_ _39_/a_129_47# 0.00175f
C1473 VGND _30_/a_215_297# 0.00693f
C1474 b[2] net5 7.33e-20
C1475 _19_ _49_/a_208_47# 7.12e-20
C1476 th03_0/m1_890_n844# p[1] 0.00745f
C1477 net14 net19 0.148f
C1478 _01_ _22_ 0.15f
C1479 _20_ net7 0.0257f
C1480 VPWR input12/a_27_47# 0.0648f
C1481 _02_ _30_/a_109_53# 5.03e-22
C1482 _08_ _34_/a_129_47# 3.29e-19
C1483 _45_/a_109_297# _12_ 0.00587f
C1484 net15 net1 7.44e-20
C1485 _43_/a_369_47# _17_ 5.87e-19
C1486 _04_ _50_/a_27_47# 2.07e-21
C1487 VGND _38_/a_109_47# 2.3e-19
C1488 _55_/a_217_297# net5 8.84e-20
C1489 _19_ th11_0/m1_577_n654# 3.11e-19
C1490 _36_/a_197_47# _06_ 6.18e-19
C1491 b[1] _52_/a_93_21# 2.82e-19
C1492 VPWR b[3] 0.129f
C1493 VPWR _45_/a_205_47# -1.62e-19
C1494 VPWR th12_0/m1_529_n42# 0.0444f
C1495 net2 input2/a_27_47# 0.024f
C1496 net10 net8 2.05e-21
C1497 net1 _29_/a_29_53# 9.76e-19
C1498 _10_ net8 5.86e-19
C1499 net3 _10_ 3.89e-19
C1500 _23_ net13 4.11e-19
C1501 net1 _06_ 0.0115f
C1502 _44_/a_93_21# _14_ 0.04f
C1503 _44_/a_250_297# _15_ 0.00517f
C1504 net15 input5/a_841_47# 0.00585f
C1505 _18_ net8 1.15e-21
C1506 _18_ net3 7.34e-20
C1507 _19_ _02_ 0.213f
C1508 p[3] p[2] 0.0558f
C1509 _45_/a_465_47# net6 6.06e-20
C1510 VGND _50_/a_615_93# -5.19e-19
C1511 _20_ net6 9.69e-20
C1512 _21_ _22_ 0.00314f
C1513 _11_ _25_ 7.05e-19
C1514 _35_/a_226_47# net10 0.018f
C1515 VPWR _41_/a_59_75# 0.0186f
C1516 net5 input4/a_75_212# 0.0104f
C1517 net10 _07_ 0.0605f
C1518 input5/a_62_47# p[11] 0.00153f
C1519 _35_/a_226_47# _10_ 1.25e-19
C1520 _00_ net2 0.00732f
C1521 _10_ _07_ 2.19e-19
C1522 _22_ _42_/a_109_93# 1.21e-19
C1523 th01_0/m1_991_n1219# VGND 6.29e-19
C1524 VPWR VGND 0.267f
C1525 p[7] p[3] 0.0834f
C1526 _24_ _02_ 0.0232f
C1527 input5/a_841_47# _06_ 1.66e-19
C1528 net14 b[1] 0.00256f
C1529 p[3] _30_/a_109_53# 5.57e-19
C1530 _31_/a_285_297# b[1] 0.0101f
C1531 th04_0/m1_892_n998# b[1] 2.07e-20
C1532 _26_/a_29_53# _00_ 0.0466f
C1533 _32_/a_303_47# _20_ 1.54e-19
C1534 net15 _37_/a_27_47# 0.0541f
C1535 net4 _38_/a_27_47# 0.0119f
C1536 _43_/a_27_47# _02_ 1.88e-21
C1537 p[5] VPWR 0.165f
C1538 net10 p[4] 0.00273f
C1539 _53_/a_29_53# net6 2.11e-20
C1540 th14_0/m1_641_n318# th15_0/Vin 7.77e-19
C1541 _35_/a_489_413# b[1] 0.00104f
C1542 p[7] net13 0.00514f
C1543 th15_0/Vin input5/a_664_47# 2.16e-19
C1544 th03_0/m1_890_n844# net7 2.87e-19
C1545 _03_ net12 0.0268f
C1546 VPWR _50_/a_223_47# -0.00601f
C1547 _30_/a_109_53# net13 1.05e-19
C1548 p[12] _41_/a_59_75# 0.0048f
C1549 net19 _16_ 0.206f
C1550 net11 _22_ 6.82e-21
C1551 _20_ _55_/a_80_21# 0.0291f
C1552 b[1] input8/a_27_47# 0.00172f
C1553 _37_/a_27_47# _06_ 2.5e-20
C1554 _33_/a_209_311# net9 4.33e-20
C1555 VGND p[12] 0.359f
C1556 _28_/a_109_297# net9 3.7e-19
C1557 net4 _52_/a_93_21# 7.93e-20
C1558 _20_ _47_/a_384_47# 1.72e-19
C1559 p[13] _32_/a_27_47# 6.49e-20
C1560 net6 _50_/a_343_93# 0.00214f
C1561 net15 _11_ 0.145f
C1562 VGND b[2] 0.0779f
C1563 _08_ Vin 2.97e-19
C1564 th15_0/Vin th01_0/m1_571_n501# 0.00971f
C1565 net17 _42_/a_209_311# 1.04e-21
C1566 _52_/a_93_21# _33_/a_109_93# 2.89e-21
C1567 _04_ _03_ 0.586f
C1568 _19_ net13 4.45e-20
C1569 output18/a_27_47# _53_/a_29_53# 9.46e-19
C1570 VGND _55_/a_217_297# -0.00342f
C1571 _11_ _06_ 0.493f
C1572 _36_/a_109_47# _25_ 3.76e-21
C1573 _04_ input3/a_27_47# 3.55e-19
C1574 net4 b[0] 0.0024f
C1575 _04_ _14_ 2.04e-21
C1576 input5/a_558_47# _42_/a_209_311# 7.85e-20
C1577 _43_/a_193_413# _12_ 7.94e-22
C1578 Vin input7/a_27_47# 0.0085f
C1579 p[8] net14 0.01f
C1580 net4 net14 2.21e-21
C1581 b[1] _16_ 2.21e-19
C1582 _43_/a_369_47# VPWR -3.75e-19
C1583 _41_/a_59_75# input4/a_75_212# 0.00153f
C1584 th15_0/Vin input14/a_27_47# 0.00489f
C1585 _17_ input5/a_558_47# 2.13e-21
C1586 _45_/a_465_47# _10_ 3.32e-19
C1587 net10 _20_ 3.23e-19
C1588 _44_/a_93_21# input5/a_664_47# 1.88e-20
C1589 _52_/a_93_21# _52_/a_250_297# -6.97e-22
C1590 _20_ _10_ 0.179f
C1591 VGND input4/a_75_212# 0.0528f
C1592 _20_ _18_ 0.0151f
C1593 VGND th04_0/m1_620_n488# 0.00107f
C1594 _44_/a_346_47# net2 1.64e-19
C1595 net3 p[11] 0.00765f
C1596 p[0] output17/a_27_47# 0.00839f
C1597 net1 p[0] 0.00473f
C1598 _43_/a_469_47# net6 4.85e-21
C1599 th14_0/m1_641_n318# _42_/a_296_53# 8.45e-21
C1600 _35_/a_226_47# _33_/a_209_311# 1.31e-19
C1601 _33_/a_368_53# _06_ 1.7e-19
C1602 _33_/a_209_311# _07_ 0.00859f
C1603 net16 _53_/a_29_53# 2.04e-20
C1604 _29_/a_183_297# net11 3.64e-19
C1605 _10_ _41_/a_145_75# 0.00148f
C1606 net10 _53_/a_29_53# 7.88e-22
C1607 _22_ net7 2.73e-20
C1608 p[3] th07_0/m1_808_n892# 6.45e-21
C1609 th15_0/m1_597_n912# net5 1.17e-19
C1610 _10_ _53_/a_29_53# 0.00779f
C1611 _08_ p[6] 5.04e-19
C1612 Vin th11_0/m1_577_n654# 0.0926f
C1613 _12_ _15_ 0.00833f
C1614 _40_/a_297_297# net2 0.00101f
C1615 _27_/a_27_297# net14 0.0118f
C1616 _27_/a_109_297# net3 5.45e-19
C1617 _27_/a_277_297# net15 1.93e-19
C1618 net17 _30_/a_215_297# 4.69e-20
C1619 _04_ _49_/a_201_297# 0.0253f
C1620 _47_/a_81_21# net6 2.14e-19
C1621 _21_ _38_/a_27_47# 3.87e-19
C1622 _36_/a_109_47# _06_ 0.00168f
C1623 _13_ _12_ 0.462f
C1624 _10_ _50_/a_343_93# 0.0284f
C1625 _52_/a_584_47# _06_ 0.00218f
C1626 th13_0/m1_559_n458# b[0] 5.75e-19
C1627 Vin _02_ 1.03e-20
C1628 _18_ _50_/a_343_93# 0.0276f
C1629 _22_ net6 0.163f
C1630 _45_/a_193_297# _11_ 0.0292f
C1631 net4 _16_ 2.73e-20
C1632 Vin p[14] 0.143f
C1633 _52_/a_93_21# _21_ 9.4e-19
C1634 net14 _01_ 8.29e-19
C1635 _31_/a_285_297# _01_ 1.92e-19
C1636 _52_/a_346_47# net5 7.03e-19
C1637 th15_0/Vin net5 0.00138f
C1638 _17_ net9 2.89e-23
C1639 _04_ input5/a_664_47# 6.73e-21
C1640 net11 _38_/a_27_47# 1.68e-20
C1641 VPWR net17 0.037f
C1642 _44_/a_250_297# net15 8.86e-20
C1643 b[1] input13/a_27_47# 0.00624f
C1644 _01_ input8/a_27_47# 1.43e-19
C1645 output18/a_27_47# _22_ 7.51e-19
C1646 _55_/a_472_297# _14_ 0.00192f
C1647 _55_/a_300_47# _15_ 1.42e-20
C1648 _55_/a_80_21# _22_ 0.00926f
C1649 _00_ _45_/a_27_47# 4.84e-20
C1650 net2 th02_0/m1_983_133# 3.55e-19
C1651 Vin p[3] 0.359f
C1652 _35_/a_556_47# _07_ 0.00128f
C1653 VPWR _49_/a_75_199# 0.0154f
C1654 _43_/a_469_47# _10_ 0.00124f
C1655 net14 _21_ 7.17e-21
C1656 _28_/a_109_297# _20_ 0.00221f
C1657 net11 _52_/a_93_21# 2.8e-19
C1658 VPWR input5/a_558_47# 0.0083f
C1659 _43_/a_469_47# _18_ 1.59e-19
C1660 net8 _42_/a_209_311# 7.7e-21
C1661 net3 _42_/a_209_311# 0.029f
C1662 net14 _42_/a_109_93# 0.00351f
C1663 _27_/a_27_297# _16_ 3.74e-22
C1664 _11_ _50_/a_27_47# 0.0592f
C1665 _08_ _05_ 0.00897f
C1666 VGND th15_0/m1_597_n912# 0.051f
C1667 _03_ output17/a_27_47# 1.94e-19
C1668 _03_ net1 0.298f
C1669 th03_0/m1_890_n844# th02_0/m1_571_144# 1.09e-20
C1670 _35_/a_489_413# _21_ 0.0448f
C1671 _02_ p[6] 0.00164f
C1672 Vin net13 0.00366f
C1673 _17_ net3 0.0698f
C1674 _17_ net8 4.52e-20
C1675 input10/a_27_47# net12 0.00115f
C1676 net15 _40_/a_109_297# 0.0016f
C1677 _19_ net2 0.101f
C1678 _33_/a_296_53# VGND -1.43e-19
C1679 _08_ _09_ 0.106f
C1680 input3/a_27_47# output17/a_27_47# 3.15e-19
C1681 input2/a_27_47# _30_/a_109_53# 1.54e-20
C1682 _47_/a_81_21# _10_ 0.0061f
C1683 th15_0/Vin b[3] 0.106f
C1684 _44_/a_93_21# net5 3.61e-20
C1685 _18_ _47_/a_81_21# 7.96e-20
C1686 _30_/a_215_297# net9 0.0456f
C1687 _37_/a_27_47# input6/a_27_47# 9.35e-19
C1688 VPWR input5/a_62_47# 0.0601f
C1689 _01_ _16_ 3.24e-19
C1690 th15_0/Vin th12_0/m1_529_n42# 0.0693f
C1691 net11 net14 9.95e-19
C1692 net16 _22_ 0.00606f
C1693 _40_/a_109_297# _06_ 0.00175f
C1694 net4 _50_/a_429_93# 4.16e-19
C1695 _00_ _30_/a_109_53# 3.67e-20
C1696 th03_0/m1_638_n591# th02_0/m1_983_133# 0.00168f
C1697 th11_0/m1_705_187# th01_0/m1_991_n1219# 7.73e-20
C1698 _10_ _22_ 0.0904f
C1699 VPWR th11_0/m1_705_187# 0.0375f
C1700 net14 p[1] 0.0025f
C1701 _26_/a_29_53# _24_ 2.11e-20
C1702 _18_ _22_ 0.0211f
C1703 _43_/a_27_47# net2 0.01f
C1704 _19_ input2/a_27_47# 5.26e-20
C1705 th15_0/Vin _41_/a_59_75# 0.00218f
C1706 Vin _34_/a_377_297# 1.75e-19
C1707 p[10] net15 0.00989f
C1708 _52_/a_346_47# VGND -0.00175f
C1709 th15_0/Vin VGND 1.04f
C1710 p[3] p[6] 8.32e-22
C1711 _09_ _39_/a_47_47# 7.7e-21
C1712 _27_/a_205_297# VGND -3.36e-19
C1713 Vin th10_0/m1_536_174# 0.102f
C1714 _35_/a_76_199# net12 0.0132f
C1715 _33_/a_109_93# input13/a_27_47# 0.00348f
C1716 b[1] net19 1e-19
C1717 input8/a_27_47# p[1] 5.13e-20
C1718 _04_ _31_/a_35_297# 1.89e-20
C1719 _12_ _25_ 1.23e-20
C1720 b[1] input1/a_75_212# 0.0074f
C1721 _37_/a_27_47# _14_ 0.00137f
C1722 VPWR net9 0.496f
C1723 net8 _30_/a_215_297# 8.14e-21
C1724 _09_ _49_/a_208_47# 5.43e-21
C1725 net5 net12 0.0674f
C1726 _12_ _36_/a_27_47# 0.00178f
C1727 _49_/a_201_297# net1 0.00304f
C1728 _04_ _35_/a_76_199# 0.0269f
C1729 _44_/a_93_21# b[3] 7.07e-20
C1730 _44_/a_93_21# th12_0/m1_529_n42# 7.97e-20
C1731 _32_/a_197_47# net5 5.61e-21
C1732 _43_/a_27_47# _00_ 0.0431f
C1733 _05_ _02_ 0.00163f
C1734 _11_ _14_ 0.0415f
C1735 _29_/a_111_297# net11 8.27e-19
C1736 _20_ _42_/a_209_311# 1.66e-20
C1737 Vin output19/a_27_47# 0.00177f
C1738 _04_ net5 0.00476f
C1739 _52_/a_93_21# net6 2.33e-19
C1740 net14 net7 2.23e-19
C1741 _31_/a_285_297# net7 0.00227f
C1742 p[8] th09_0/m1_485_n505# 0.00223f
C1743 _09_ _02_ 0.297f
C1744 _03_ _30_/a_392_297# 6.33e-19
C1745 net14 _50_/a_515_93# 1.39e-20
C1746 _44_/a_93_21# VGND -0.0223f
C1747 _29_/a_183_297# _10_ 6.24e-20
C1748 p[6] _34_/a_377_297# 6.3e-19
C1749 _17_ _20_ 0.102f
C1750 net4 _47_/a_299_297# 3.28e-19
C1751 _12_ net15 8.14e-21
C1752 _34_/a_47_47# _25_ 1.08e-19
C1753 net1 input5/a_664_47# 2.41e-19
C1754 output18/a_27_47# _38_/a_27_47# 8.6e-19
C1755 VPWR net8 0.701f
C1756 VPWR net3 0.351f
C1757 VPWR _31_/a_117_297# 5.04e-19
C1758 p[13] net15 0.00241f
C1759 input12/a_27_47# net12 0.0297f
C1760 _43_/a_369_47# th15_0/Vin 1.11e-19
C1761 b[1] _48_/a_27_47# 0.00666f
C1762 net6 b[0] 2.52e-19
C1763 _45_/a_27_47# _23_ 1.74e-19
C1764 p[8] net19 0.00885f
C1765 input15/a_27_47# Vin 0.00251f
C1766 net4 net19 2.65e-20
C1767 Vin th14_0/m1_891_419# 0.101f
C1768 input8/a_27_47# net7 1.47e-19
C1769 _12_ _06_ 0.136f
C1770 VPWR _35_/a_226_47# 0.00159f
C1771 VPWR _07_ 0.0728f
C1772 net14 net6 2.82e-21
C1773 _05_ p[3] 9.91e-20
C1774 _22_ p[11] 3.13e-20
C1775 _36_/a_303_47# _25_ 2.03e-21
C1776 _09_ p[3] 5.82e-20
C1777 _05_ net13 0.192f
C1778 _45_/a_109_297# _02_ 8.44e-19
C1779 _03_ _27_/a_277_297# 2.1e-20
C1780 VPWR p[4] 0.145f
C1781 VPWR th08_0/m1_477_n803# 0.0276f
C1782 Vin net2 0.0132f
C1783 net16 _38_/a_27_47# 0.114f
C1784 _17_ _50_/a_343_93# 0.0015f
C1785 VGND net12 0.344f
C1786 th15_0/m1_849_n157# b[3] 2.83e-20
C1787 _10_ _38_/a_27_47# 0.0133f
C1788 _09_ net13 0.0379f
C1789 net2 _37_/a_303_47# 4.41e-19
C1790 _20_ _30_/a_215_297# 6.08e-19
C1791 net7 _16_ 7.5e-20
C1792 th04_0/m1_892_n998# input9/a_75_212# 3.16e-20
C1793 p[10] p[0] 0.00247f
C1794 net3 _55_/a_217_297# 5.78e-20
C1795 net14 _55_/a_80_21# 4.7e-19
C1796 _27_/a_27_297# net19 1.98e-19
C1797 net15 _55_/a_300_47# 1.09e-19
C1798 _32_/a_197_47# VGND 8.12e-20
C1799 _34_/a_47_47# _06_ 0.0391f
C1800 p[5] net12 0.00294f
C1801 b[1] _33_/a_109_93# 0.00411f
C1802 _04_ VGND 0.135f
C1803 net10 _52_/a_93_21# 7.84e-20
C1804 _55_/a_300_47# _06_ 2.5e-20
C1805 Vin input2/a_27_47# 0.00133f
C1806 th15_0/m1_849_n157# _41_/a_59_75# 0.00112f
C1807 _10_ _52_/a_93_21# 0.00534f
C1808 _12_ _39_/a_285_47# 0.0221f
C1809 input8/a_27_47# input9/a_75_212# 3.09e-20
C1810 _18_ _52_/a_93_21# 1.97e-19
C1811 VGND th15_0/m1_849_n157# 0.0514f
C1812 p[2] th02_0/m1_983_133# 9.44e-20
C1813 _01_ net19 4.9e-19
C1814 net16 b[0] 0.0306f
C1815 net6 _16_ 1.62e-20
C1816 _20_ _50_/a_615_93# 8.8e-19
C1817 _08_ _34_/a_285_47# 0.00414f
C1818 Vin th03_0/m1_638_n591# 1.78e-19
C1819 _48_/a_181_47# b[1] 3.46e-19
C1820 _45_/a_27_47# _24_ 4.57e-19
C1821 _45_/a_193_297# _12_ 0.0103f
C1822 _31_/a_35_297# net1 0.0111f
C1823 VGND _38_/a_197_47# 2.29e-19
C1824 _43_/a_469_47# _17_ 0.00177f
C1825 _04_ _50_/a_223_47# 7.89e-22
C1826 VPWR _45_/a_465_47# -5.05e-19
C1827 _36_/a_303_47# _06_ 5.3e-19
C1828 _24_ _23_ 0.012f
C1829 VPWR _20_ 0.34f
C1830 _27_/a_27_297# b[1] 0.00644f
C1831 _44_/a_250_297# input3/a_27_47# 2.07e-19
C1832 _32_/a_27_47# _02_ 0.00247f
C1833 _31_/a_285_297# net10 1.68e-19
C1834 _19_ p[2] 1.1e-21
C1835 net14 _10_ 2.4e-19
C1836 net10 th04_0/m1_892_n998# 8.54e-21
C1837 _44_/a_250_297# _14_ 4.82e-19
C1838 _18_ net14 0.0147f
C1839 Vin output16/a_27_47# 3.69e-19
C1840 th15_0/Vin input5/a_558_47# 2.18e-19
C1841 _36_/a_197_47# net5 0.00254f
C1842 _35_/a_489_413# net10 0.00225f
C1843 VPWR _41_/a_145_75# -2.41e-19
C1844 _48_/a_109_47# p[6] 3.39e-21
C1845 _17_ _47_/a_81_21# 0.0456f
C1846 _35_/a_489_413# _10_ 3.41e-19
C1847 th08_0/m1_477_n803# th04_0/m1_620_n488# 6.4e-19
C1848 net19 _42_/a_109_93# 0.0448f
C1849 _55_/a_80_21# _16_ 0.0143f
C1850 _22_ _42_/a_209_311# 1.72e-19
C1851 VPWR _53_/a_29_53# 0.00821f
C1852 _01_ b[1] 0.00233f
C1853 input14/a_27_47# _11_ 1.42e-19
C1854 net1 net5 0.0772f
C1855 net5 output17/a_27_47# 5.01e-20
C1856 _31_/a_285_47# b[1] 8.76e-19
C1857 p[13] p[0] 2.15e-19
C1858 p[3] _30_/a_297_297# 3.04e-20
C1859 _26_/a_111_297# _00_ 3.7e-19
C1860 _17_ _22_ 0.00334f
C1861 _40_/a_109_297# _14_ -1.78e-33
C1862 _43_/a_193_413# _02_ 9.4e-21
C1863 _49_/a_315_47# _02_ 0.00134f
C1864 _12_ _50_/a_27_47# 0.00354f
C1865 _35_/a_226_297# b[1] 1.03e-19
C1866 _54_/a_75_212# _25_ 0.0247f
C1867 th15_0/Vin input5/a_62_47# 9.04e-19
C1868 net5 input5/a_841_47# 0.0221f
C1869 VPWR _50_/a_343_93# -0.0126f
C1870 _13_ _39_/a_47_47# 0.00117f
C1871 _30_/a_297_297# net13 3.27e-20
C1872 p[12] _41_/a_145_75# 4.82e-19
C1873 _43_/a_193_413# p[14] 1.34e-20
C1874 _20_ _55_/a_217_297# 0.0013f
C1875 th11_0/m1_705_187# th15_0/Vin 0.0346f
C1876 _03_ p[10] 8.74e-20
C1877 VPWR th03_0/m1_890_n844# 0.037f
C1878 b[1] _21_ 0.00892f
C1879 net4 _52_/a_250_297# 0.00136f
C1880 _53_/a_29_53# b[2] 6.22e-19
C1881 net6 _50_/a_429_93# 6.18e-19
C1882 b[1] _42_/a_109_93# 2.38e-19
C1883 _52_/a_250_297# _33_/a_109_93# 5.17e-22
C1884 input1/a_75_212# p[1] 0.0023f
C1885 _03_ _49_/a_544_297# 0.00568f
C1886 _44_/a_93_21# input5/a_558_47# 2.71e-19
C1887 net1 input12/a_27_47# 7.44e-20
C1888 _10_ _16_ 0.00486f
C1889 _37_/a_27_47# net5 1.13e-20
C1890 _02_ _34_/a_285_47# 7.14e-19
C1891 VGND _55_/a_472_297# -0.00188f
C1892 _18_ _16_ 0.144f
C1893 _35_/a_76_199# _11_ 6.99e-22
C1894 _21_ _48_/a_27_47# 0.0121f
C1895 _05_ net2 4.03e-20
C1896 _02_ _15_ 0.101f
C1897 p[7] th07_0/m1_808_n892# 0.012f
C1898 p[14] p[9] 0.0624f
C1899 p[14] _15_ 0.00339f
C1900 net11 b[1] 0.0777f
C1901 _30_/a_215_297# _22_ 2.46e-21
C1902 _43_/a_469_47# VPWR -2.75e-19
C1903 _13_ _02_ 0.0676f
C1904 _36_/a_197_47# VGND -3.75e-19
C1905 _52_/a_93_21# _52_/a_256_47# -6.6e-20
C1906 _44_/a_93_21# input5/a_62_47# 5.05e-20
C1907 _11_ net5 0.207f
C1908 net17 net12 2.11e-21
C1909 b[1] p[1] 0.00395f
C1910 _44_/a_584_47# net2 0.0053f
C1911 _54_/a_75_212# _06_ 0.00727f
C1912 net14 p[11] 4.35e-19
C1913 VGND output17/a_27_47# 0.00246f
C1914 net1 VGND 0.513f
C1915 net11 _48_/a_27_47# 0.0179f
C1916 th14_0/m1_641_n318# _42_/a_368_53# 2.53e-20
C1917 input9/a_75_212# input13/a_27_47# 0.00732f
C1918 _05_ input2/a_27_47# 1.83e-19
C1919 _35_/a_489_413# _33_/a_209_311# 2.77e-20
C1920 _12_ _03_ 2.76e-20
C1921 VPWR _47_/a_81_21# 0.0089f
C1922 net4 _21_ 0.00535f
C1923 _04_ net17 0.0218f
C1924 VGND input5/a_841_47# 0.0943f
C1925 input1/a_75_212# net7 3.77e-19
C1926 _00_ _05_ 5.03e-22
C1927 _21_ _33_/a_109_93# 1.62e-20
C1928 net3 th15_0/Vin 0.00715f
C1929 net8 th15_0/Vin 1.56e-21
C1930 _12_ _14_ 1.98e-20
C1931 _34_/a_285_47# net13 4.11e-20
C1932 _27_/a_27_297# _01_ 8.04e-19
C1933 _27_/a_109_297# net14 1.32e-19
C1934 _27_/a_205_297# net3 4.37e-19
C1935 VPWR _22_ 1.4f
C1936 p[13] input3/a_27_47# 0.00527f
C1937 _47_/a_299_297# net6 3.63e-19
C1938 th03_0/m1_890_n844# th04_0/m1_620_n488# 0.00138f
C1939 _04_ _49_/a_75_199# 0.0782f
C1940 _00_ _09_ 9.35e-21
C1941 Vin p[2] 0.165f
C1942 _04_ input5/a_558_47# 1.25e-20
C1943 _10_ _50_/a_429_93# 0.00167f
C1944 _44_/a_250_297# input14/a_27_47# 8.25e-21
C1945 net19 net6 0.00346f
C1946 VGND _37_/a_27_47# -0.0147f
C1947 _13_ net13 4e-21
C1948 p[7] Vin 0.474f
C1949 Vin _30_/a_109_53# 1.09e-19
C1950 Vin th02_0/m1_983_133# 0.062f
C1951 _36_/a_109_47# net5 0.00144f
C1952 net10 input13/a_27_47# 8.86e-20
C1953 _03_ _34_/a_47_47# 4.5e-20
C1954 th10_0/m1_502_n495# VGND 0.0046f
C1955 net11 _33_/a_109_93# 5.14e-19
C1956 _31_/a_285_47# _01_ 3.36e-19
C1957 b[1] net7 0.0783f
C1958 p[12] _22_ 4.34e-21
C1959 _52_/a_584_47# net5 0.0022f
C1960 _28_/a_109_297# _16_ 1.26e-19
C1961 _16_ p[11] 1.76e-19
C1962 _04_ input5/a_62_47# 0.00345f
C1963 _27_/a_27_297# _42_/a_109_93# 1.35e-20
C1964 _11_ _41_/a_59_75# 8.7e-19
C1965 _22_ b[2] 0.0043f
C1966 _00_ _39_/a_129_47# 1.63e-20
C1967 VGND _11_ 0.091f
C1968 th10_0/m1_536_174# p[9] 0.185f
C1969 p[10] th01_0/m1_571_n501# 0.006f
C1970 _19_ Vin 0.00421f
C1971 _44_/a_93_21# net3 0.0102f
C1972 _55_/a_80_21# net19 0.00423f
C1973 _55_/a_300_47# _14_ 8.09e-19
C1974 _00_ _45_/a_109_297# 4.86e-20
C1975 _08_ _06_ 0.0343f
C1976 _01_ _21_ 7.94e-19
C1977 p[13] _49_/a_201_297# 6.25e-20
C1978 net9 net12 0.0596f
C1979 net11 _52_/a_250_297# 1.2e-19
C1980 net11 _27_/a_27_297# 1.58e-20
C1981 net15 input7/a_27_47# 1.88e-19
C1982 net14 _42_/a_209_311# 0.0238f
C1983 net3 _42_/a_296_53# 1.81e-19
C1984 _11_ _50_/a_223_47# 0.0329f
C1985 _32_/a_197_47# net9 6.06e-19
C1986 VPWR _29_/a_183_297# -8.13e-19
C1987 VGND _30_/a_392_297# 3.41e-19
C1988 net15 _39_/a_47_47# 9.44e-22
C1989 _27_/a_27_297# p[1] 2.87e-19
C1990 _43_/a_193_413# input15/a_27_47# 1.62e-20
C1991 _17_ net14 0.104f
C1992 _02_ _25_ 0.0156f
C1993 net15 _40_/a_191_297# 8.41e-19
C1994 p[7] p[6] 0.196f
C1995 _04_ net9 0.0213f
C1996 _33_/a_368_53# VGND 2.38e-19
C1997 _47_/a_299_297# _10_ 0.0134f
C1998 _44_/a_250_297# net5 3.11e-20
C1999 output19/a_27_47# p[9] 0.0933f
C2000 _02_ _36_/a_27_47# 9.37e-20
C2001 _39_/a_47_47# _06_ 1.44e-19
C2002 net11 _01_ 3.82e-20
C2003 b[1] input9/a_75_212# 0.00598f
C2004 th14_0/m1_641_n318# p[13] 0.00188f
C2005 p[13] input5/a_664_47# 0.0024f
C2006 b[1] _55_/a_80_21# 6.03e-19
C2007 _40_/a_191_297# _06_ 5.84e-19
C2008 b[1] output18/a_27_47# 9.26e-19
C2009 _10_ net19 3.43e-19
C2010 net8 net12 0.00458f
C2011 VGND th13_0/m1_831_275# 0.0456f
C2012 _18_ net19 4.89e-20
C2013 _43_/a_193_413# net2 1.52e-19
C2014 VGND _36_/a_109_47# 3.56e-19
C2015 th15_0/Vin _41_/a_145_75# 1.73e-19
C2016 _32_/a_197_47# net8 3.39e-20
C2017 _31_/a_35_297# p[10] 3.66e-19
C2018 _52_/a_584_47# VGND -0.00112f
C2019 Vin th07_0/m1_808_n892# 0.0314f
C2020 _27_/a_277_297# VGND -4.65e-19
C2021 input15/a_27_47# p[9] 0.0194f
C2022 _00_ _32_/a_27_47# 0.00228f
C2023 _35_/a_226_47# net12 8.29e-19
C2024 _45_/a_27_47# _05_ 9.34e-23
C2025 input15/a_27_47# _15_ 2.15e-20
C2026 net12 _07_ 0.18f
C2027 _33_/a_209_311# input13/a_27_47# 5.85e-20
C2028 net11 _21_ 0.586f
C2029 net15 _02_ 0.0806f
C2030 p[8] net6 1.3e-20
C2031 VPWR _38_/a_27_47# -0.0142f
C2032 _04_ net8 0.02f
C2033 _04_ net3 0.113f
C2034 net4 net6 0.713f
C2035 _12_ net18 8.24e-19
C2036 _02_ _53_/a_111_297# 9.57e-20
C2037 net17 output17/a_27_47# 0.0149f
C2038 net17 net1 2.89e-19
C2039 _42_/a_209_311# _16_ 0.00129f
C2040 _37_/a_197_47# _15_ 3.02e-19
C2041 _45_/a_27_47# _09_ 0.00823f
C2042 net15 p[14] 0.00328f
C2043 _27_/a_27_297# net7 1.22e-19
C2044 _09_ _23_ 0.207f
C2045 net13 _25_ 0.00297f
C2046 _02_ _29_/a_29_53# 6.76e-21
C2047 th04_0/m1_892_n998# _30_/a_215_297# 6.06e-21
C2048 th08_0/m1_477_n803# net12 1.46e-19
C2049 p[4] net12 5.75e-19
C2050 _44_/a_250_297# b[3] 3.45e-19
C2051 _04_ _35_/a_226_47# 0.00551f
C2052 _02_ _06_ 0.85f
C2053 net10 b[1] 0.117f
C2054 _17_ _16_ 0.242f
C2055 _04_ _07_ 9.74e-20
C2056 net1 _49_/a_75_199# 0.00799f
C2057 b[1] _10_ 2.37e-20
C2058 _05_ p[2] 5.07e-19
C2059 net2 p[9] 0.00112f
C2060 VPWR _52_/a_93_21# -0.00838f
C2061 net1 input5/a_558_47# 1.1e-19
C2062 p[13] input14/a_27_47# 3.88e-19
C2063 th03_0/m1_890_n844# th15_0/Vin 4.95e-20
C2064 p[10] net5 5.12e-21
C2065 _36_/a_27_47# net13 0.0488f
C2066 net2 _15_ 9.8e-19
C2067 p[14] _06_ 2.49e-19
C2068 _43_/a_193_413# _00_ 0.00721f
C2069 net10 _48_/a_27_47# 0.00377f
C2070 _26_/a_29_53# _15_ 0.00192f
C2071 net4 _55_/a_80_21# 1.06e-19
C2072 _10_ _48_/a_27_47# 4.55e-19
C2073 Vin th09_0/m1_962_372# 0.00142f
C2074 _01_ net7 0.233f
C2075 _05_ _30_/a_109_53# 0.033f
C2076 _52_/a_250_297# net6 0.00133f
C2077 _31_/a_285_47# net7 0.00132f
C2078 _45_/a_193_297# _39_/a_47_47# 1.4e-20
C2079 net14 _50_/a_615_93# 1.69e-20
C2080 VPWR b[0] 0.166f
C2081 p[6] _34_/a_129_47# 2.45e-20
C2082 _44_/a_250_297# VGND -0.00591f
C2083 _03_ _54_/a_75_212# 5.45e-21
C2084 p[7] _09_ 1.85e-20
C2085 input5/a_62_47# output17/a_27_47# 1.02e-19
C2086 net1 input5/a_62_47# 7.59e-20
C2087 p[6] th07_0/m1_808_n892# 0.0192f
C2088 VPWR net14 0.182f
C2089 input2/a_27_47# _15_ 3.18e-20
C2090 VPWR _31_/a_285_297# 0.013f
C2091 p[3] _29_/a_29_53# 4.58e-19
C2092 th09_0/m1_485_n505# p[11] 1.22e-20
C2093 VPWR th04_0/m1_892_n998# 0.0709f
C2094 p[0] input7/a_27_47# 5.13e-20
C2095 VGND _42_/a_368_53# -4.05e-19
C2096 p[3] _06_ 3.66e-20
C2097 _43_/a_469_47# th15_0/Vin 2.09e-19
C2098 net15 net13 8.84e-19
C2099 _52_/a_93_21# b[2] 1.63e-19
C2100 th11_0/m1_705_187# output17/a_27_47# 0.00103f
C2101 th11_0/m1_705_187# net1 5.27e-20
C2102 _12_ _35_/a_76_199# 6.84e-20
C2103 VPWR _35_/a_489_413# -0.00725f
C2104 _21_ net7 3e-19
C2105 _00_ _15_ 0.207f
C2106 _03_ _30_/a_465_297# 7.72e-19
C2107 net13 _29_/a_29_53# 0.00104f
C2108 _20_ net12 0.00437f
C2109 _40_/a_109_297# VGND -0.00181f
C2110 _02_ _39_/a_285_47# 0.0019f
C2111 _19_ _09_ 4.8e-21
C2112 net13 _06_ 0.0758f
C2113 VPWR input8/a_27_47# 0.0863f
C2114 net4 net16 0.155f
C2115 net19 p[11] 0.00647f
C2116 b[2] b[0] 0.183f
C2117 net4 net10 8.28e-22
C2118 net4 _10_ 0.183f
C2119 _47_/a_81_21# th15_0/Vin 6.76e-20
C2120 _13_ _00_ 3.77e-20
C2121 _12_ net5 0.983f
C2122 _32_/a_303_47# _01_ 8.58e-19
C2123 net10 _33_/a_109_93# 0.0336f
C2124 _45_/a_193_297# _02_ 0.00988f
C2125 _24_ _09_ 0.0202f
C2126 net4 _18_ 0.023f
C2127 _04_ _20_ 0.0677f
C2128 net1 net9 0.47f
C2129 p[13] net5 0.012f
C2130 _21_ net6 2.92e-20
C2131 _20_ th15_0/m1_849_n157# 2.76e-21
C2132 net11 net7 1.77e-19
C2133 _01_ _55_/a_80_21# 0.0121f
C2134 net14 _55_/a_217_297# 2.1e-19
C2135 p[10] VGND 0.388f
C2136 _13_ output16/a_27_47# 4.58e-19
C2137 b[1] _33_/a_209_311# 0.0129f
C2138 _34_/a_377_297# _06_ 0.00427f
C2139 net9 input5/a_841_47# 2.7e-19
C2140 net7 p[1] 0.00514f
C2141 _49_/a_544_297# VGND -0.00256f
C2142 VPWR _16_ 0.126f
C2143 VPWR _29_/a_111_297# -5.85e-19
C2144 net10 _52_/a_250_297# 2.86e-21
C2145 b[1] p[11] 2.45e-20
C2146 Vin p[6] 0.353f
C2147 _10_ _52_/a_250_297# 0.00368f
C2148 _18_ _52_/a_250_297# 1.77e-19
C2149 _08_ _03_ 0.0144f
C2150 _21_ input9/a_75_212# 1.17e-21
C2151 net11 net6 1.08e-19
C2152 net8 output17/a_27_47# 0.0043f
C2153 output18/a_27_47# _21_ 0.00103f
C2154 net3 net1 4.25e-20
C2155 _45_/a_205_47# _12_ 7.46e-19
C2156 net1 net8 0.381f
C2157 net3 output17/a_27_47# 0.00248f
C2158 _02_ _50_/a_27_47# 2.09e-19
C2159 VGND _38_/a_303_47# 1.78e-19
C2160 output19/a_27_47# net15 6.88e-19
C2161 b[1] _52_/a_256_47# 8.49e-20
C2162 net16 th13_0/m1_559_n458# 6.79e-20
C2163 _27_/a_109_297# b[1] 8.35e-20
C2164 th15_0/m1_849_n157# _50_/a_343_93# 2.76e-21
C2165 p[13] th12_0/m1_529_n42# 3.34e-20
C2166 _35_/a_226_47# net1 1.3e-20
C2167 _01_ _10_ 2.22e-19
C2168 net1 _07_ 6.08e-22
C2169 _44_/a_256_47# _14_ 0.00124f
C2170 net8 input5/a_841_47# 0.025f
C2171 net15 input5/a_381_47# 7.15e-19
C2172 _18_ _01_ 6.1e-20
C2173 output19/a_27_47# _06_ 1.53e-19
C2174 _12_ _41_/a_59_75# 0.00101f
C2175 _32_/a_27_47# _30_/a_109_53# 1.51e-19
C2176 _36_/a_303_47# net5 0.00256f
C2177 _03_ _39_/a_47_47# 1.47e-19
C2178 _35_/a_226_297# net10 2.48e-19
C2179 _11_ net9 5.39e-19
C2180 _12_ VGND 0.816f
C2181 net11 input9/a_75_212# 1.1e-20
C2182 _55_/a_217_297# _16_ 0.0017f
C2183 net19 _42_/a_209_311# 0.0766f
C2184 net11 output18/a_27_47# 6.84e-20
C2185 input15/a_27_47# net15 0.00325f
C2186 net15 th14_0/m1_891_419# 3.54e-21
C2187 input5/a_381_47# _06_ 1.6e-19
C2188 _34_/a_47_47# input12/a_27_47# 2.17e-19
C2189 p[13] VGND 0.153f
C2190 net16 _21_ 1.89e-19
C2191 _26_/a_29_53# _36_/a_27_47# 1.6e-19
C2192 _26_/a_183_297# _00_ 4.53e-19
C2193 _49_/a_315_47# p[2] 8.45e-20
C2194 net8 _37_/a_27_47# 6.66e-21
C2195 net10 _21_ 0.0275f
C2196 net3 _37_/a_27_47# 0.094f
C2197 _17_ net19 0.0269f
C2198 net15 _37_/a_197_47# 1.78e-19
C2199 p[8] p[11] 0.00322f
C2200 _10_ _21_ 0.00421f
C2201 _40_/a_191_297# _14_ 2.4e-19
C2202 _03_ _49_/a_208_47# 3.86e-19
C2203 input15/a_27_47# _06_ 4.73e-19
C2204 _12_ _50_/a_223_47# 0.00327f
C2205 _35_/a_556_47# b[1] 3.23e-19
C2206 _30_/a_392_297# net9 9.92e-19
C2207 _54_/a_75_212# net18 0.0143f
C2208 VPWR _50_/a_429_93# -3.61e-19
C2209 _20_ _55_/a_472_297# 0.00212f
C2210 net13 _50_/a_27_47# 7.27e-21
C2211 p[14] input6/a_27_47# 0.0235f
C2212 _05_ Vin 8.25e-21
C2213 th07_0/m1_808_n892# input11/a_27_47# 1.85e-20
C2214 net15 net2 0.324f
C2215 _22_ net12 5.73e-20
C2216 _13_ _45_/a_27_47# 0.0703f
C2217 net8 _11_ 1.81e-20
C2218 net3 _11_ 0.165f
C2219 input10/a_27_47# _54_/a_75_212# 1.17e-22
C2220 net6 _50_/a_515_93# 4.7e-19
C2221 net16 net11 4.43e-22
C2222 VPWR input13/a_27_47# 0.0699f
C2223 b[1] _42_/a_209_311# 5.21e-19
C2224 _43_/a_27_47# _32_/a_27_47# 2.01e-20
C2225 _34_/a_47_47# VGND 0.0892f
C2226 _26_/a_29_53# net15 9.06e-21
C2227 _03_ _02_ 0.00474f
C2228 _13_ _23_ 2.08e-20
C2229 net11 net10 0.592f
C2230 net11 _10_ 0.0109f
C2231 net2 _06_ 0.0108f
C2232 _43_/a_193_413# _19_ 4.85e-21
C2233 _19_ _49_/a_315_47# 1.33e-19
C2234 VGND _55_/a_300_47# -0.00109f
C2235 _47_/a_81_21# th15_0/m1_849_n157# 4.9e-19
C2236 p[7] _34_/a_285_47# 5.01e-20
C2237 _26_/a_29_53# _29_/a_29_53# 0.00121f
C2238 _26_/a_29_53# _06_ 0.0135f
C2239 _02_ _14_ 0.0316f
C2240 _04_ _22_ 1.76e-20
C2241 net15 input2/a_27_47# 1.61e-19
C2242 _20_ net1 0.363f
C2243 _48_/a_109_47# _06_ 9.47e-19
C2244 p[14] _14_ 1.13e-19
C2245 _55_/a_80_21# net7 0.00163f
C2246 _36_/a_303_47# VGND 8.14e-19
C2247 _44_/a_250_297# input5/a_62_47# 2.45e-20
C2248 _52_/a_93_21# _52_/a_346_47# -5.12e-20
C2249 _00_ net15 0.00147f
C2250 _27_/a_27_297# _27_/a_109_297# -3.68e-20
C2251 _03_ p[3] 0.00387f
C2252 p[10] net17 0.183f
C2253 input7/a_27_47# input5/a_664_47# 1.08e-21
C2254 VPWR th09_0/m1_485_n505# 0.0937f
C2255 _00_ _06_ 0.1f
C2256 _19_ _15_ 1.46e-20
C2257 VPWR _47_/a_299_297# 0.0643f
C2258 Vin input11/a_27_47# 0.00547f
C2259 _03_ net13 0.271f
C2260 p[10] input5/a_558_47# 1.09e-19
C2261 net14 th15_0/Vin 0.0111f
C2262 th02_0/m1_571_144# p[1] 1.08e-20
C2263 _27_/a_277_297# net8 7.99e-20
C2264 _27_/a_205_297# net14 3.63e-19
C2265 _27_/a_277_297# net3 2.71e-19
C2266 b[1] _30_/a_215_297# 0.0176f
C2267 VPWR net19 0.189f
C2268 net10 net7 1.65e-36
C2269 net4 _17_ 7.52e-21
C2270 VPWR input1/a_75_212# 0.0788f
C2271 _10_ net7 6.22e-20
C2272 net1 th03_0/m1_890_n844# 2.78e-20
C2273 _13_ _24_ 2.47e-19
C2274 _43_/a_27_47# _15_ 8.96e-20
C2275 _42_/a_109_93# p[11] 3.74e-19
C2276 _10_ _50_/a_515_93# 0.00129f
C2277 _18_ net7 2.58e-20
C2278 th14_0/m1_641_n318# th11_0/m1_577_n654# 2.63e-20
C2279 _29_/a_183_297# _04_ 0.0015f
C2280 VGND _37_/a_109_47# -7.9e-19
C2281 _20_ _11_ 0.268f
C2282 _43_/a_27_47# _13_ 1.66e-20
C2283 _03_ _34_/a_377_297# 3.13e-20
C2284 net11 _33_/a_209_311# 2.49e-19
C2285 net16 net6 8.27e-20
C2286 p[10] th11_0/m1_705_187# 0.0622f
C2287 net10 net6 1.35e-20
C2288 _02_ input5/a_664_47# 0.00187f
C2289 _27_/a_27_297# _42_/a_209_311# 4.7e-20
C2290 _10_ net6 0.0965f
C2291 _00_ _39_/a_285_47# 1.47e-21
C2292 _18_ net6 0.166f
C2293 VPWR b[1] 1.11f
C2294 _53_/a_29_53# _11_ 2.33e-20
C2295 p[6] input11/a_27_47# 7.64e-20
C2296 p[13] net17 8.11e-20
C2297 _44_/a_93_21# net14 0.0646f
C2298 _44_/a_250_297# net3 0.0088f
C2299 _23_ _25_ 0.00465f
C2300 _17_ _27_/a_27_297# 6.78e-22
C2301 output19/a_27_47# input6/a_27_47# 0.107f
C2302 _35_/a_76_199# _08_ 0.0061f
C2303 _00_ _45_/a_193_297# 4.38e-20
C2304 _49_/a_201_297# net13 3.31e-19
C2305 _23_ _36_/a_27_47# 0.00118f
C2306 th15_0/Vin _16_ 5.12e-19
C2307 VPWR _48_/a_27_47# 0.0158f
C2308 p[13] _49_/a_75_199# 1.23e-19
C2309 _01_ _42_/a_209_311# 1.58e-19
C2310 net3 _42_/a_368_53# 3.82e-19
C2311 net14 _42_/a_296_53# 2.18e-19
C2312 p[13] input5/a_558_47# 0.00363f
C2313 net16 output18/a_27_47# 3.45e-19
C2314 _11_ _50_/a_343_93# 0.0384f
C2315 net10 input9/a_75_212# 0.00699f
C2316 _09_ _05_ 0.0683f
C2317 _47_/a_81_21# net1 1.58e-21
C2318 _26_/a_29_53# _50_/a_27_47# 5.56e-19
C2319 _10_ input9/a_75_212# 5.49e-21
C2320 _33_/a_109_93# _30_/a_215_297# 0.00104f
C2321 VGND _54_/a_75_212# 0.053f
C2322 _35_/a_556_47# _21_ 2.69e-19
C2323 _10_ _55_/a_80_21# 5.49e-19
C2324 _17_ _01_ 1.46e-20
C2325 net4 _38_/a_109_47# 7.32e-19
C2326 net15 _40_/a_297_297# 4.08e-19
C2327 net3 _40_/a_109_297# 3.14e-19
C2328 _02_ net18 8.53e-20
C2329 _18_ _55_/a_80_21# 1.44e-20
C2330 input15/a_27_47# input6/a_27_47# 5.3e-19
C2331 b[1] b[2] 5.48e-19
C2332 _47_/a_384_47# _10_ 3.53e-19
C2333 net1 _22_ 0.0129f
C2334 input3/a_27_47# output19/a_27_47# 4.77e-21
C2335 _39_/a_377_297# _06_ 8.76e-20
C2336 output19/a_27_47# _14_ 1.43e-19
C2337 th09_0/m1_962_372# p[9] 5.57e-19
C2338 _04_ _52_/a_93_21# 2.35e-19
C2339 p[13] input5/a_62_47# 0.0281f
C2340 _40_/a_297_297# _06_ 1.64e-19
C2341 VGND _30_/a_465_297# 6.42e-19
C2342 _14_ input5/a_381_47# 5.68e-20
C2343 th04_0/m1_892_n998# net12 1.19e-21
C2344 _45_/a_27_47# _06_ 0.0021f
C2345 _00_ _50_/a_27_47# 0.00197f
C2346 p[13] th11_0/m1_705_187# 0.0061f
C2347 VPWR p[8] 0.267f
C2348 net4 VPWR 1.07f
C2349 net2 input6/a_27_47# 0.0047f
C2350 p[10] net8 0.00619f
C2351 _39_/a_47_47# net5 0.0389f
C2352 _23_ _06_ 0.218f
C2353 p[10] net3 3.61e-19
C2354 _31_/a_117_297# p[10] 1.09e-19
C2355 VPWR _33_/a_109_93# -0.00817f
C2356 net16 _10_ 0.0338f
C2357 _44_/a_93_21# _16_ 0.00354f
C2358 _17_ _42_/a_109_93# 7.83e-20
C2359 input3/a_27_47# th14_0/m1_891_419# 3.77e-20
C2360 Vin p[9] 0.112f
C2361 _35_/a_489_413# net12 3.97e-20
C2362 _45_/a_109_297# _05_ 2.79e-22
C2363 input15/a_27_47# _14_ 9.48e-21
C2364 net16 _18_ 8.17e-21
C2365 net10 _10_ 4.45e-19
C2366 net10 _18_ 1.47e-21
C2367 _31_/a_35_297# _02_ 0.00316f
C2368 _04_ net14 0.0863f
C2369 _18_ _10_ 0.133f
C2370 _04_ th04_0/m1_892_n998# 4.5e-20
C2371 _12_ net9 4.39e-22
C2372 _03_ net2 1.89e-19
C2373 p[13] net9 1.72e-19
C2374 net4 p[12] 0.0242f
C2375 _35_/a_76_199# _02_ 5.73e-19
C2376 VPWR _48_/a_181_47# -3.35e-19
C2377 _47_/a_81_21# _11_ 0.0454f
C2378 input3/a_27_47# net2 0.0229f
C2379 _26_/a_29_53# _03_ 7.93e-21
C2380 VPWR _52_/a_250_297# 0.019f
C2381 p[7] _06_ 0.00878f
C2382 _30_/a_109_53# _29_/a_29_53# 0.0103f
C2383 _04_ input8/a_27_47# 2.36e-22
C2384 net2 _14_ 0.0104f
C2385 VPWR _27_/a_27_297# 0.0329f
C2386 _30_/a_109_53# _06_ 1.96e-19
C2387 _43_/a_297_47# _00_ 1.26e-19
C2388 _11_ _22_ 0.15f
C2389 _08_ VGND 0.161f
C2390 _19_ net15 0.00628f
C2391 _02_ net5 0.233f
C2392 net4 _55_/a_217_297# 1.13e-19
C2393 _26_/a_29_53# _14_ 3.67e-19
C2394 _03_ input2/a_27_47# 2.71e-19
C2395 _21_ _30_/a_215_297# 1.48e-19
C2396 p[7] th05_0/m1_752_n794# 2.37e-19
C2397 _44_/a_256_47# VGND -0.00184f
C2398 _29_/a_111_297# net12 1.21e-19
C2399 _28_/a_109_297# _55_/a_80_21# 2.05e-20
C2400 p[6] _34_/a_285_47# 4.63e-19
C2401 _39_/a_285_47# _23_ 1.9e-20
C2402 _20_ _40_/a_109_297# 2.35e-20
C2403 _12_ net3 3.09e-20
C2404 th12_0/m1_394_n856# Vin 8.07e-19
C2405 _55_/a_80_21# p[11] 9.25e-20
C2406 _34_/a_47_47# net9 1.41e-20
C2407 VPWR th13_0/m1_559_n458# 0.0186f
C2408 _52_/a_250_297# p[12] 1.84e-20
C2409 VPWR _01_ 0.521f
C2410 _24_ _53_/a_111_297# 9.08e-21
C2411 VPWR _31_/a_285_47# -2.91e-19
C2412 _05_ _32_/a_27_47# 2.2e-20
C2413 _35_/a_76_199# p[3] 2.23e-19
C2414 _00_ _03_ 2.31e-20
C2415 p[13] net8 0.00375f
C2416 p[13] net3 9.08e-19
C2417 VGND input7/a_27_47# 0.0575f
C2418 _32_/a_109_47# net5 5.69e-21
C2419 _31_/a_35_297# net13 1.86e-20
C2420 net4 input4/a_75_212# 0.0178f
C2421 _52_/a_250_297# b[2] 1.6e-19
C2422 _45_/a_193_297# _23_ 4.13e-19
C2423 _12_ _35_/a_226_47# 8.38e-20
C2424 _24_ _06_ 0.113f
C2425 _12_ _07_ 2.94e-23
C2426 _04_ _29_/a_111_297# 9.25e-19
C2427 _39_/a_47_47# VGND 0.0665f
C2428 VPWR _35_/a_226_297# -8.54e-19
C2429 _00_ _14_ 0.133f
C2430 _40_/a_191_297# VGND -9.29e-19
C2431 _35_/a_76_199# net13 0.0337f
C2432 net11 _30_/a_215_297# 1.04e-19
C2433 _43_/a_27_47# _06_ 0.0329f
C2434 _02_ input12/a_27_47# 1.88e-19
C2435 th09_0/m1_485_n505# th15_0/Vin 0.00438f
C2436 th13_0/m1_559_n458# p[12] 2.29e-19
C2437 VPWR _21_ 0.869f
C2438 _47_/a_299_297# th15_0/Vin 8.81e-20
C2439 th14_0/m1_891_419# input5/a_664_47# 2.08e-20
C2440 net10 _33_/a_209_311# 0.0426f
C2441 _49_/a_208_47# VGND -0.00164f
C2442 VPWR _42_/a_109_93# -0.00115f
C2443 _28_/a_109_297# _10_ 4.34e-19
C2444 net13 net5 0.127f
C2445 _10_ p[11] 9.81e-21
C2446 VGND th11_0/m1_577_n654# 0.0025f
C2447 p[14] b[3] 0.0451f
C2448 _52_/a_584_47# _22_ 6.24e-19
C2449 th15_0/Vin net19 0.00574f
C2450 _18_ p[11] 1.24e-19
C2451 _09_ _49_/a_315_47# 1.11e-20
C2452 _45_/a_27_47# _50_/a_27_47# 0.109f
C2453 _01_ _55_/a_217_297# 0.00112f
C2454 input1/a_75_212# th15_0/Vin 0.00156f
C2455 net6 _42_/a_209_311# 1.32e-20
C2456 output19/a_27_47# input14/a_27_47# 0.0101f
C2457 _34_/a_47_47# _07_ 0.011f
C2458 b[1] _33_/a_296_53# 2.69e-20
C2459 _34_/a_129_47# _06_ 5.3e-19
C2460 th14_0/m1_641_n318# net2 4.8e-19
C2461 net2 input5/a_664_47# 8.11e-20
C2462 _02_ VGND 1.63f
C2463 VPWR net11 1f
C2464 net10 _52_/a_256_47# 8.13e-20
C2465 _17_ net6 3.12e-19
C2466 p[14] _41_/a_59_75# 5.52e-19
C2467 _10_ _52_/a_256_47# 1.65e-19
C2468 _05_ _34_/a_285_47# 7.85e-21
C2469 _21_ b[2] 2.14e-19
C2470 VGND p[14] 0.619f
C2471 th01_0/m1_991_n1219# p[1] 5.78e-20
C2472 p[0] th02_0/m1_983_133# 0.0563f
C2473 VPWR p[1] 0.135f
C2474 th08_0/m1_477_n803# _34_/a_47_47# 3.25e-20
C2475 input13/a_27_47# net12 0.0163f
C2476 _45_/a_465_47# _12_ 0.00211f
C2477 net14 net1 6.64e-20
C2478 _31_/a_285_297# net1 5.85e-19
C2479 _02_ _50_/a_223_47# 2.51e-20
C2480 _32_/a_109_47# VGND 1.05e-19
C2481 _12_ _20_ 3.9e-19
C2482 _55_/a_80_21# _42_/a_209_311# 0.0175f
C2483 b[1] _52_/a_346_47# 6.37e-20
C2484 b[1] th15_0/Vin 7.03e-19
C2485 input2/a_27_47# input5/a_664_47# 4.47e-21
C2486 _27_/a_205_297# b[1] 1.41e-19
C2487 _13_ _05_ 2.57e-20
C2488 _02_ _53_/a_183_297# 4.14e-19
C2489 _44_/a_93_21# net19 0.0074f
C2490 _44_/a_346_47# _14_ 3.76e-19
C2491 _17_ _55_/a_80_21# 7.64e-21
C2492 _11_ _38_/a_27_47# 0.071f
C2493 net11 b[2] 1.46e-19
C2494 p[3] VGND 0.526f
C2495 _13_ _09_ 0.0927f
C2496 net1 input8/a_27_47# 0.0347f
C2497 _35_/a_556_47# net10 5.59e-19
C2498 net4 th15_0/m1_597_n912# 2.43e-20
C2499 _12_ _53_/a_29_53# 3.46e-20
C2500 _17_ _47_/a_384_47# 1.1e-20
C2501 net2 input14/a_27_47# 0.0235f
C2502 _26_/a_29_53# net18 2.57e-21
C2503 _55_/a_472_297# _16_ 3.71e-19
C2504 net19 _42_/a_296_53# 2.71e-19
C2505 Vin net15 0.0041f
C2506 VGND net13 0.142f
C2507 _30_/a_215_297# net6 3.3e-21
C2508 _45_/a_27_47# _03_ 2.06e-20
C2509 net14 _37_/a_27_47# 0.0584f
C2510 net15 _37_/a_303_47# 0.00118f
C2511 net3 _37_/a_109_47# 0.00212f
C2512 _40_/a_297_297# _14_ 1.58e-19
C2513 Vin _29_/a_29_53# 1.71e-21
C2514 _03_ _23_ 0.0564f
C2515 _12_ _50_/a_343_93# 5.63e-20
C2516 Vin _06_ 0.00141f
C2517 VPWR net7 0.786f
C2518 th10_0/m1_536_174# b[3] 0.00833f
C2519 net5 input5/a_381_47# 0.0546f
C2520 p[5] net13 1.05e-19
C2521 VPWR _50_/a_515_93# -5.03e-19
C2522 _18_ _42_/a_209_311# 3.21e-19
C2523 _31_/a_35_297# net2 0.0635f
C2524 _17_ _10_ 0.0233f
C2525 p[8] th15_0/Vin 0.167f
C2526 _17_ _18_ 0.271f
C2527 th14_0/m1_891_419# net5 0.00243f
C2528 Vin th05_0/m1_752_n794# 0.117f
C2529 _03_ p[2] 2.16e-20
C2530 net4 th15_0/Vin 3.6e-19
C2531 input9/a_75_212# _30_/a_215_297# 6.24e-21
C2532 th04_0/m1_620_n488# p[1] 1.03e-21
C2533 net6 _50_/a_615_93# 1.43e-19
C2534 net14 _11_ 5e-19
C2535 _34_/a_47_47# _53_/a_29_53# 5.88e-22
C2536 _34_/a_377_297# VGND -0.00102f
C2537 net17 input7/a_27_47# 4.99e-20
C2538 b[1] _42_/a_296_53# 2.38e-20
C2539 _30_/a_465_297# net9 0.00138f
C2540 VGND th10_0/m1_536_174# 0.0658f
C2541 p[7] _03_ 4.51e-22
C2542 input5/a_841_47# _16_ 8.62e-19
C2543 VPWR net6 0.999f
C2544 _03_ _30_/a_109_53# 0.0189f
C2545 _26_/a_111_297# _06_ 9e-19
C2546 input7/a_27_47# input5/a_558_47# 1.22e-20
C2547 _04_ net19 2.07e-20
C2548 _31_/a_35_297# input2/a_27_47# 0.00136f
C2549 output19/a_27_47# b[3] 0.0274f
C2550 net2 net5 0.0616f
C2551 VPWR _32_/a_303_47# 6.03e-19
C2552 _55_/a_217_297# net7 1.04e-19
C2553 p[6] _06_ 0.00365f
C2554 _37_/a_27_47# _16_ 2.07e-19
C2555 _26_/a_29_53# net5 0.0237f
C2556 _19_ _03_ 0.0019f
C2557 p[12] net6 0.0439f
C2558 b[1] net12 0.12f
C2559 VPWR input9/a_75_212# 0.0643f
C2560 VPWR _55_/a_80_21# 0.0289f
C2561 _32_/a_27_47# _15_ 1.19e-19
C2562 VPWR output18/a_27_47# 0.0689f
C2563 net10 _30_/a_215_297# 0.0512f
C2564 _10_ _30_/a_215_297# 5.66e-20
C2565 output19/a_27_47# VGND 0.0024f
C2566 _12_ _47_/a_81_21# 0.00158f
C2567 input15/a_27_47# b[3] 1.77e-19
C2568 _24_ _03_ 9.46e-20
C2569 _19_ _14_ 2.71e-21
C2570 net16 _38_/a_109_47# 4.17e-19
C2571 p[6] th05_0/m1_752_n794# 0.00131f
C2572 VPWR _47_/a_384_47# -1.45e-19
C2573 th14_0/m1_891_419# th12_0/m1_529_n42# 0.00211f
C2574 _48_/a_27_47# net12 0.0126f
C2575 th11_0/m1_705_187# input7/a_27_47# 1.5e-20
C2576 _02_ net17 0.0608f
C2577 _04_ b[1] 0.0568f
C2578 _10_ _38_/a_109_47# 5.44e-19
C2579 VGND input5/a_381_47# -0.00305f
C2580 _49_/a_201_297# p[2] 8.68e-20
C2581 _11_ _16_ 4.42e-20
C2582 _05_ _36_/a_27_47# 3.67e-21
C2583 th15_0/Vin th13_0/m1_559_n458# 1.16e-21
C2584 _09_ _25_ 1.49e-19
C2585 _08_ net9 7.71e-21
C2586 _12_ _22_ 0.196f
C2587 _27_/a_277_297# net14 5.1e-19
C2588 _00_ net5 0.00954f
C2589 input15/a_27_47# _41_/a_59_75# 3.96e-20
C2590 _02_ _49_/a_75_199# 0.0354f
C2591 _43_/a_193_413# p[9] 1.09e-19
C2592 Vin p[0] 0.134f
C2593 input15/a_27_47# VGND 0.0158f
C2594 th14_0/m1_891_419# VGND 0.00531f
C2595 net2 b[3] 0.00419f
C2596 _43_/a_27_47# _14_ 0.00938f
C2597 _43_/a_193_413# _15_ 4.86e-19
C2598 _42_/a_209_311# p[11] 4.19e-19
C2599 _10_ _50_/a_615_93# 8.82e-19
C2600 net1 input13/a_27_47# 1.9e-19
C2601 output18/a_27_47# b[2] 0.0141f
C2602 VPWR net16 0.518f
C2603 net2 th12_0/m1_529_n42# 0.0122f
C2604 net6 input4/a_75_212# 0.0271f
C2605 VGND _37_/a_197_47# -4.58e-19
C2606 VPWR net10 0.375f
C2607 VPWR _10_ 0.577f
C2608 _17_ p[11] 0.00765f
C2609 _43_/a_193_413# _13_ 5.58e-21
C2610 net5 output16/a_27_47# 4.14e-19
C2611 _55_/a_80_21# _55_/a_217_297# 1.42e-32
C2612 VPWR _18_ 0.0721f
C2613 th11_0/m1_705_187# th11_0/m1_577_n654# -1.6e-19
C2614 th15_0/Vin _42_/a_109_93# 9.71e-20
C2615 net4 net12 2.57e-20
C2616 net2 VGND 0.852f
C2617 _33_/a_109_93# net12 0.0435f
C2618 _05_ _29_/a_29_53# 3.79e-20
C2619 _34_/a_47_47# _22_ 3.9e-21
C2620 _05_ _06_ 0.00724f
C2621 _09_ _53_/a_111_297# 3.4e-19
C2622 _26_/a_29_53# VGND 0.0381f
C2623 _15_ p[9] 2.06e-19
C2624 _44_/a_256_47# net3 0.00101f
C2625 _44_/a_250_297# net14 4.24e-20
C2626 _23_ net18 -4.05e-24
C2627 net17 net13 5.21e-20
C2628 input9/a_75_212# th04_0/m1_620_n488# 8.03e-20
C2629 _10_ p[12] 0.0134f
C2630 _48_/a_109_47# VGND 9.44e-19
C2631 _55_/a_300_47# _22_ 2.08e-19
C2632 _09_ _29_/a_29_53# 0.00488f
C2633 _35_/a_226_47# _08_ 0.00117f
C2634 _18_ p[12] 2.17e-19
C2635 _09_ _06_ 0.0965f
C2636 _08_ _07_ 0.348f
C2637 _04_ _33_/a_109_93# 0.0299f
C2638 net13 _49_/a_75_199# 3.2e-19
C2639 net8 input7/a_27_47# 2.03e-21
C2640 net14 _42_/a_368_53# 7.39e-19
C2641 _13_ _15_ 3.69e-20
C2642 input2/a_27_47# VGND -0.0137f
C2643 _26_/a_29_53# _50_/a_223_47# 0.00124f
C2644 VPWR th02_0/m1_571_144# 0.0143f
C2645 _19_ input5/a_664_47# 2.19e-21
C2646 _33_/a_209_311# _30_/a_215_297# 1.56e-19
C2647 th01_0/m1_991_n1219# th02_0/m1_571_144# 0.00603f
C2648 th01_0/m1_571_n501# th02_0/m1_983_133# 7.11e-20
C2649 th15_0/Vin p[1] 2.84e-19
C2650 _10_ _55_/a_217_297# 1.43e-19
C2651 net3 _39_/a_47_47# 1.66e-20
C2652 net4 _38_/a_197_47# 7.64e-19
C2653 _00_ _41_/a_59_75# 2.43e-20
C2654 net3 _40_/a_191_297# 1.89e-19
C2655 Vin input6/a_27_47# 0.00242f
C2656 _02_ net9 0.00611f
C2657 th03_0/m1_638_n591# VGND 0.00103f
C2658 _00_ VGND 0.139f
C2659 _44_/a_93_21# _42_/a_109_93# 1.25e-19
C2660 input1/a_75_212# output17/a_27_47# 0.0101f
C2661 input1/a_75_212# net1 0.00208f
C2662 _49_/a_208_47# net8 1.4e-19
C2663 _04_ _52_/a_250_297# 3.98e-21
C2664 _04_ _27_/a_27_297# 0.0526f
C2665 _10_ input4/a_75_212# 0.00346f
C2666 _32_/a_109_47# net9 6.44e-19
C2667 _01_ net12 1.67e-21
C2668 _18_ input4/a_75_212# 4.36e-19
C2669 th12_0/m1_394_n856# p[9] 1.33e-19
C2670 _45_/a_27_47# _35_/a_76_199# 2.04e-21
C2671 p[7] input10/a_27_47# 3.04e-19
C2672 _03_ Vin 5.94e-19
C2673 VGND output16/a_27_47# 0.0728f
C2674 _45_/a_109_297# _06_ 0.0023f
C2675 _00_ _50_/a_223_47# 0.00738f
C2676 p[10] net14 1.59e-20
C2677 _39_/a_377_297# net5 0.00234f
C2678 _32_/a_197_47# _01_ 0.00156f
C2679 _31_/a_285_297# p[10] 4.45e-20
C2680 VPWR _33_/a_209_311# -0.0131f
C2681 _17_ _42_/a_209_311# 1.22e-19
C2682 _44_/a_250_297# _16_ 3.25e-19
C2683 _32_/a_27_47# _36_/a_27_47# 0.011f
C2684 VPWR _28_/a_109_297# -1.71e-19
C2685 th09_0/m1_485_n505# th10_0/m1_502_n495# 7.17e-20
C2686 _45_/a_193_297# _05_ 4.84e-22
C2687 _31_/a_35_297# p[2] 0.00277f
C2688 Vin _14_ 3.46e-19
C2689 _12_ _38_/a_27_47# 0.0527f
C2690 th15_0/m1_597_n912# net6 1.34e-20
C2691 p[3] net9 0.0376f
C2692 VPWR p[11] 0.401f
C2693 _02_ net8 0.334f
C2694 net3 _02_ 9.52e-20
C2695 _45_/a_27_47# net5 0.0288f
C2696 _04_ _01_ 0.119f
C2697 _24_ net18 5.57e-21
C2698 b[1] output17/a_27_47# 0.0373f
C2699 b[1] net1 0.0593f
C2700 _37_/a_27_47# net19 0.0105f
C2701 _45_/a_193_297# _09_ 0.00961f
C2702 th15_0/Vin net7 1.02e-19
C2703 _23_ net5 0.0052f
C2704 input11/a_27_47# th05_0/m1_752_n794# 2.38e-19
C2705 net3 p[14] 0.00504f
C2706 _21_ net12 0.23f
C2707 _31_/a_35_297# _30_/a_109_53# 2.89e-20
C2708 th06_0/m1_904_n796# th07_0/m1_808_n892# 2.38e-19
C2709 _35_/a_226_47# _02_ 2.21e-19
C2710 net13 net9 0.035f
C2711 _04_ _35_/a_226_297# 4.51e-19
C2712 _02_ _07_ 0.0083f
C2713 _12_ _52_/a_93_21# 0.0157f
C2714 _47_/a_299_297# _11_ 0.00738f
C2715 _32_/a_109_47# net8 0.0011f
C2716 VPWR _52_/a_256_47# -9.47e-19
C2717 net17 input5/a_381_47# 1.37e-20
C2718 b[1] input5/a_841_47# 7.07e-19
C2719 VPWR _27_/a_109_297# -2.45e-19
C2720 _11_ net19 2.19e-19
C2721 _04_ _21_ 0.39f
C2722 _19_ _31_/a_35_297# 1.47e-19
C2723 _12_ b[0] 2.61e-20
C2724 _04_ _42_/a_109_93# 5.77e-22
C2725 th15_0/Vin net6 0.00781f
C2726 p[3] net8 0.0015f
C2727 _32_/a_27_47# _06_ 0.00663f
C2728 _20_ _39_/a_47_47# 2.3e-20
C2729 _44_/a_346_47# VGND -0.00198f
C2730 net11 net12 0.358f
C2731 _30_/a_109_53# net5 5.84e-22
C2732 _20_ _40_/a_191_297# 2.07e-20
C2733 _55_/a_217_297# p[11] 1.6e-20
C2734 th14_0/m1_891_419# input5/a_558_47# 3.96e-20
C2735 _09_ _50_/a_27_47# 1.3e-19
C2736 p[13] net14 5.58e-19
C2737 net3 net13 3.25e-21
C2738 net8 net13 7.51e-20
C2739 _43_/a_193_413# net15 0.00169f
C2740 _04_ net11 0.078f
C2741 VPWR _35_/a_556_47# -7.24e-19
C2742 net17 net2 0.261f
C2743 _39_/a_377_297# VGND -6.28e-19
C2744 _19_ net5 6.41e-21
C2745 _40_/a_297_297# VGND -5.1e-19
C2746 _35_/a_226_47# net13 0.00709f
C2747 net13 _07_ 0.00686f
C2748 _04_ p[1] 9.99e-21
C2749 th08_0/m1_477_n803# p[3] 3.99e-19
C2750 _43_/a_193_413# _06_ 0.0138f
C2751 _45_/a_27_47# VGND -0.029f
C2752 th14_0/m1_641_n318# Vin 0.00276f
C2753 th06_0/m1_904_n796# Vin 0.0135f
C2754 _24_ net5 5.83e-20
C2755 net2 input5/a_558_47# 5.99e-21
C2756 th14_0/m1_891_419# input5/a_62_47# 0.00116f
C2757 p[7] input12/a_27_47# 1.65e-19
C2758 net10 _33_/a_296_53# 8.22e-20
C2759 _23_ VGND 0.16f
C2760 VPWR _42_/a_209_311# -0.00753f
C2761 _44_/a_93_21# net6 1.08e-20
C2762 _20_ _02_ 0.1f
C2763 net13 p[4] 2.34e-20
C2764 net17 input2/a_27_47# 0.0398f
C2765 th11_0/m1_705_187# th14_0/m1_891_419# 1.31e-19
C2766 b[1] _30_/a_392_297# 3.99e-19
C2767 net15 p[9] 0.00302f
C2768 VPWR _17_ 0.306f
C2769 net15 _15_ 0.156f
C2770 _01_ _55_/a_472_297# 6.28e-19
C2771 Vin th01_0/m1_571_n501# 0.00112f
C2772 _34_/a_285_47# _06_ 0.00598f
C2773 _34_/a_377_297# _07_ 5.8e-19
C2774 p[2] VGND 0.29f
C2775 p[8] _37_/a_27_47# 9.82e-21
C2776 net9 input5/a_381_47# 3.4e-19
C2777 _27_/a_27_297# net1 6.05e-21
C2778 b[1] _33_/a_368_53# 4.19e-19
C2779 net2 input5/a_62_47# 0.0197f
C2780 input2/a_27_47# input5/a_558_47# 2.04e-20
C2781 net7 net12 1.57e-19
C2782 _02_ _53_/a_29_53# 0.0388f
C2783 p[9] _06_ 0.00205f
C2784 _05_ _03_ 0.135f
C2785 _15_ _06_ 0.22f
C2786 p[8] th10_0/m1_502_n495# 1.22e-20
C2787 _10_ th15_0/Vin 0.00935f
C2788 p[14] _41_/a_145_75# 1.12e-19
C2789 p[7] VGND 0.323f
C2790 th11_0/m1_705_187# net2 1.39e-19
C2791 _18_ th15_0/Vin 6.4e-19
C2792 VGND _30_/a_109_53# -0.0072f
C2793 VGND th02_0/m1_983_133# 0.0729f
C2794 _09_ _03_ 0.326f
C2795 p[3] _20_ 7.36e-19
C2796 _13_ _06_ 0.00188f
C2797 Vin input14/a_27_47# 4.64e-19
C2798 _04_ net7 0.0602f
C2799 p[8] _11_ 6.68e-20
C2800 _01_ net1 0.0509f
C2801 p[5] p[7] 2.33e-19
C2802 _02_ _50_/a_343_93# 6.94e-19
C2803 net4 _11_ 0.0858f
C2804 th06_0/m1_904_n796# p[6] 0.00406f
C2805 output19/a_27_47# net3 0.00356f
C2806 Vin input10/a_27_47# 0.00453f
C2807 net12 net6 0.00643f
C2808 _27_/a_277_297# b[1] 1.24e-19
C2809 _20_ net13 5.95e-19
C2810 _19_ VGND 0.379f
C2811 th11_0/m1_705_187# input2/a_27_47# 3e-19
C2812 _44_/a_250_297# net19 0.00592f
C2813 net8 input5/a_381_47# 7.48e-19
C2814 net3 input5/a_381_47# 0.0299f
C2815 net2 net9 3.64e-20
C2816 VPWR _30_/a_215_297# -0.00548f
C2817 _24_ VGND -0.00863f
C2818 _26_/a_29_53# net9 0.00343f
C2819 _04_ net6 2.61e-20
C2820 net1 _21_ 0.0252f
C2821 net19 _42_/a_368_53# 5.12e-19
C2822 th15_0/Vin th02_0/m1_571_144# 8.16e-21
C2823 th14_0/m1_891_419# net8 2.46e-21
C2824 input15/a_27_47# net3 8.74e-20
C2825 net3 th14_0/m1_891_419# 2.08e-19
C2826 _31_/a_35_297# Vin 5.96e-19
C2827 VPWR _38_/a_109_47# -4.66e-19
C2828 _44_/a_93_21# _10_ 2.48e-19
C2829 _42_/a_109_93# output17/a_27_47# 8.6e-21
C2830 th15_0/m1_849_n157# net6 3.87e-20
C2831 _43_/a_27_47# VGND -0.0153f
C2832 _44_/a_93_21# _18_ 0.00485f
C2833 _54_/a_75_212# _38_/a_27_47# 2.67e-19
C2834 net14 _37_/a_109_47# 1.71e-19
C2835 net3 _37_/a_197_47# 0.0028f
C2836 _35_/a_76_199# Vin 5.98e-21
C2837 _21_ input5/a_841_47# 1.59e-21
C2838 VPWR _50_/a_615_93# -5.34e-19
C2839 p[3] th03_0/m1_890_n844# 2.56e-19
C2840 _13_ _39_/a_285_47# 0.00451f
C2841 net4 th13_0/m1_831_275# 3.27e-19
C2842 _09_ _49_/a_201_297# 1.74e-20
C2843 _04_ input9/a_75_212# 7.69e-22
C2844 _36_/a_27_47# _25_ 2.34e-20
C2845 net2 net8 0.0525f
C2846 net3 net2 0.519f
C2847 _00_ net9 0.00501f
C2848 net11 net1 1.13e-19
C2849 p[6] input10/a_27_47# 0.00459f
C2850 VPWR th01_0/m1_991_n1219# 0.0681f
C2851 b[1] _42_/a_368_53# 5.32e-20
C2852 _26_/a_29_53# net3 2.83e-21
C2853 _34_/a_129_47# VGND -8.76e-20
C2854 _02_ _47_/a_81_21# 1.59e-20
C2855 net1 p[1] 0.0291f
C2856 p[10] net19 1.26e-21
C2857 _37_/a_27_47# _42_/a_109_93# 2.55e-20
C2858 th07_0/m1_808_n892# VGND 0.0127f
C2859 th15_0/Vin p[11] 0.186f
C2860 p[10] input1/a_75_212# 0.00136f
C2861 _47_/a_81_21# p[14] 1.42e-21
C2862 _03_ _30_/a_297_297# 0.00117f
C2863 net10 net12 0.539f
C2864 _02_ _22_ 0.552f
C2865 _26_/a_183_297# _06_ 3.16e-19
C2866 _10_ net12 0.00257f
C2867 input2/a_27_47# net8 0.0207f
C2868 VPWR p[12] 0.144f
C2869 _48_/a_109_47# _07_ 3.01e-19
C2870 _18_ net12 2.25e-21
C2871 p[5] th07_0/m1_808_n892# 0.00441f
C2872 _21_ _11_ 9.98e-20
C2873 _03_ _32_/a_27_47# 1.9e-19
C2874 VPWR b[2] 0.262f
C2875 _15_ _50_/a_27_47# 5.65e-19
C2876 _00_ net3 2.12e-19
C2877 _00_ net8 3.23e-19
C2878 _04_ net10 0.121f
C2879 Vin input12/a_27_47# 0.00444f
C2880 _04_ _10_ 9.24e-20
C2881 _25_ _06_ 0.144f
C2882 _04_ _18_ 1.94e-21
C2883 VPWR _55_/a_217_297# -0.00133f
C2884 _13_ _50_/a_27_47# 0.00169f
C2885 _36_/a_27_47# _29_/a_29_53# 6.92e-20
C2886 p[10] b[1] 0.114f
C2887 Vin b[3] 0.0166f
C2888 _10_ th15_0/m1_849_n157# 1.54e-19
C2889 _12_ _47_/a_299_297# 0.00805f
C2890 _36_/a_27_47# _06_ 0.0501f
C2891 net16 _38_/a_197_47# 5.89e-19
C2892 Vin th12_0/m1_529_n42# 0.0341f
C2893 _49_/a_544_297# b[1] 8.23e-19
C2894 _10_ _38_/a_197_47# 6.29e-19
C2895 net7 output17/a_27_47# 0.0018f
C2896 net1 net7 0.0712f
C2897 _44_/a_93_21# p[11] 7.91e-19
C2898 _09_ net18 1.97e-21
C2899 _03_ _49_/a_315_47# 9.22e-19
C2900 p[2] _49_/a_75_199# 2.21e-19
C2901 VPWR input4/a_75_212# 0.0608f
C2902 net17 _30_/a_109_53# 4.18e-20
C2903 net17 th02_0/m1_983_133# 1.59e-19
C2904 VPWR th04_0/m1_620_n488# 0.00264f
C2905 net13 _22_ 4.63e-20
C2906 Vin VGND 1.48f
C2907 p[9] input6/a_27_47# 0.0756f
C2908 _43_/a_193_413# _14_ 0.0297f
C2909 net7 input5/a_841_47# 0.00193f
C2910 p[13] input1/a_75_212# 4.16e-19
C2911 _36_/a_197_47# net6 6.94e-20
C2912 _20_ net2 8.83e-19
C2913 _15_ input6/a_27_47# 4.43e-19
C2914 net15 _06_ 0.033f
C2915 VGND _37_/a_303_47# -1.63e-19
C2916 _53_/a_111_297# _06_ 3.82e-19
C2917 p[5] Vin 0.335f
C2918 _26_/a_29_53# _20_ 0.00447f
C2919 _55_/a_80_21# _55_/a_472_297# 1.78e-33
C2920 _19_ net17 0.0211f
C2921 p[6] input12/a_27_47# 0.0225f
C2922 p[12] input4/a_75_212# 0.0278f
C2923 _29_/a_29_53# _06_ 0.00111f
C2924 _31_/a_35_297# _05_ 0.00649f
C2925 th15_0/Vin _42_/a_209_311# 2.47e-20
C2926 _03_ _15_ 7.39e-20
C2927 _19_ _49_/a_75_199# 0.0206f
C2928 _12_ b[1] 3.18e-21
C2929 _33_/a_209_311# net12 0.0769f
C2930 _32_/a_303_47# net1 1.45e-19
C2931 _35_/a_76_199# _05_ 0.00238f
C2932 _52_/a_93_21# _39_/a_47_47# 1.44e-20
C2933 _17_ th15_0/Vin 0.00232f
C2934 input3/a_27_47# _15_ 7.53e-19
C2935 p[13] b[1] 0.00201f
C2936 _26_/a_111_297# VGND -2.75e-19
C2937 _14_ p[9] 2.62e-21
C2938 _44_/a_256_47# net14 0.00379f
C2939 _44_/a_346_47# net3 8.04e-19
C2940 _13_ _03_ 1.74e-20
C2941 _23_ net9 1.21e-19
C2942 _15_ _14_ 0.148f
C2943 net1 input9/a_75_212# 0.002f
C2944 _35_/a_489_413# _08_ 5.56e-19
C2945 _35_/a_76_199# _09_ 0.047f
C2946 _00_ _20_ 0.271f
C2947 net2 _50_/a_343_93# 1.25e-20
C2948 net1 _55_/a_80_21# 1.8e-19
C2949 _04_ _33_/a_209_311# 0.00133f
C2950 _39_/a_47_47# b[0] 2.04e-19
C2951 net14 input7/a_27_47# 3.48e-19
C2952 _13_ _14_ 1.47e-20
C2953 p[6] VGND 0.251f
C2954 _37_/a_27_47# net6 4.3e-20
C2955 input10/a_27_47# input11/a_27_47# 5.3e-19
C2956 _26_/a_29_53# _50_/a_343_93# 2.61e-19
C2957 _02_ _38_/a_27_47# 0.00103f
C2958 _19_ input5/a_62_47# 0.00159f
C2959 p[2] net9 1.4e-20
C2960 _10_ _55_/a_472_297# 7.35e-21
C2961 _27_/a_277_297# p[1] 1.66e-20
C2962 _09_ net5 5.18e-19
C2963 net4 _38_/a_303_47# 5.95e-19
C2964 net3 _40_/a_297_297# 2.54e-19
C2965 p[5] p[6] 0.348f
C2966 p[10] _27_/a_27_297# 1.63e-19
C2967 b[1] _34_/a_47_47# 0.0197f
C2968 p[7] net9 8.26e-19
C2969 _44_/a_93_21# _42_/a_209_311# 2.21e-19
C2970 _44_/a_250_297# _42_/a_109_93# 6.38e-19
C2971 input8/a_27_47# input7/a_27_47# 3.2e-20
C2972 _30_/a_109_53# net9 0.0191f
C2973 _39_/a_285_47# _06_ 1.23e-20
C2974 _02_ _52_/a_93_21# 0.0962f
C2975 b[1] _55_/a_300_47# 1.1e-19
C2976 _11_ net6 0.0257f
C2977 _36_/a_197_47# _10_ 1.54e-19
C2978 _04_ _27_/a_109_297# 7.2e-20
C2979 _44_/a_93_21# _17_ 0.0646f
C2980 _34_/a_47_47# _48_/a_27_47# 4.45e-21
C2981 VPWR th15_0/m1_597_n912# 2.46e-19
C2982 _45_/a_27_47# _35_/a_226_47# 5.71e-21
C2983 net10 output17/a_27_47# 1.31e-20
C2984 net4 _12_ 0.105f
C2985 _36_/a_27_47# _50_/a_27_47# 6.08e-19
C2986 _45_/a_27_47# _07_ 1.02e-20
C2987 _45_/a_193_297# _06_ 0.00201f
C2988 _00_ _50_/a_343_93# 0.102f
C2989 net10 net1 0.00388f
C2990 net1 _10_ 4.34e-19
C2991 _12_ _33_/a_109_93# 9.75e-20
C2992 _35_/a_226_47# _23_ 4.21e-19
C2993 _39_/a_129_47# net5 0.00344f
C2994 p[13] p[8] 0.00239f
C2995 _23_ _07_ 1.27e-19
C2996 _31_/a_285_47# p[10] 2.16e-20
C2997 VPWR _33_/a_296_53# -1.15e-19
C2998 net8 p[2] 0.0146f
C2999 net14 _02_ 0.00952f
C3000 _01_ _49_/a_544_297# 0.00109f
C3001 _45_/a_109_297# net5 0.0184f
C3002 _31_/a_285_297# _02_ 5.86e-20
C3003 _37_/a_109_47# net19 1.16e-20
C3004 p[12] th15_0/m1_597_n912# 0.0395f
C3005 _47_/a_81_21# net2 4.95e-19
C3006 net8 _30_/a_109_53# 1.76e-20
C3007 net14 p[14] 0.00278f
C3008 _35_/a_489_413# _02_ 3.86e-19
C3009 _44_/a_584_47# b[3] 1.27e-19
C3010 _12_ _52_/a_250_297# 0.0139f
C3011 _47_/a_384_47# _11_ 7.23e-20
C3012 _15_ input5/a_664_47# 9.15e-22
C3013 p[7] _35_/a_226_47# 2.84e-19
C3014 _44_/a_584_47# th12_0/m1_529_n42# 1.38e-20
C3015 _05_ VGND 0.754f
C3016 VPWR _52_/a_346_47# -0.00109f
C3017 p[7] _07_ 0.00283f
C3018 th15_0/Vin th01_0/m1_991_n1219# -8.41e-19
C3019 VPWR th15_0/Vin 0.945f
C3020 net2 _22_ 1.93e-20
C3021 _02_ input8/a_27_47# 5.08e-20
C3022 p[10] _42_/a_109_93# 1.82e-21
C3023 VPWR _27_/a_205_297# 1.05e-19
C3024 _31_/a_35_297# _32_/a_27_47# 9.17e-20
C3025 _52_/a_93_21# net13 7.21e-19
C3026 _29_/a_29_53# _50_/a_27_47# 1.44e-20
C3027 th08_0/m1_477_n803# p[2] 3.32e-21
C3028 p[13] _27_/a_27_297# 2.6e-19
C3029 _06_ _50_/a_27_47# 0.00972f
C3030 _18_ _37_/a_27_47# 3.31e-20
C3031 _09_ VGND 0.397f
C3032 _19_ net8 0.0322f
C3033 _19_ net3 0.0129f
C3034 _26_/a_29_53# _22_ 0.09f
C3035 _26_/a_183_297# _14_ 6.98e-22
C3036 Vin net17 0.00133f
C3037 _04_ _42_/a_209_311# 9.84e-22
C3038 p[7] p[4] 7.8e-20
C3039 p[7] th08_0/m1_477_n803# 0.0155f
C3040 _44_/a_584_47# VGND -0.00145f
C3041 _03_ _25_ 0.00422f
C3042 p[3] th04_0/m1_892_n998# 0.0241f
C3043 net16 _11_ 0.172f
C3044 _20_ _40_/a_297_297# 9.18e-21
C3045 _17_ _04_ 4.34e-19
C3046 th15_0/Vin p[12] 0.175f
C3047 _10_ _11_ 0.176f
C3048 _00_ _47_/a_81_21# 0.0258f
C3049 th15_0/m1_597_n912# input4/a_75_212# 8.81e-20
C3050 p[13] _01_ 4.28e-19
C3051 _18_ _11_ 0.484f
C3052 net14 net13 2.21e-21
C3053 _17_ th15_0/m1_849_n157# 8.52e-20
C3054 _31_/a_285_297# net13 3.85e-20
C3055 _32_/a_27_47# net5 0.0961f
C3056 _12_ _35_/a_226_297# 3.35e-20
C3057 th04_0/m1_892_n998# net13 2.29e-19
C3058 p[10] p[1] 9.56e-19
C3059 net15 input6/a_27_47# 0.00115f
C3060 _02_ _16_ 0.00564f
C3061 _24_ _07_ 5.67e-19
C3062 _09_ _53_/a_183_297# 4.18e-19
C3063 p[3] input8/a_27_47# 0.0023f
C3064 input14/a_27_47# p[9] 8.53e-21
C3065 _39_/a_129_47# VGND -0.00126f
C3066 th14_0/m1_641_n318# th12_0/m1_394_n856# 1.54e-19
C3067 _00_ _22_ 0.477f
C3068 _35_/a_489_413# net13 7.36e-20
C3069 p[14] _16_ 1.74e-21
C3070 VPWR _44_/a_93_21# 0.005f
C3071 net10 _30_/a_392_297# 3.4e-19
C3072 _43_/a_297_47# _06_ 4.81e-20
C3073 _12_ _21_ 7.99e-20
C3074 _06_ input6/a_27_47# 2.85e-19
C3075 _45_/a_109_297# VGND -0.00179f
C3076 _30_/a_215_297# net12 0.00676f
C3077 net10 _33_/a_368_53# 0.00171f
C3078 _20_ p[2] 3.01e-20
C3079 _03_ net15 4.26e-20
C3080 input11/a_27_47# VGND 0.0274f
C3081 VPWR _42_/a_296_53# -6.37e-20
C3082 th11_0/m1_705_187# Vin 0.0585f
C3083 _43_/a_193_413# net5 1.39e-20
C3084 th15_0/Vin input4/a_75_212# 0.00104f
C3085 input3/a_27_47# net15 6.19e-20
C3086 b[1] _54_/a_75_212# 0.0023f
C3087 _03_ _29_/a_29_53# 0.0414f
C3088 _20_ _30_/a_109_53# 8.12e-19
C3089 net16 th13_0/m1_831_275# 1.81e-20
C3090 net15 _14_ 0.0538f
C3091 _01_ _55_/a_300_47# 0.00113f
C3092 p[5] input11/a_27_47# 0.0506f
C3093 _03_ _06_ 0.00635f
C3094 _04_ _30_/a_215_297# 0.00225f
C3095 _10_ th13_0/m1_831_275# 7.72e-20
C3096 net11 _12_ 0.00799f
C3097 _14_ _06_ 0.0556f
C3098 _40_/a_109_297# net6 2.53e-20
C3099 p[10] net7 0.00695f
C3100 _21_ _34_/a_47_47# 8.93e-19
C3101 VGND _30_/a_297_297# -5.13e-19
C3102 _19_ _20_ 0.00734f
C3103 Vin net9 5.21e-19
C3104 VPWR net12 0.82f
C3105 b[1] _30_/a_465_297# 4.8e-19
C3106 _13_ _35_/a_76_199# 3.01e-21
C3107 _49_/a_544_297# net7 2.72e-19
C3108 th08_0/m1_477_n803# th07_0/m1_808_n892# 6.27e-19
C3109 th07_0/m1_808_n892# p[4] 1.11e-20
C3110 VPWR _32_/a_197_47# 0.00146f
C3111 _15_ net5 0.0352f
C3112 output19/a_27_47# net14 0.00142f
C3113 _32_/a_27_47# VGND 0.0233f
C3114 th03_0/m1_890_n844# p[2] 0.0404f
C3115 _28_/a_109_297# _11_ 6.29e-19
C3116 VPWR _04_ 0.456f
C3117 _13_ net5 0.0381f
C3118 _43_/a_27_47# _20_ 0.0124f
C3119 net14 input5/a_381_47# 0.00479f
C3120 net15 _49_/a_201_297# 1.41e-19
C3121 p[7] th03_0/m1_890_n844# 1.48e-20
C3122 net11 _34_/a_47_47# 0.0309f
C3123 VPWR th15_0/m1_849_n157# 0.0316f
C3124 th03_0/m1_890_n844# th02_0/m1_983_133# 0.0135f
C3125 _24_ _53_/a_29_53# 0.0835f
C3126 Vin net8 0.00767f
C3127 Vin net3 0.00372f
C3128 net14 th14_0/m1_891_419# 4.02e-21
C3129 _31_/a_117_297# Vin 3.9e-19
C3130 VPWR _38_/a_197_47# -5.24e-19
C3131 input1/a_75_212# input7/a_27_47# 3.2e-20
C3132 _05_ net17 0.0111f
C3133 _43_/a_193_413# VGND -0.0147f
C3134 _45_/a_193_297# _03_ 2.57e-20
C3135 _49_/a_315_47# VGND -0.0034f
C3136 net3 _37_/a_303_47# 0.00133f
C3137 net14 _37_/a_197_47# 7e-19
C3138 Vin _07_ 2.86e-19
C3139 _08_ b[1] 0.0127f
C3140 _25_ net18 0.0594f
C3141 p[12] th15_0/m1_849_n157# 0.0103f
C3142 p[9] b[3] 0.134f
C3143 th14_0/m1_641_n318# net15 4.16e-20
C3144 net11 _36_/a_303_47# 7.63e-20
C3145 net15 input5/a_664_47# 0.0216f
C3146 _45_/a_27_47# _22_ 0.0131f
C3147 p[13] net7 4.55e-19
C3148 p[3] input13/a_27_47# 0.00107f
C3149 _23_ _22_ 0.0187f
C3150 net14 net2 0.151f
C3151 _09_ _49_/a_75_199# 2.93e-19
C3152 th15_0/Vin th15_0/m1_597_n912# 0.00183f
C3153 _08_ _48_/a_27_47# 2.58e-19
C3154 Vin p[4] 0.0788f
C3155 th08_0/m1_477_n803# Vin 0.0494f
C3156 _13_ _45_/a_205_47# 7.51e-20
C3157 input10/a_27_47# _25_ 2.03e-20
C3158 input5/a_664_47# _06_ 3.21e-19
C3159 _34_/a_285_47# VGND -0.00301f
C3160 b[1] input7/a_27_47# 0.00663f
C3161 _26_/a_29_53# net14 1.33e-20
C3162 p[9] _41_/a_59_75# 1.02e-19
C3163 _12_ net6 0.0891f
C3164 input13/a_27_47# net13 0.00139f
C3165 _15_ _41_/a_59_75# 0.0143f
C3166 _38_/a_27_47# output16/a_27_47# 9.02e-19
C3167 th09_0/m1_485_n505# p[14] 1.95e-20
C3168 VGND p[9] 0.443f
C3169 _37_/a_27_47# _42_/a_209_311# 1.59e-20
C3170 VGND _15_ 0.15f
C3171 th06_0/m1_904_n796# th05_0/m1_752_n794# 9.46e-19
C3172 _02_ net19 0.0474f
C3173 net14 input2/a_27_47# 0.0102f
C3174 _17_ _37_/a_27_47# 0.00277f
C3175 input15/a_27_47# _16_ 7.13e-19
C3176 _13_ VGND 0.363f
C3177 _30_/a_109_53# _22_ 3.67e-21
C3178 p[14] net19 0.06f
C3179 _49_/a_208_47# b[1] 2.93e-19
C3180 _15_ _50_/a_223_47# 0.00698f
C3181 p[6] _07_ 4.16e-19
C3182 net1 _30_/a_215_297# 0.00375f
C3183 _00_ net14 4.11e-20
C3184 _43_/a_193_413# _43_/a_369_47# -1.25e-19
C3185 net18 _06_ 0.0211f
C3186 th12_0/m1_394_n856# th12_0/m1_529_n42# 1.78e-33
C3187 VPWR _55_/a_472_297# 0.00488f
C3188 _13_ _50_/a_223_47# 8.2e-20
C3189 output16/a_27_47# b[0] 0.014f
C3190 _17_ _11_ 0.197f
C3191 _35_/a_76_199# _36_/a_27_47# 3.22e-19
C3192 _12_ _47_/a_384_47# 9.51e-20
C3193 _05_ net9 0.124f
C3194 Vin _20_ 6.26e-20
C3195 net16 _38_/a_303_47# 6.47e-19
C3196 net2 _16_ 0.00654f
C3197 p[6] p[4] 0.00576f
C3198 th08_0/m1_477_n803# p[6] 4.52e-19
C3199 _25_ net5 6.42e-19
C3200 _02_ b[1] 0.00718f
C3201 _10_ _38_/a_303_47# 7.36e-19
C3202 th12_0/m1_394_n856# VGND 0.0134f
C3203 _44_/a_250_297# p[11] 0.00177f
C3204 _24_ _22_ 0.0846f
C3205 _09_ net9 2.62e-19
C3206 VPWR _36_/a_197_47# -5.24e-19
C3207 _36_/a_27_47# net5 0.0163f
C3208 net4 _39_/a_47_47# 0.0202f
C3209 VPWR output17/a_27_47# 0.0268f
C3210 _02_ _48_/a_27_47# 0.00435f
C3211 VPWR net1 1.17f
C3212 input10/a_27_47# th05_0/m1_752_n794# 1.29e-19
C3213 net16 _12_ 0.131f
C3214 _43_/a_27_47# _22_ 0.091f
C3215 _43_/a_297_47# _14_ 9.11e-19
C3216 _14_ input6/a_27_47# 3.75e-21
C3217 _36_/a_303_47# net6 1.25e-19
C3218 _12_ net10 7.82e-20
C3219 _12_ _10_ 0.19f
C3220 _44_/a_93_21# th15_0/Vin 0.00197f
C3221 net11 _54_/a_75_212# 0.00956f
C3222 _12_ _18_ 0.0115f
C3223 VPWR input5/a_841_47# 0.0775f
C3224 _35_/a_76_199# _29_/a_29_53# 9.88e-19
C3225 th09_0/m1_485_n505# th10_0/m1_536_174# 0.00429f
C3226 _05_ net8 0.0146f
C3227 _35_/a_76_199# _06_ 0.00425f
C3228 _00_ _16_ 0.00613f
C3229 p[3] b[1] 0.00473f
C3230 th15_0/Vin _42_/a_296_53# 7.75e-21
C3231 net15 net5 0.0226f
C3232 _27_/a_27_297# input7/a_27_47# 0.00119f
C3233 _33_/a_296_53# net12 1.23e-20
C3234 Vin th03_0/m1_890_n844# 0.0269f
C3235 _35_/a_226_47# _05_ 0.0134f
C3236 _05_ _07_ 1.21e-19
C3237 _26_/a_183_297# VGND 2.42e-19
C3238 b[1] net13 0.0495f
C3239 net5 _29_/a_29_53# 8.1e-20
C3240 _44_/a_346_47# net14 0.00464f
C3241 VPWR _37_/a_27_47# -0.0178f
C3242 th01_0/m1_571_n501# p[0] 2.36e-19
C3243 net5 _06_ 0.41f
C3244 _35_/a_226_47# _09_ 0.0599f
C3245 net4 _02_ 0.00376f
C3246 p[10] p[11] 0.00389f
C3247 _09_ _07_ 0.0416f
C3248 _45_/a_27_47# _52_/a_93_21# 1.18e-19
C3249 th15_0/m1_597_n912# th15_0/m1_849_n157# -5.55e-35
C3250 VPWR th10_0/m1_502_n495# 0.0291f
C3251 net10 _34_/a_47_47# 0.0507f
C3252 _02_ _33_/a_109_93# 1.54e-21
C3253 p[8] p[14] 1.91e-20
C3254 _52_/a_93_21# _23_ 0.0166f
C3255 VGND _25_ 0.199f
C3256 _08_ _21_ 0.00139f
C3257 VPWR _11_ 0.352f
C3258 _36_/a_27_47# VGND 0.0211f
C3259 b[1] _34_/a_377_297# 0.00115f
C3260 _48_/a_181_47# _02_ 3.9e-19
C3261 net15 b[3] 0.00264f
C3262 _03_ _49_/a_201_297# 0.00842f
C3263 _30_/a_297_297# net9 7.53e-19
C3264 output19/a_27_47# net19 0.0273f
C3265 _02_ _52_/a_250_297# 0.0128f
C3266 net15 th12_0/m1_529_n42# 2.01e-21
C3267 _01_ _49_/a_208_47# 2.13e-19
C3268 input12/a_27_47# _06_ 5.3e-22
C3269 _36_/a_303_47# _10_ 4.09e-19
C3270 _27_/a_27_297# _02_ 0.00179f
C3271 _04_ _27_/a_205_297# 6.42e-19
C3272 _44_/a_250_297# _17_ 0.0336f
C3273 p[3] _33_/a_109_93# 1.64e-19
C3274 th15_0/Vin th15_0/m1_849_n157# 0.173f
C3275 _45_/a_27_47# _35_/a_489_413# 3.89e-21
C3276 _45_/a_109_297# _35_/a_226_47# 1.59e-21
C3277 net19 input5/a_381_47# 0.00173f
C3278 _36_/a_27_47# _50_/a_223_47# 1.27e-20
C3279 _49_/a_201_297# _14_ 4.76e-21
C3280 b[3] _06_ 9.96e-21
C3281 net11 _08_ 8.83e-19
C3282 _32_/a_27_47# net9 0.0136f
C3283 p[12] _11_ 3.66e-20
C3284 _12_ _33_/a_209_311# 2.88e-20
C3285 _39_/a_285_47# net5 0.05f
C3286 net15 _41_/a_59_75# 1.16e-20
C3287 _15_ input5/a_558_47# 0.00166f
C3288 net4 net13 2.48e-19
C3289 input12/a_27_47# th05_0/m1_752_n794# 4.98e-20
C3290 VPWR _33_/a_368_53# -4.26e-19
C3291 net15 VGND 0.222f
C3292 _31_/a_285_297# p[2] 0.00165f
C3293 input15/a_27_47# net19 0.00231f
C3294 _33_/a_109_93# net13 0.0254f
C3295 th04_0/m1_892_n998# p[2] 0.0503f
C3296 _05_ _20_ 6.79e-19
C3297 _53_/a_111_297# VGND -2.89e-19
C3298 _01_ _02_ 0.106f
C3299 _45_/a_193_297# net5 0.00935f
C3300 p[13] p[11] 0.0167f
C3301 _06_ _41_/a_59_75# 0.0457f
C3302 _17_ _40_/a_109_297# 9.67e-19
C3303 _45_/a_465_47# _09_ 2.77e-19
C3304 VGND _29_/a_29_53# 0.0544f
C3305 p[7] th04_0/m1_892_n998# 0.00187f
C3306 _47_/a_299_297# net2 1.18e-19
C3307 input11/a_27_47# p[4] 0.0648f
C3308 net8 _30_/a_297_297# 2.42e-21
C3309 VGND _06_ 1.1f
C3310 _09_ _20_ 7.11e-19
C3311 th14_0/m1_641_n318# input3/a_27_47# 4.43e-19
C3312 VPWR th13_0/m1_831_275# 0.0295f
C3313 th04_0/m1_892_n998# _30_/a_109_53# 2.97e-20
C3314 th04_0/m1_892_n998# th02_0/m1_983_133# 8.54e-21
C3315 VPWR _36_/a_109_47# -4.66e-19
C3316 input7/a_27_47# p[1] 0.0164f
C3317 _24_ _52_/a_93_21# 0.0211f
C3318 p[2] input8/a_27_47# 0.0217f
C3319 p[7] _35_/a_489_413# 3.02e-20
C3320 VPWR _52_/a_584_47# -9.47e-19
C3321 _32_/a_109_47# _01_ 0.00129f
C3322 b[1] input5/a_381_47# 0.0023f
C3323 net2 net19 0.599f
C3324 _44_/a_93_21# _04_ 4.47e-21
C3325 p[10] _42_/a_209_311# 2.37e-20
C3326 VPWR _27_/a_277_297# -3.63e-19
C3327 _32_/a_27_47# net8 0.0275f
C3328 _29_/a_29_53# _50_/a_223_47# 1.45e-20
C3329 VGND th05_0/m1_752_n794# 0.0192f
C3330 p[8] th10_0/m1_536_174# 0.0134f
C3331 _06_ _50_/a_223_47# 0.0481f
C3332 _02_ _21_ 0.397f
C3333 _34_/a_47_47# _33_/a_209_311# 0.017f
C3334 output18/a_27_47# _54_/a_75_212# 2.28e-19
C3335 _09_ _53_/a_29_53# 0.00642f
C3336 _19_ net14 0.0512f
C3337 _26_/a_111_297# _22_ 0.00137f
C3338 _19_ _31_/a_285_297# 1.34e-19
C3339 _53_/a_183_297# _06_ 0.00146f
C3340 p[12] th13_0/m1_831_275# 0.00668f
C3341 _20_ _39_/a_129_47# 1.71e-20
C3342 _03_ net18 2.07e-21
C3343 p[5] th05_0/m1_752_n794# 0.00925f
C3344 net5 _50_/a_27_47# 0.0169f
C3345 _08_ net7 9.54e-25
C3346 input2/a_27_47# net19 2.9e-23
C3347 _00_ _47_/a_299_297# 7.59e-21
C3348 _05_ th03_0/m1_890_n844# 9.65e-20
C3349 _01_ net13 0.00228f
C3350 net9 _15_ 0.00113f
C3351 _43_/a_193_413# net8 1.62e-20
C3352 _43_/a_193_413# net3 5.65e-20
C3353 _43_/a_27_47# net14 4.87e-20
C3354 net11 _02_ 0.0327f
C3355 input3/a_27_47# input14/a_27_47# 5.08e-20
C3356 _39_/a_285_47# VGND -0.0046f
C3357 b[1] net2 0.0389f
C3358 net16 _54_/a_75_212# 1.69e-21
C3359 p[8] output19/a_27_47# 0.0094f
C3360 _35_/a_226_297# net13 6.88e-19
C3361 p[3] _21_ 2.13e-20
C3362 net7 input7/a_27_47# 0.00318f
C3363 VPWR _44_/a_250_297# 0.0233f
C3364 _04_ net12 0.267f
C3365 net10 _54_/a_75_212# 7.43e-19
C3366 _43_/a_369_47# _06_ -2.02e-19
C3367 _26_/a_29_53# b[1] 9.93e-21
C3368 _45_/a_193_297# VGND -0.00241f
C3369 _48_/a_109_47# b[1] 9.32e-20
C3370 _31_/a_35_297# _03_ 0.00749f
C3371 _21_ net13 0.13f
C3372 VPWR _42_/a_368_53# -3.03e-19
C3373 b[1] input2/a_27_47# 0.014f
C3374 _17_ _12_ 0.0109f
C3375 net3 p[9] 1.63e-19
C3376 _35_/a_76_199# _03_ 0.0733f
C3377 net8 _15_ 1.79e-19
C3378 net3 _15_ 0.224f
C3379 th04_0/m1_892_n998# th07_0/m1_808_n892# 2.34e-19
C3380 VPWR _40_/a_109_297# -4.23e-19
C3381 net10 _30_/a_465_297# 0.00106f
C3382 th15_0/Vin output17/a_27_47# 1.87e-20
C3383 net11 p[3] 5.73e-20
C3384 _49_/a_208_47# net7 0.00312f
C3385 net1 th15_0/Vin 4.02e-19
C3386 p[0] VGND 0.423f
C3387 _34_/a_285_47# _07_ 0.00975f
C3388 Vin _38_/a_27_47# 5.31e-19
C3389 _39_/a_47_47# net6 0.0249f
C3390 _32_/a_27_47# _20_ 0.0069f
C3391 _40_/a_191_297# net6 1.16e-20
C3392 net11 net13 0.093f
C3393 _21_ _34_/a_377_297# 2.37e-19
C3394 th15_0/Vin input5/a_841_47# 9.9e-20
C3395 _03_ net5 1.04e-19
C3396 _50_/a_27_47# _41_/a_59_75# 9.59e-22
C3397 _43_/a_27_47# _16_ 2.47e-19
C3398 _27_/a_27_297# input5/a_381_47# 1.47e-19
C3399 p[8] net2 0.0279f
C3400 _13_ _35_/a_226_47# 5.62e-21
C3401 VGND _50_/a_27_47# -0.00432f
C3402 _05_ _22_ 3.33e-21
C3403 _13_ _07_ 3.22e-23
C3404 _02_ net7 0.445f
C3405 p[10] th01_0/m1_991_n1219# 0.00424f
C3406 VPWR p[10] 0.433f
C3407 _14_ net5 3.89e-19
C3408 _26_/a_29_53# net4 0.00412f
C3409 _09_ _22_ 0.0279f
C3410 net15 net17 5.19e-19
C3411 VPWR _49_/a_544_297# 0.00504f
C3412 th15_0/Vin _37_/a_27_47# 0.00332f
C3413 _44_/a_346_47# net19 0.00124f
C3414 _43_/a_193_413# _20_ 0.00161f
C3415 b[3] input6/a_27_47# 4.02e-19
C3416 _31_/a_35_297# _49_/a_201_297# 5.52e-20
C3417 Vin b[0] 1.65e-19
C3418 th10_0/m1_502_n495# th15_0/Vin 0.0036f
C3419 net15 _49_/a_75_199# 5.13e-20
C3420 p[7] input13/a_27_47# 0.0171f
C3421 net15 input5/a_558_47# 0.00672f
C3422 _08_ net10 0.194f
C3423 _32_/a_27_47# _50_/a_343_93# 6.48e-20
C3424 _08_ _10_ 1.51e-19
C3425 _02_ net6 0.00427f
C3426 _12_ _38_/a_109_47# 0.00179f
C3427 Vin net14 0.00129f
C3428 _31_/a_285_297# Vin 3.61e-19
C3429 VPWR _38_/a_303_47# -4.83e-19
C3430 Vin th04_0/m1_892_n998# 0.0366f
C3431 _49_/a_75_199# _29_/a_29_53# 1.28e-19
C3432 _27_/a_27_297# net2 0.0131f
C3433 th15_0/Vin _11_ 0.00308f
C3434 p[14] net6 0.00518f
C3435 net4 _00_ 0.0166f
C3436 _43_/a_297_47# VGND -1.33e-19
C3437 input5/a_558_47# _06_ 3.55e-19
C3438 net14 _37_/a_303_47# 0.00112f
C3439 output19/a_27_47# _42_/a_109_93# 1.56e-20
C3440 VGND input6/a_27_47# -0.00236f
C3441 _32_/a_303_47# _02_ 1.15e-20
C3442 input3/a_27_47# b[3] 1.4e-19
C3443 th13_0/m1_831_275# th15_0/m1_597_n912# 0.0186f
C3444 net16 _39_/a_47_47# 7.7e-20
C3445 input5/a_381_47# _42_/a_109_93# 0.00763f
C3446 _45_/a_109_297# _22_ 0.0426f
C3447 Vin input8/a_27_47# 0.00586f
C3448 net13 net7 1.72e-19
C3449 _20_ _15_ 0.691f
C3450 net10 _39_/a_47_47# 4.72e-22
C3451 VPWR _12_ 0.28f
C3452 _10_ _39_/a_47_47# 0.00824f
C3453 net4 output16/a_27_47# 0.00706f
C3454 _36_/a_27_47# net9 0.00493f
C3455 _01_ net2 2.72e-19
C3456 _02_ _55_/a_80_21# 0.164f
C3457 _02_ output18/a_27_47# 4.13e-19
C3458 _36_/a_197_47# net12 4.67e-20
C3459 _27_/a_27_297# input2/a_27_47# 1.16e-19
C3460 _18_ _39_/a_47_47# 1.23e-19
C3461 _44_/a_93_21# _37_/a_27_47# 3.19e-19
C3462 _13_ _45_/a_465_47# 0.00134f
C3463 _03_ VGND 0.119f
C3464 p[13] VPWR 0.318f
C3465 input10/a_27_47# net18 4.16e-20
C3466 th14_0/m1_891_419# _42_/a_109_93# 1.58e-19
C3467 _13_ _20_ 7.38e-21
C3468 _29_/a_183_297# _09_ 4.51e-20
C3469 net1 net12 1.17e-19
C3470 input3/a_27_47# VGND 0.0414f
C3471 VGND _14_ 0.226f
C3472 _32_/a_197_47# net1 0.00142f
C3473 net13 net6 0.00188f
C3474 _12_ p[12] 0.00589f
C3475 _03_ _50_/a_223_47# 1.41e-21
C3476 input5/a_664_47# net5 0.0536f
C3477 _44_/a_93_21# _11_ 4.78e-20
C3478 _17_ _37_/a_109_47# 8.86e-21
C3479 th04_0/m1_892_n998# p[6] 9.47e-20
C3480 th15_0/Vin th13_0/m1_831_275# 0.00711f
C3481 _13_ _53_/a_29_53# 9.05e-19
C3482 net15 net9 8.49e-20
C3483 Vin _16_ 6.65e-20
C3484 _04_ net1 0.018f
C3485 _04_ output17/a_27_47# 0.027f
C3486 _12_ b[2] 3.89e-20
C3487 _32_/a_27_47# _47_/a_81_21# 5.06e-21
C3488 net2 _42_/a_109_93# 0.00507f
C3489 p[3] input9/a_75_212# 0.0171f
C3490 net16 _02_ 8.94e-19
C3491 b[1] _23_ 7.65e-19
C3492 _15_ _50_/a_343_93# 0.0098f
C3493 net8 _36_/a_27_47# 1.52e-19
C3494 VPWR _34_/a_47_47# 0.0372f
C3495 input1/a_75_212# th02_0/m1_983_133# 5.8e-20
C3496 _00_ _01_ 0.00124f
C3497 net10 _02_ 6.74e-19
C3498 net9 _29_/a_29_53# 0.0205f
C3499 _02_ _10_ 0.0537f
C3500 net9 _06_ 0.0505f
C3501 _18_ _02_ 2.96e-20
C3502 VPWR _55_/a_300_47# -4.61e-19
C3503 _32_/a_27_47# _22_ 1.76e-19
C3504 th04_0/m1_892_n998# 0 0.832f
C3505 p[3] 0 0.52f
C3506 th04_0/m1_620_n488# 0 0.0632f
C3507 Vin 0 15.9f
C3508 th11_0/m1_705_187# 0 0.602f
C3509 p[10] 0 0.502f
C3510 th11_0/m1_577_n654# 0 0.286f
C3511 th06_0/m1_904_n796# 0 0.495f
C3512 p[5] 0 0.861f
C3513 th13_0/m1_831_275# 0 1.05f
C3514 p[12] 0 0.639f
C3515 th13_0/m1_559_n458# 0 0.286f
C3516 th08_0/m1_477_n803# 0 0.577f
C3517 p[7] 0 0.583f
C3518 _03_ 0 0.36f
C3519 net10 0 0.418f
C3520 _30_/a_109_53# 0 0.159f
C3521 _30_/a_215_297# 0 0.142f
C3522 p[14] 0 0.608f
C3523 th15_0/m1_849_n157# 0 1.28f
C3524 th15_0/m1_597_n912# 0 0.19f
C3525 _05_ 0 0.152f
C3526 _31_/a_285_297# 0 0.00137f
C3527 _31_/a_35_297# 0 0.255f
C3528 _32_/a_27_47# 0 0.175f
C3529 _50_/a_343_93# 0 0.172f
C3530 _50_/a_223_47# 0 0.141f
C3531 _50_/a_27_47# 0 0.259f
C3532 _07_ 0 0.285f
C3533 _06_ 0 0.779f
C3534 _33_/a_209_311# 0 0.143f
C3535 _33_/a_109_93# 0 0.158f
C3536 _34_/a_285_47# 0 0.0174f
C3537 _34_/a_47_47# 0 0.199f
C3538 _23_ 0 0.106f
C3539 _09_ 0 0.142f
C3540 _08_ 0 0.128f
C3541 _35_/a_489_413# 0 0.0254f
C3542 _35_/a_226_47# 0 0.162f
C3543 _35_/a_76_199# 0 0.141f
C3544 input15/a_27_47# 0 0.208f
C3545 _24_ 0 0.135f
C3546 _12_ 0 0.378f
C3547 _52_/a_250_297# 0 0.0278f
C3548 _52_/a_93_21# 0 0.151f
C3549 _10_ 0 0.624f
C3550 _36_/a_27_47# 0 0.175f
C3551 _53_/a_29_53# 0 0.18f
C3552 input14/a_27_47# 0 0.208f
C3553 VGND 0 23.9f
C3554 p[0] 0 0.808f
C3555 th01_0/m1_991_n1219# 0 1.24f
C3556 th01_0/m1_571_n501# 0 0.194f
C3557 th15_0/Vin 0 6.95f
C3558 _11_ 0 0.265f
C3559 _37_/a_27_47# 0 0.175f
C3560 net13 0 0.38f
C3561 input13/a_27_47# 0 0.208f
C3562 net18 0 0.207f
C3563 _25_ 0 0.191f
C3564 _54_/a_75_212# 0 0.21f
C3565 _38_/a_27_47# 0 0.175f
C3566 net19 0 0.165f
C3567 _22_ 0 0.215f
C3568 _14_ 0 0.225f
C3569 _15_ 0 0.331f
C3570 _55_/a_217_297# 0 0.00117f
C3571 _55_/a_80_21# 0 0.21f
C3572 input12/a_27_47# 0 0.208f
C3573 net9 0 0.285f
C3574 input9/a_75_212# 0 0.21f
C3575 _39_/a_285_47# 0 0.0174f
C3576 _39_/a_47_47# 0 0.199f
C3577 input11/a_27_47# 0 0.208f
C3578 net8 0 0.386f
C3579 input8/a_27_47# 0 0.208f
C3580 p[2] 0 0.487f
C3581 th03_0/m1_890_n844# 0 1.05f
C3582 th03_0/m1_638_n591# 0 0.224f
C3583 input10/a_27_47# 0 0.208f
C3584 net7 0 0.449f
C3585 input7/a_27_47# 0 0.208f
C3586 p[9] 0 0.698f
C3587 th10_0/m1_536_174# 0 0.825f
C3588 th10_0/m1_502_n495# 0 0.146f
C3589 input6/a_27_47# 0 0.208f
C3590 net5 0 0.817f
C3591 input5/a_841_47# 0 0.0929f
C3592 input5/a_664_47# 0 0.13f
C3593 input5/a_558_47# 0 0.164f
C3594 input5/a_381_47# 0 0.11f
C3595 input5/a_62_47# 0 0.169f
C3596 p[4] 0 0.515f
C3597 th05_0/m1_752_n794# 0 0.788f
C3598 input4/a_75_212# 0 0.21f
C3599 th12_0/m1_529_n42# 0 0.861f
C3600 p[11] 0 0.505f
C3601 th12_0/m1_394_n856# 0 0.215f
C3602 input3/a_27_47# 0 0.208f
C3603 net2 0 0.68f
C3604 input2/a_27_47# 0 0.208f
C3605 th07_0/m1_808_n892# 0 0.511f
C3606 p[6] 0 0.61f
C3607 net1 0 0.337f
C3608 input1/a_75_212# 0 0.21f
C3609 th14_0/m1_891_419# 0 1.48f
C3610 p[13] 0 0.763f
C3611 th14_0/m1_641_n318# 0 0.241f
C3612 b[3] 0 0.136f
C3613 output19/a_27_47# 0 0.543f
C3614 th09_0/m1_485_n505# 0 1.18f
C3615 p[8] 0 0.623f
C3616 th09_0/m1_962_372# 0 0.118f
C3617 b[2] 0 0.515f
C3618 output18/a_27_47# 0 0.543f
C3619 b[1] 0 0.204f
C3620 net17 0 0.169f
C3621 output17/a_27_47# 0 0.543f
C3622 _41_/a_59_75# 0 0.177f
C3623 b[0] 0 0.501f
C3624 output16/a_27_47# 0 0.543f
C3625 _16_ 0 0.125f
C3626 _42_/a_209_311# 0 0.143f
C3627 _42_/a_109_93# 0 0.158f
C3628 net6 0 0.533f
C3629 net4 0 0.315f
C3630 _26_/a_29_53# 0 0.18f
C3631 _43_/a_193_413# 0 0.136f
C3632 _43_/a_27_47# 0 0.224f
C3633 _01_ 0 0.15f
C3634 net14 0 0.502f
C3635 net3 0 0.453f
C3636 net15 0 0.446f
C3637 _27_/a_27_297# 0 0.163f
C3638 _18_ 0 0.143f
C3639 _17_ 0 0.242f
C3640 _44_/a_250_297# 0 0.0278f
C3641 _44_/a_93_21# 0 0.151f
C3642 net16 0 0.23f
C3643 _13_ 0 0.133f
C3644 _45_/a_193_297# 0 0.0011f
C3645 _45_/a_109_297# 0 7.11e-19
C3646 _45_/a_27_47# 0 0.216f
C3647 _00_ 0 0.377f
C3648 net11 0 0.762f
C3649 net12 0 0.512f
C3650 _29_/a_29_53# 0 0.18f
C3651 _19_ 0 0.113f
C3652 _04_ 0 0.334f
C3653 p[1] 0 0.451f
C3654 th02_0/m1_983_133# 0 1.44f
C3655 th02_0/m1_571_144# 0 0.252f
C3656 _47_/a_299_297# 0 0.0348f
C3657 _47_/a_81_21# 0 0.147f
C3658 VPWR 0 96f
C3659 _48_/a_27_47# 0 0.177f
C3660 _21_ 0 0.29f
C3661 _20_ 0 0.237f
C3662 _02_ 0 0.447f
C3663 _49_/a_201_297# 0 0.00345f
C3664 _49_/a_75_199# 0 0.205f
.ends

