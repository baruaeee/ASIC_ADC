magic
tech sky130A
magscale 1 2
timestamp 1702941821
<< checkpaint >>
rect -774 2329 2168 2374
rect -1313 2268 2168 2329
rect -1313 2107 3076 2268
rect -1313 -713 3445 2107
rect -1260 -925 3445 -713
rect -1260 -2460 1460 -925
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_WV9GCW  XM1
timestamp 0
transform 1 0 1151 0 1 702
box -296 -261 296 261
use sky130_fd_pr__nfet_01v8_KPA4J6  XM2
timestamp 0
transform 1 0 1974 0 1 591
box -211 -256 211 256
use sky130_fd_pr__nfet_01v8_648S5X  XM3
timestamp 0
transform 1 0 1605 0 1 698
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_WV9GCW  XM7
timestamp 0
transform 1 0 243 0 1 808
box -296 -261 296 261
use sky130_fd_pr__nfet_01v8_648S5X  XM10
timestamp 0
transform 1 0 697 0 1 804
box -211 -310 211 310
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
