magic
tech sky130A
magscale 1 2
timestamp 1706224144
<< error_p >>
rect -29 123 29 129
rect -29 89 -17 123
rect -29 83 29 89
rect -29 -89 29 -83
rect -29 -123 -17 -89
rect -29 -129 29 -123
<< nwell >>
rect -218 -261 218 261
<< pmos >>
rect -22 -42 22 42
<< pdiff >>
rect -80 30 -22 42
rect -80 -30 -68 30
rect -34 -30 -22 30
rect -80 -42 -22 -30
rect 22 30 80 42
rect 22 -30 34 30
rect 68 -30 80 30
rect 22 -42 80 -30
<< pdiffc >>
rect -68 -30 -34 30
rect 34 -30 68 30
<< nsubdiff >>
rect -148 191 -86 225
rect 86 191 148 225
<< nsubdiffcont >>
rect -86 191 86 225
<< poly >>
rect -33 123 33 139
rect -33 89 -17 123
rect 17 89 33 123
rect -33 73 33 89
rect -22 42 22 73
rect -22 -73 22 -42
rect -33 -89 33 -73
rect -33 -123 -17 -89
rect 17 -123 33 -89
rect -33 -139 33 -123
<< polycont >>
rect -17 89 17 123
rect -17 -123 17 -89
<< locali >>
rect -148 191 -86 225
rect 86 191 148 225
rect -33 89 -17 123
rect 17 89 33 123
rect -68 30 -34 46
rect -68 -46 -34 -30
rect 34 30 68 46
rect 34 -46 68 -30
rect -33 -123 -17 -89
rect 17 -123 33 -89
<< viali >>
rect -17 89 17 123
rect -68 -30 -34 30
rect 34 -30 68 30
rect -17 -123 17 -89
<< metal1 >>
rect -29 123 29 129
rect -29 89 -17 123
rect 17 89 29 123
rect -29 83 29 89
rect -74 30 -28 42
rect -74 -30 -68 30
rect -34 -30 -28 30
rect -74 -42 -28 -30
rect 28 30 74 42
rect 28 -30 34 30
rect 68 -30 74 30
rect 28 -42 74 -30
rect -29 -89 29 -83
rect -29 -123 -17 -89
rect 17 -123 29 -89
rect -29 -129 29 -123
<< properties >>
string FIXED_BBOX -165 -208 165 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.22 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
