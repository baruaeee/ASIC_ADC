VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO oaTaper STRING ;
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO div_fixed
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN div_fixed 0 0 ;
  SIZE 1.68 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
        RECT 0.275 -0.2 0.505 0.73 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT -0.095 2.335 0.345 3.715 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.185 1.045 1.515 2.805 ;
        RECT 0.495 1.045 1.515 1.735 ;
    END
  END Y
  OBS
    LAYER mcon ;
      RECT 1.265 2.605 1.435 2.775 ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.525 1.125 0.695 1.295 ;
      RECT 0.525 1.485 0.695 1.655 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.305 0.5 0.475 0.67 ;
      RECT 0.06 2.71 0.23 2.88 ;
      RECT 0.06 3.17 0.23 3.34 ;
  END
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END div_fixed

MACRO inv01f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv01f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.95 2.86 1.47 3.55 ;
        RECT 1.245 0.525 1.47 3.55 ;
        RECT 0.97 0.525 1.47 0.855 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.39 1.35 0.76 2.2 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 1 0.61 1.17 0.78 ;
      RECT 0.98 2.94 1.15 3.11 ;
      RECT 0.98 3.3 1.15 3.47 ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.49 1.545 0.66 1.715 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv01f

MACRO inv02f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv02f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.61 2.72 1.355 3.41 ;
        RECT 1.125 0.685 1.355 3.41 ;
        RECT 0.625 0.685 1.355 1.015 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.275 1.35 0.645 2.2 ;
    END
  END A
  OBS
    LAYER mcon ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.655 0.765 0.825 0.935 ;
      RECT 0.64 2.8 0.81 2.97 ;
      RECT 0.64 3.16 0.81 3.33 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 1.545 0.545 1.715 ;
      RECT 0.375 4.055 0.545 4.225 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv02f

MACRO inv03f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv03f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.705 2.81 1.49 3.5 ;
        RECT 1.26 0.665 1.49 3.5 ;
        RECT 0.685 0.665 1.49 1.355 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.325 1.675 0.695 2.045 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.735 2.89 0.905 3.06 ;
      RECT 0.735 3.25 0.905 3.42 ;
      RECT 0.715 0.745 0.885 0.915 ;
      RECT 0.715 1.105 0.885 1.275 ;
      RECT 0.425 1.775 0.595 1.945 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv03f

MACRO inv04f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv04f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.54 2.81 1.445 3.5 ;
        RECT 1.215 0.615 1.445 3.5 ;
        RECT 0.88 0.615 1.445 1.305 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.555 1.675 0.925 2.045 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 0.91 0.695 1.08 0.865 ;
      RECT 0.91 1.055 1.08 1.225 ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.655 1.775 0.825 1.945 ;
      RECT 0.57 2.89 0.74 3.06 ;
      RECT 0.57 3.25 0.74 3.42 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv04f

MACRO inv05f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv05f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.54 2.81 1.445 3.5 ;
        RECT 1.215 0.615 1.445 3.5 ;
        RECT 0.88 0.615 1.445 1.305 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.25 1.675 0.62 2.045 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 0.91 0.695 1.08 0.865 ;
      RECT 0.91 1.055 1.08 1.225 ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.57 2.89 0.74 3.06 ;
      RECT 0.57 3.25 0.74 3.42 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
      RECT 0.35 1.775 0.52 1.945 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv05f

MACRO inv06f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv06f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.37 2.135 0.74 2.505 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.795 3.12 1.44 3.45 ;
        RECT 1.21 0.69 1.44 3.45 ;
        RECT 0.74 0.69 1.44 1.38 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  OBS
    LAYER mcon ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.825 3.2 0.995 3.37 ;
      RECT 0.77 0.77 0.94 0.94 ;
      RECT 0.77 1.13 0.94 1.3 ;
      RECT 0.47 2.235 0.64 2.405 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv06f

MACRO inv07f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv07f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.54 3.07 1.34 3.4 ;
        RECT 1.11 0.595 1.34 3.4 ;
        RECT 0.64 0.595 1.34 1.285 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.25 2.135 0.62 2.505 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.67 0.675 0.84 0.845 ;
      RECT 0.67 1.035 0.84 1.205 ;
      RECT 0.57 3.15 0.74 3.32 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
      RECT 0.35 2.235 0.52 2.405 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv07f

MACRO inv08f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv08f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.55 2.825 1.2 3.515 ;
        RECT 0.87 1.755 1.2 3.515 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT -0.03 1.56 0.34 1.93 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 0.95 1.785 1.12 1.955 ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.58 2.905 0.75 3.075 ;
      RECT 0.58 3.265 0.75 3.435 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
      RECT 0.07 1.66 0.24 1.83 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv08f

MACRO inv09f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv09f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.505 2.19 1.435 2.45 ;
        RECT 0.505 1.82 0.835 2.45 ;
        RECT 0.575 1.82 0.805 3.39 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT -0.165 1.89 0.205 2.26 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.34 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.605 3.14 0.775 3.31 ;
      RECT 0.585 1.85 0.755 2.02 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
      RECT -0.065 1.99 0.105 2.16 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv09f

MACRO inv10f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv10f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.655 2.745 1.355 3.435 ;
        RECT 1.095 0.69 1.355 3.435 ;
        RECT 0.605 0.69 1.355 1.38 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.315 1.675 0.685 2.045 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.685 2.825 0.855 2.995 ;
      RECT 0.685 3.185 0.855 3.355 ;
      RECT 0.635 0.77 0.805 0.94 ;
      RECT 0.635 1.13 0.805 1.3 ;
      RECT 0.415 1.775 0.585 1.945 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv10f

MACRO inv11f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv11f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.635 2.7 1.45 3.39 ;
        RECT 1.19 0.745 1.45 3.39 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.295 1.58 0.665 1.95 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.34 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 1.22 0.825 1.39 0.995 ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.665 2.78 0.835 2.95 ;
      RECT 0.665 3.14 0.835 3.31 ;
      RECT 0.395 1.68 0.565 1.85 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv11f

MACRO inv12f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv12f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.56 2.825 1.185 3.515 ;
        RECT 0.925 0.62 1.185 3.515 ;
        RECT 0.695 0.62 1.185 1.31 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.28 2 0.65 2.37 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.725 0.7 0.895 0.87 ;
      RECT 0.725 1.06 0.895 1.23 ;
      RECT 0.59 2.885 0.76 3.055 ;
      RECT 0.59 3.245 0.76 3.415 ;
      RECT 0.38 2.1 0.55 2.27 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv12f

MACRO inv13f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv13f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.57 2.775 1.165 3.465 ;
        RECT 0.935 0.72 1.165 3.465 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.28 1.605 0.65 1.975 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 0.965 0.83 1.135 1 ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.6 2.855 0.77 3.025 ;
      RECT 0.6 3.215 0.77 3.385 ;
      RECT 0.38 1.705 0.55 1.875 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv13f

MACRO inv14f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv14f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.62 2.75 1.28 3.44 ;
        RECT 1.05 0.72 1.28 3.44 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.335 1.56 0.705 1.93 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.38 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 1.08 0.83 1.25 1 ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.65 2.83 0.82 3 ;
      RECT 0.65 3.19 0.82 3.36 ;
      RECT 0.435 1.66 0.605 1.83 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
  END
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
  PROPERTY CatenaDesignType "deviceLevel" ;
END inv14f

MACRO inv15f
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN inv15f 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.795 2.725 1.45 3.415 ;
        RECT 1.19 0.745 1.45 3.415 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.515 1.58 0.885 1.95 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.34 ;
    END
  END VDD
  OBS
    LAYER mcon ;
      RECT 1.22 0.825 1.39 0.995 ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.825 2.805 0.995 2.975 ;
      RECT 0.825 3.165 0.995 3.335 ;
      RECT 0.615 1.68 0.785 1.85 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END inv15f

MACRO preampF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN preampF 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT -0.125 3.94 1.38 4.38 ;
        RECT -0.125 0.47 0.245 1.52 ;
        RECT -0.125 0.47 0.075 4.38 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.23 1.855 0.6 2.705 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.955 0.47 1.245 3.685 ;
        RECT 0.455 0.47 1.245 1.52 ;
    END
  END Y
  OBS
    LAYER mcon ;
      RECT 1.015 3.485 1.185 3.655 ;
      RECT 0.835 -0.085 1.005 0.085 ;
      RECT 0.835 4.055 1.005 4.225 ;
      RECT 0.485 0.55 0.655 0.72 ;
      RECT 0.485 0.91 0.655 1.08 ;
      RECT 0.485 1.27 0.655 1.44 ;
      RECT 0.375 -0.085 0.545 0.085 ;
      RECT 0.375 4.055 0.545 4.225 ;
      RECT 0.33 2.05 0.5 2.22 ;
      RECT 0.045 0.55 0.215 0.72 ;
      RECT 0.045 0.91 0.215 1.08 ;
      RECT 0.045 1.27 0.215 1.44 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
  PROPERTY oaTaper "virtuosoDefaultSetup" ;
END preampF

MACRO preampF_comm_B
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN preampF_comm_B 0 0 ;
  SIZE 1.38 BY 4.14 ;
  SYMMETRY X Y ;
  SITE MACRO ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 3.94 1.38 4.34 ;
        RECT 0 2.735 0.31 3.785 ;
        RECT 0 2.735 0.165 4.34 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.13 2.19 0.78 2.56 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0 -0.2 1.38 0.2 ;
        RECT 0.24 -0.2 0.57 0.645 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.51 2.735 0.74 3.785 ;
    END
  END Y
  OBS
    LAYER mcon ;
      RECT 1.08 0.57 1.25 0.74 ;
      RECT 1.08 0.93 1.25 1.1 ;
      RECT 1.08 1.29 1.25 1.46 ;
      RECT 1.08 1.65 1.25 1.82 ;
      RECT 1.08 2.995 1.25 3.165 ;
      RECT 1.08 3.355 1.25 3.525 ;
      RECT 0.54 2.815 0.71 2.985 ;
      RECT 0.54 3.175 0.71 3.345 ;
      RECT 0.54 3.535 0.71 3.705 ;
      RECT 0.325 2.29 0.495 2.46 ;
      RECT 0.32 0.445 0.49 0.615 ;
      RECT 0.11 2.815 0.28 2.985 ;
      RECT 0.11 3.175 0.28 3.345 ;
      RECT 0.11 3.535 0.28 3.705 ;
    LAYER met1 ;
      RECT 1.03 0.415 1.3 1.975 ;
      RECT 1.03 2.75 1.3 3.77 ;
  END
END preampF_comm_B

END LIBRARY
