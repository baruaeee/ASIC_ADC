magic
tech sky130A
magscale 1 2
timestamp 1706270854
<< psubdiff >>
rect 710 -1088 807 -1054
<< locali >>
rect 451 78 493 112
rect 707 -1088 767 -1054
rect 801 -1088 825 -1054
<< viali >>
rect 417 78 451 112
rect 981 -156 1015 -122
rect 767 -1088 801 -1054
<< metal1 >>
rect 411 113 457 124
rect 399 112 461 113
rect 399 78 417 112
rect 451 79 461 112
rect 451 78 457 79
rect 399 66 457 78
rect 399 -209 433 66
rect 616 53 668 59
rect 952 48 1052 148
rect 616 -5 668 1
rect 504 -98 556 -36
rect 399 -243 513 -209
rect 479 -485 513 -243
rect 479 -543 545 -485
rect 620 -488 654 -97
rect 728 -124 734 -72
rect 786 -124 792 -72
rect 979 -110 1013 48
rect 975 -122 1021 -110
rect 975 -156 981 -122
rect 1015 -156 1021 -122
rect 975 -168 1021 -156
rect 979 -328 1013 -168
rect 1088 -214 1150 -212
rect 1086 -262 1150 -214
rect 1086 -264 1148 -262
rect 979 -362 1084 -328
rect 1151 -371 1293 -337
rect 1052 -434 1104 -428
rect 707 -542 741 -485
rect 1104 -486 1133 -435
rect 1052 -492 1133 -486
rect 650 -543 741 -542
rect 479 -577 741 -543
rect 1099 -643 1133 -492
rect 1259 -622 1293 -371
rect 489 -677 1133 -643
rect 489 -701 523 -677
rect 457 -735 523 -701
rect 906 -681 1133 -677
rect 457 -842 491 -735
rect 566 -758 572 -706
rect 624 -758 630 -706
rect 906 -795 940 -681
rect 1234 -722 1334 -622
rect 457 -876 562 -842
rect 631 -890 894 -856
rect 1259 -860 1293 -722
rect 376 -954 476 -910
rect 376 -988 615 -954
rect 376 -1010 476 -988
rect 771 -1042 805 -890
rect 954 -894 1293 -860
rect 892 -998 954 -944
rect 761 -1054 807 -1042
rect 761 -1088 767 -1054
rect 801 -1085 807 -1054
rect 1154 -1085 1254 -1022
rect 801 -1088 1254 -1085
rect 761 -1100 1254 -1088
rect 771 -1119 1254 -1100
rect 1154 -1122 1254 -1119
<< via1 >>
rect 616 1 668 53
rect 734 -124 786 -72
rect 1052 -486 1104 -434
rect 572 -758 624 -706
<< metal2 >>
rect 610 1 616 53
rect 668 44 674 53
rect 668 10 923 44
rect 668 1 674 10
rect 734 -72 786 -66
rect 734 -130 786 -124
rect 743 -187 777 -130
rect 743 -221 844 -187
rect 810 -693 844 -221
rect 889 -443 923 10
rect 1046 -443 1052 -434
rect 889 -477 1052 -443
rect 1046 -486 1052 -477
rect 1104 -486 1110 -434
rect 581 -700 844 -693
rect 572 -706 844 -700
rect 624 -727 844 -706
rect 572 -764 624 -758
use sky130_fd_pr__nfet_01v8_42G4RD  XM0
timestamp 1706224144
transform 1 0 596 0 1 -872
box -218 -252 218 252
use sky130_fd_pr__pfet_01v8_DDPLQ8  XM1
timestamp 1706224144
transform 0 -1 641 1 0 -67
box -215 -261 215 261
use sky130_fd_pr__nfet_01v8_VWP3K3  XM2
timestamp 1706224144
transform 0 -1 626 1 0 -515
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_LZD9A4  XM3
timestamp 1706224144
transform 1 0 1118 0 1 -347
box -218 -261 218 261
use sky130_fd_pr__nfet_01v8_VRD6K3  XM4
timestamp 1706224144
transform 1 0 923 0 1 -874
box -215 -252 215 252
<< labels >>
flabel metal1 1154 -1122 1254 -1022 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 1234 -722 1334 -622 0 FreeSans 256 0 0 0 V04
port 1 nsew
flabel metal1 952 48 1052 148 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 376 -1010 476 -910 0 FreeSans 256 0 0 0 Vin
port 2 nsew
<< end >>
