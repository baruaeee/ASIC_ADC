magic
tech sky130A
magscale 1 2
timestamp 1705195269
<< error_s >>
rect -8720 -8186 -8696 -8054
rect -8660 -8126 -8636 -8054
<< locali >>
rect -9082 -1852 -9034 -1784
<< viali >>
rect -9082 -1888 -9034 -1852
<< metal1 >>
rect -2393 1473 -2341 1479
rect -9426 1421 -2393 1470
rect -9426 480 -9377 1421
rect -2393 1412 -2341 1418
rect -3707 988 -3626 1078
rect -3707 958 -3693 988
rect -6831 909 -3693 958
rect -3641 909 -3626 988
rect -6831 908 -3626 909
rect -6831 903 -3641 908
rect -6831 900 -3647 903
rect -2666 250 -2466 450
rect -2619 222 -2491 250
rect -2619 138 -2533 222
rect -2673 132 -2533 138
rect -2683 55 -2673 130
rect -2619 55 -2533 132
rect -2673 47 -2619 53
rect -2501 -72 -2438 -66
rect -2438 -135 -2303 -72
rect -2501 -141 -2438 -135
rect -1995 -142 -1932 629
rect -2001 -205 -1995 -142
rect -1932 -205 -1926 -142
rect -1854 -359 -1848 -296
rect -1785 -359 -1779 -296
rect -9639 -472 -9121 -414
rect -9639 -1849 -9581 -472
rect -1848 -521 -1785 -359
rect -5182 -616 -5124 -610
rect -5124 -678 -4089 -620
rect -5182 -687 -5124 -681
rect -3496 -1368 -3296 -1168
rect -1847 -1252 -1784 -1036
rect -1847 -1315 -1533 -1252
rect -3418 -1652 -3354 -1368
rect -1906 -1542 -1900 -1506
rect -1976 -1570 -1900 -1542
rect -1836 -1570 -1830 -1506
rect -1976 -1642 -1836 -1570
rect -8697 -1745 -7715 -1687
rect -3424 -1716 -3418 -1652
rect -3354 -1716 -3348 -1652
rect -1968 -1682 -1836 -1642
rect -7773 -1831 -7715 -1745
rect -2788 -1812 -2724 -1766
rect -11037 -1907 -9581 -1849
rect -11037 -2165 -10979 -1907
rect -10091 -1975 -10085 -1971
rect -10588 -2033 -10085 -1975
rect -10588 -2287 -10530 -2033
rect -10091 -2039 -10085 -2033
rect -10017 -2039 -10011 -1971
rect -9639 -2483 -9581 -1907
rect -9094 -1852 -9022 -1846
rect -9094 -1888 -9082 -1852
rect -9034 -1860 -9022 -1852
rect -9034 -1888 -9020 -1860
rect -9094 -1912 -9020 -1888
rect -7773 -1889 -7293 -1831
rect -9368 -1971 -9316 -1965
rect -9368 -2044 -9316 -2039
rect -9094 -1973 -9029 -1912
rect -7351 -1967 -7293 -1889
rect -2898 -1962 -2724 -1812
rect -2844 -1970 -2724 -1962
rect -9094 -2003 -8940 -1973
rect -7822 -1981 -7764 -1975
rect -8158 -1985 -7958 -1984
rect -9094 -2044 -8924 -2003
rect -8158 -2043 -7822 -1985
rect -9368 -2045 -9029 -2044
rect -9360 -2080 -9029 -2045
rect -9360 -2446 -9324 -2080
rect -8158 -2184 -7958 -2043
rect -7822 -2052 -7764 -2046
rect -9639 -2541 -9177 -2483
rect -10068 -2718 -9868 -2646
rect -8530 -2709 -8330 -2648
rect -10068 -2776 -9830 -2718
rect -9762 -2776 -9756 -2718
rect -8530 -2734 -8170 -2709
rect -10068 -2846 -9868 -2776
rect -8530 -2792 -8290 -2734
rect -8170 -2792 -8164 -2734
rect -8530 -2817 -8170 -2792
rect -8530 -2848 -8330 -2817
rect -8604 -3104 -7388 -3068
rect -8604 -3336 -8568 -3104
rect -8864 -3372 -8568 -3336
rect -10150 -3842 -8748 -3806
rect -1751 -5475 -1688 -5469
rect -1596 -5475 -1533 -1315
rect -9576 -5700 -9376 -5500
rect -8104 -5684 -7904 -5484
rect -1688 -5538 -1533 -5475
rect -1418 -5516 -1348 -5506
rect -1751 -5544 -1688 -5538
rect -1418 -5570 -1410 -5516
rect -1354 -5570 -1348 -5516
rect -1418 -5608 -1348 -5570
rect -2563 -5735 -2557 -5712
rect -2572 -5764 -2557 -5735
rect -2505 -5764 -2499 -5712
rect -2572 -5776 -2507 -5764
rect -2689 -5827 -2507 -5776
rect -10006 -6114 -9806 -5914
rect -2051 -5981 -2045 -5911
rect -1975 -5973 -1969 -5911
rect -1975 -5981 -1907 -5973
rect -2045 -6079 -1907 -5981
rect -813 -5992 -722 -5938
rect -666 -5992 -660 -5938
rect -9945 -6172 -9883 -6114
rect -9952 -6234 -9946 -6172
rect -9882 -6234 -9876 -6172
rect -10900 -6500 -10700 -6300
rect -9776 -6374 -9576 -6174
rect -1737 -6192 -1683 -6186
rect -1811 -6246 -1737 -6192
rect -1737 -6252 -1683 -6246
rect -900 -6300 -700 -6100
rect -1541 -6667 -1471 -6653
rect -1457 -6667 -1205 -6653
rect -1541 -6723 -1205 -6667
rect -1541 -6740 -1387 -6723
rect -10560 -6896 -10554 -6836
rect -10490 -6896 -10484 -6836
rect -10552 -6938 -10492 -6896
rect -10642 -6998 -10492 -6938
rect -10259 -7038 -10221 -6855
rect -10272 -7090 -10266 -7038
rect -10214 -7090 -10208 -7038
rect -5069 -7271 -2635 -7200
rect -4566 -7486 -4495 -7271
rect -10272 -7544 -10266 -7492
rect -10214 -7544 -10208 -7492
rect -10259 -7637 -10221 -7544
rect -4566 -7557 -3849 -7486
rect -3920 -7881 -3849 -7557
rect -1910 -7568 -1710 -7550
rect -1910 -7569 -1768 -7568
rect -1931 -7619 -1768 -7569
rect -1910 -7620 -1768 -7619
rect -1712 -7620 -1706 -7568
rect -3014 -7732 -3008 -7656
rect -2932 -7732 -2856 -7656
rect -1910 -7750 -1710 -7620
rect -9458 -8012 -9397 -8007
rect -9462 -8064 -9456 -8012
rect -9400 -8064 -9394 -8012
rect -9458 -8150 -9397 -8064
rect -9532 -8350 -9332 -8150
rect -1541 -8305 -1471 -6740
rect -1143 -6775 -1073 -6769
rect -1073 -6839 -937 -6780
rect -1143 -6851 -1073 -6845
rect -996 -6951 -937 -6839
rect -378 -7863 -170 -7798
rect -2233 -8375 -1460 -8305
rect -2544 -8410 -2296 -8380
rect -3020 -8462 -2256 -8410
rect -9982 -8588 -9946 -8560
rect -10010 -8702 -9946 -8588
rect -9306 -8644 -8716 -8643
rect -9306 -8720 -8568 -8644
rect -9306 -8726 -8502 -8720
rect -5618 -8722 -5418 -8522
rect -3378 -8552 -3178 -8512
rect -3378 -8604 -3124 -8552
rect -3072 -8604 -3066 -8552
rect -3378 -8712 -3178 -8604
rect -9306 -8782 -8554 -8726
rect -9306 -8788 -8502 -8782
rect -9306 -8843 -8568 -8788
rect -3020 -8804 -2968 -8462
rect -1042 -8566 -842 -8474
rect -1042 -8650 -992 -8566
rect -908 -8650 -842 -8566
rect -1042 -8674 -842 -8650
rect -8768 -8844 -8568 -8843
rect -3208 -8856 -2968 -8804
rect -235 -8830 -170 -7863
rect -4779 -8939 -4579 -8931
rect -4787 -8991 -4781 -8939
rect -4711 -8991 -4579 -8939
rect -4779 -8998 -4579 -8991
rect -10028 -9422 -9964 -9392
rect -10028 -9599 -9920 -9422
rect -8943 -9488 -8937 -9436
rect -8881 -9488 -8875 -9436
rect -8354 -9524 -8318 -9252
rect -3208 -9340 -3156 -8856
rect -1447 -8895 -170 -8830
rect -1888 -8981 -1688 -8946
rect -1888 -8987 -1641 -8981
rect -1888 -9039 -1693 -8987
rect -1888 -9045 -1641 -9039
rect -3017 -9100 -3011 -9048
rect -2955 -9100 -2848 -9048
rect -1888 -9146 -1688 -9045
rect -4288 -9524 -4252 -9368
rect -3540 -9392 -3156 -9340
rect -8354 -9560 -4252 -9524
rect -10028 -9605 -9907 -9599
rect -10028 -9670 -9959 -9605
rect -3348 -9603 -3296 -9597
rect -9907 -9670 -9901 -9606
rect -3354 -9671 -3348 -9606
rect -9959 -9677 -9907 -9671
rect -1447 -9606 -1382 -8895
rect -3296 -9671 -1382 -9606
rect -3348 -9682 -3296 -9676
<< via1 >>
rect -2393 1418 -2341 1473
rect -3693 909 -3641 988
rect -2673 53 -2619 132
rect -2501 -135 -2438 -72
rect -1995 -205 -1932 -142
rect -1848 -359 -1785 -296
rect -5182 -681 -5124 -616
rect -1900 -1570 -1836 -1506
rect -3418 -1716 -3354 -1652
rect -10085 -2039 -10017 -1971
rect -9368 -2039 -9316 -1971
rect -7822 -2046 -7764 -1981
rect -9830 -2776 -9762 -2718
rect -8290 -2792 -8170 -2734
rect -1751 -5538 -1688 -5475
rect -1410 -5570 -1354 -5516
rect -2557 -5764 -2505 -5712
rect -2045 -5981 -1975 -5911
rect -722 -5992 -666 -5938
rect -9946 -6234 -9882 -6172
rect -1737 -6246 -1683 -6192
rect -10554 -6896 -10490 -6836
rect -10266 -7090 -10214 -7038
rect -10266 -7544 -10214 -7492
rect -1768 -7620 -1712 -7568
rect -3008 -7732 -2932 -7656
rect -9456 -8064 -9400 -8012
rect -1143 -6845 -1073 -6775
rect -3124 -8604 -3072 -8552
rect -8554 -8782 -8502 -8726
rect -992 -8650 -908 -8566
rect -4781 -8991 -4711 -8939
rect -8937 -9488 -8881 -9436
rect -1693 -9039 -1641 -8987
rect -3011 -9100 -2955 -9048
rect -9959 -9671 -9907 -9605
rect -3348 -9676 -3296 -9603
<< metal2 >>
rect -2399 1418 -2393 1473
rect -2341 1418 -1793 1473
rect -3764 988 -3695 992
rect -3769 983 -3693 988
rect -3769 914 -3764 983
rect -3695 914 -3693 983
rect -3769 909 -3693 914
rect -3641 909 -3635 988
rect -3764 905 -3695 909
rect -2841 53 -2673 132
rect -2619 53 -2613 132
rect -2554 -72 -2498 -67
rect -2554 -76 -2501 -72
rect -2554 -135 -2501 -132
rect -2438 -135 -2432 -72
rect -2554 -141 -2498 -135
rect -1995 -142 -1932 -136
rect -1995 -211 -1932 -205
rect -5993 -681 -5182 -616
rect -5124 -681 -5118 -616
rect -1986 -620 -1942 -211
rect -1848 -241 -1793 1418
rect -1848 -296 -1785 -241
rect -1848 -365 -1785 -359
rect -1986 -664 -1846 -620
rect -5993 -1616 -5928 -681
rect -1890 -1500 -1846 -664
rect -1900 -1506 -1836 -1500
rect -1900 -1576 -1836 -1570
rect -7575 -1681 -5928 -1616
rect -3418 -1652 -3354 -1646
rect -10085 -1971 -10017 -1965
rect -10017 -2039 -9368 -1971
rect -9316 -2039 -9310 -1971
rect -7575 -1981 -7510 -1681
rect -3418 -1722 -3354 -1716
rect -3414 -1852 -3358 -1722
rect -7828 -1982 -7822 -1981
rect -10085 -2045 -10017 -2039
rect -7870 -2046 -7822 -1982
rect -7764 -2046 -7510 -1981
rect -7870 -2089 -7510 -2046
rect -7575 -2154 -7510 -2089
rect -9830 -2718 -9762 -2712
rect -9830 -3898 -9762 -2776
rect -8290 -2734 -8170 -2548
rect -8290 -2798 -8170 -2792
rect -9830 -3966 -8288 -3898
rect -1476 -5416 -666 -5360
rect -1757 -5482 -1751 -5475
rect -2035 -5532 -1751 -5482
rect -2564 -5684 -2555 -5628
rect -2499 -5684 -2490 -5628
rect -2564 -5712 -2491 -5684
rect -2564 -5762 -2557 -5712
rect -2505 -5762 -2491 -5712
rect -2557 -5770 -2505 -5764
rect -2035 -5905 -1985 -5532
rect -1757 -5538 -1751 -5532
rect -1688 -5538 -1682 -5475
rect -1419 -5508 -1410 -5452
rect -1354 -5508 -1345 -5452
rect -1410 -5516 -1354 -5508
rect -1410 -5576 -1354 -5570
rect -2045 -5911 -1975 -5905
rect -2045 -5987 -1975 -5981
rect -722 -5938 -666 -5416
rect -722 -5998 -666 -5992
rect -9946 -6172 -9882 -6166
rect -9946 -6298 -9882 -6234
rect -1743 -6246 -1737 -6192
rect -1683 -6246 -1363 -6192
rect -10554 -6362 -9882 -6298
rect -10554 -6836 -10490 -6362
rect -1417 -6783 -1363 -6246
rect -1149 -6783 -1143 -6775
rect -1417 -6837 -1143 -6783
rect -1149 -6845 -1143 -6837
rect -1073 -6845 -1067 -6775
rect -10554 -6902 -10490 -6896
rect -10266 -7038 -10214 -7032
rect -10266 -7096 -10214 -7090
rect -10264 -7486 -10216 -7096
rect -10266 -7492 -10214 -7486
rect -10266 -7550 -10214 -7544
rect -1768 -7568 -1712 -6916
rect -3000 -7617 -2940 -7615
rect -9456 -8012 -9400 -7638
rect -3010 -7656 -3001 -7617
rect -2939 -7656 -2930 -7617
rect -1768 -7626 -1712 -7620
rect -3010 -7673 -3008 -7656
rect -2932 -7673 -2930 -7656
rect -3008 -7738 -2932 -7732
rect -9456 -8070 -9400 -8064
rect -3122 -8546 -3074 -8466
rect -3124 -8552 -3072 -8546
rect -3124 -8610 -3072 -8604
rect -992 -8566 -908 -8560
rect -992 -8656 -908 -8650
rect -978 -8676 -922 -8656
rect -8560 -8782 -8554 -8726
rect -8502 -8782 -8456 -8726
rect -4781 -8887 -4711 -8880
rect -4786 -8939 -4777 -8887
rect -4715 -8939 -4706 -8887
rect -4786 -8943 -4781 -8939
rect -4711 -8943 -4706 -8939
rect -4781 -8997 -4711 -8991
rect -3011 -8967 -2955 -8958
rect -3011 -9048 -2955 -9029
rect -1699 -8987 -1637 -8905
rect -1699 -9039 -1693 -8987
rect -1641 -9039 -1635 -8987
rect -3011 -9106 -2955 -9100
rect -8937 -9339 -8881 -9330
rect -8881 -9401 -8490 -9381
rect -8937 -9436 -8490 -9401
rect -8881 -9454 -8490 -9436
rect -8937 -9494 -8881 -9488
rect -9901 -9605 -9845 -9598
rect -8563 -9603 -8490 -9454
rect -9965 -9671 -9959 -9605
rect -9907 -9607 -9840 -9605
rect -9907 -9669 -9901 -9607
rect -9845 -9669 -9840 -9607
rect -9907 -9671 -9840 -9669
rect -9901 -9678 -9845 -9671
rect -8563 -9676 -3348 -9603
rect -3296 -9676 -3290 -9603
<< via2 >>
rect -3764 914 -3695 983
rect -2554 -132 -2501 -76
rect -2501 -132 -2498 -76
rect -2555 -5684 -2499 -5628
rect -1410 -5508 -1354 -5452
rect -3001 -7656 -2939 -7617
rect -3001 -7673 -2939 -7656
rect -4777 -8939 -4715 -8887
rect -4777 -8943 -4715 -8939
rect -3011 -9029 -2955 -8967
rect -8937 -9401 -8881 -9339
rect -9901 -9669 -9845 -9607
<< metal3 >>
rect -3770 983 -3638 994
rect -3770 914 -3764 983
rect -3695 981 -3638 983
rect -3695 917 -3658 981
rect -3594 917 -3588 981
rect -3695 914 -3638 917
rect -3770 902 -3638 914
rect -2559 -72 -2493 -71
rect -2559 -74 -2502 -72
rect -2594 -76 -2502 -74
rect -2594 -132 -2554 -76
rect -2594 -134 -2502 -132
rect -2559 -136 -2502 -134
rect -2438 -136 -2432 -72
rect -2559 -137 -2493 -136
rect -2558 -5301 -1351 -5239
rect -2558 -5623 -2496 -5301
rect -1413 -5447 -1351 -5301
rect -1415 -5452 -1349 -5447
rect -1415 -5508 -1410 -5452
rect -1354 -5508 -1349 -5452
rect -1415 -5513 -1349 -5508
rect -2560 -5628 -2494 -5623
rect -2560 -5684 -2555 -5628
rect -2499 -5684 -2494 -5628
rect -2560 -5689 -2494 -5684
rect -9194 -7560 -8984 -7488
rect -9056 -9334 -8984 -7560
rect -4782 -7604 -2934 -7532
rect -9056 -9339 -8876 -9334
rect -9056 -9401 -8937 -9339
rect -8881 -9401 -8876 -9339
rect -9056 -9406 -8876 -9401
rect -8768 -9602 -8696 -8054
rect -8660 -8126 -8412 -8054
rect -8484 -8202 -8412 -8126
rect -4782 -8202 -4710 -7604
rect -8484 -8274 -4710 -8202
rect -4782 -8887 -4710 -8274
rect -4782 -8943 -4777 -8887
rect -4715 -8943 -4710 -8887
rect -4782 -8948 -4710 -8943
rect -3016 -7617 -2934 -7604
rect -3016 -7673 -3001 -7617
rect -2939 -7673 -2934 -7617
rect -3016 -7678 -2934 -7673
rect -3016 -8967 -2944 -7678
rect -3016 -9029 -3011 -8967
rect -2955 -9029 -2944 -8967
rect -3016 -9034 -2944 -9029
rect -9906 -9607 -8696 -9602
rect -9906 -9669 -9901 -9607
rect -9845 -9669 -8696 -9607
rect -9906 -9674 -8696 -9669
<< via3 >>
rect -3658 917 -3594 981
rect -2502 -76 -2438 -72
rect -2502 -132 -2498 -76
rect -2498 -132 -2438 -76
rect -2502 -136 -2438 -132
<< metal4 >>
rect -3659 981 -3593 982
rect -3659 978 -3658 981
rect -3702 917 -3658 978
rect -3594 917 -3593 981
rect -3702 916 -3593 917
rect -3702 -74 -3642 916
rect -2503 -72 -2437 -71
rect -2503 -74 -2502 -72
rect -3702 -134 -2502 -74
rect -3702 -1636 -3642 -134
rect -2503 -136 -2502 -134
rect -2438 -136 -2437 -72
rect -2503 -137 -2437 -136
rect -5648 -1696 -3642 -1636
rect -5648 -1956 -5588 -1696
use th10  th10_0
timestamp 1705011335
transform 1 0 -10072 0 1 -2690
box 394 -1164 1590 790
use th02  x16
timestamp 1705010589
transform 1 0 -9326 0 1 -7538
box 1100 -1960 4395 680
use th03  x17
timestamp 1705010624
transform 1 0 -5078 0 1 -8488
box 414 -920 1840 706
use th04  x18
timestamp 1705010641
transform 0 1 -9286 1 0 -9859
box 279 -1300 1216 476
use th05  x19
timestamp 1705010690
transform 0 1 -522 -1 0 -6476
box 394 -966 2064 258
use th06  x20
timestamp 1705011040
transform 1 0 -2290 0 1 -5634
box 308 -1110 1542 62
use th07  x21
timestamp 1705011056
transform 1 0 -3192 0 -1 -9724
box 296 -1290 1462 -44
use th08  x22
timestamp 1705011074
transform 1 0 -3240 0 1 -7076
box 330 -1392 1396 54
use th09  x23
timestamp 1705011303
transform 0 -1 -3310 -1 0 2098
box 670 -1498 1918 398
use th11  x25
timestamp 1705011594
transform 0 -1 -8772 1 0 -7714
box 160 -636 1584 1464
use th12  x26
timestamp 1705011684
transform 1 0 -11565 0 1 -2790
box 375 -1092 1662 716
use th13  x27
timestamp 1705099334
transform -1 0 -1434 0 1 -630
box 240 -1200 2062 556
use th14  x28
timestamp 1705011828
transform 1 0 -12106 0 1 -4884
box 300 -1200 4172 772
use th15  x29
timestamp 1705104586
transform 1 0 -10387 0 1 -904
box 915 -950 6436 1862
use preamp  x30
timestamp 1705010541
transform 1 0 -12008 0 1 -7081
box 398 -255 1470 780
use th01  x31
timestamp 1705010572
transform 1 0 -12168 0 1 -7430
box 618 -1168 2664 -180
<< labels >>
flabel metal1 -9576 -5700 -9376 -5500 0 FreeSans 256 0 0 0 Vin
port 0 nsew
flabel metal1 -3496 -1368 -3296 -1168 0 FreeSans 256 0 0 0 V13
port 14 nsew
flabel metal1 -8158 -2184 -7958 -1984 0 FreeSans 256 0 0 0 V15
port 16 nsew
flabel metal1 -8530 -2848 -8330 -2648 0 FreeSans 256 0 0 0 V10
port 11 nsew
flabel metal1 -10068 -2846 -9868 -2646 0 FreeSans 256 0 0 0 V12
port 13 nsew
flabel metal1 -8104 -5684 -7904 -5484 0 FreeSans 256 0 0 0 V14
port 15 nsew
flabel metal1 -9776 -6374 -9576 -6174 0 FreeSans 256 0 0 0 V11
port 12 nsew
flabel metal1 -9532 -8350 -9332 -8150 0 FreeSans 256 0 0 0 V1
port 2 nsew
flabel metal1 -5618 -8722 -5418 -8522 0 FreeSans 256 0 0 0 V2
port 3 nsew
flabel metal1 -3378 -8712 -3178 -8512 0 FreeSans 256 0 0 0 V3
port 4 nsew
flabel metal1 -8768 -8844 -8568 -8644 0 FreeSans 256 0 0 0 V4
port 5 nsew
flabel metal1 -1910 -7750 -1710 -7550 0 FreeSans 256 0 0 0 V8
port 9 nsew
flabel metal1 -1888 -9146 -1688 -8946 0 FreeSans 256 0 0 0 V7
port 8 nsew
flabel metal1 -900 -6300 -700 -6100 0 FreeSans 256 0 0 0 V6
port 7 nsew
flabel metal1 -1042 -8674 -842 -8474 0 FreeSans 256 0 0 0 V5
port 6 nsew
flabel metal1 -2666 250 -2466 450 0 FreeSans 256 0 0 0 V9
port 10 nsew
flabel metal1 -10900 -6500 -10700 -6300 0 FreeSans 256 0 0 0 Vp
port 1 nsew
flabel metal1 -10006 -6114 -9806 -5914 0 FreeSans 256 0 0 0 Vn
port 17 nsew
<< end >>
