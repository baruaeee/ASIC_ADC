magic
tech sky130A
magscale 1 2
timestamp 1706466859
<< nwell >>
rect 2878 -1714 3806 -1488
rect 3808 -1708 4222 -1544
rect 4646 -1708 4894 -1528
rect 3808 -1714 4894 -1708
rect 2878 -1754 4894 -1714
rect 2878 -1756 3866 -1754
rect 2878 -1768 3824 -1756
rect 2878 -1840 3806 -1768
rect 4214 -1796 4894 -1754
rect 4214 -1912 4890 -1796
<< pwell >>
rect 4210 -758 4260 -696
<< metal1 >>
rect 1766 -545 4843 -511
rect 3028 -598 3072 -545
rect 5118 -559 5218 -528
rect 4957 -593 5443 -559
rect 1538 -1162 1638 -1062
rect 1585 -1327 1619 -1162
rect 2945 -3851 2979 -1651
rect 3028 -1871 3065 -598
rect 5118 -628 5218 -593
rect 4156 -698 4256 -660
rect 4156 -702 4308 -698
rect 4156 -754 4209 -702
rect 4261 -754 4308 -702
rect 4156 -758 4308 -754
rect 4156 -760 4256 -758
rect 5409 -769 5443 -593
rect 5144 -1135 5244 -1092
rect 4943 -1169 5244 -1135
rect 5144 -1192 5244 -1169
rect 4056 -1272 4108 -1266
rect 4056 -1330 4108 -1324
rect 3138 -1355 3190 -1349
rect 3138 -1413 3190 -1407
rect 5340 -1354 5417 -1295
rect 5340 -1391 5420 -1354
rect 5340 -1392 5404 -1391
rect 3028 -1877 3100 -1871
rect 3028 -1929 3048 -1877
rect 3028 -1935 3100 -1929
rect 3028 -1936 3065 -1935
rect 2831 -3885 2979 -3851
rect 3159 -3095 3193 -1445
rect 3581 -1591 3615 -1545
rect 3357 -1625 3615 -1591
rect 4822 -1604 4834 -1598
rect 3357 -1998 3391 -1625
rect 4814 -1636 4862 -1604
rect 4786 -1669 4886 -1636
rect 5340 -1669 5377 -1392
rect 4217 -1703 5377 -1669
rect 4786 -1736 4886 -1703
rect 3457 -1859 4085 -1825
rect 3342 -2050 3348 -1998
rect 3400 -2050 3406 -1998
rect 3457 -2777 3491 -1859
rect 3566 -2328 3572 -2276
rect 3624 -2315 3878 -2276
rect 3624 -2328 3630 -2315
rect 5064 -2360 5164 -2324
rect 4956 -2416 5286 -2360
rect 5064 -2424 5164 -2416
rect 5230 -2772 5286 -2416
rect 3389 -2811 3491 -2777
rect 3389 -2906 3423 -2811
rect 3373 -2958 3379 -2906
rect 3431 -2958 3437 -2906
rect 5315 -3005 5407 -2971
rect 5315 -3025 5349 -3005
rect 4624 -3059 5349 -3025
rect 3614 -3072 3786 -3059
rect 3159 -3129 3601 -3095
rect 3614 -3116 3788 -3072
rect 3627 -3122 3788 -3116
rect 2831 -6465 2865 -3885
rect 3159 -3955 3193 -3129
rect 4920 -3600 5020 -3500
rect 4931 -3687 4965 -3600
rect 4781 -3721 4965 -3687
rect 2917 -3989 3193 -3955
rect 2917 -5817 2951 -3989
rect 3512 -4150 3564 -4144
rect 3512 -4208 3564 -4202
rect 4112 -5022 4212 -4922
rect 3192 -5114 3244 -5108
rect 3192 -5172 3244 -5166
rect 3874 -5508 3911 -5490
rect 3012 -5596 3018 -5544
rect 3070 -5545 3076 -5544
rect 3863 -5545 3911 -5508
rect 3070 -5582 3954 -5545
rect 3070 -5596 3076 -5582
rect 3824 -5586 3911 -5582
rect 2917 -5851 3283 -5817
rect 4740 -6440 4840 -6340
rect 2831 -6499 3377 -6465
<< via1 >>
rect 4209 -754 4261 -702
rect 4056 -1324 4108 -1272
rect 3138 -1407 3190 -1355
rect 3048 -1929 3100 -1877
rect 3348 -2050 3400 -1998
rect 3572 -2328 3624 -2276
rect 3379 -2958 3431 -2906
rect 3512 -4202 3564 -4150
rect 3192 -5166 3244 -5114
rect 3018 -5596 3070 -5544
<< metal2 >>
rect 4209 -702 4261 -696
rect 4209 -760 4261 -754
rect 4218 -869 4252 -760
rect 4137 -902 4252 -869
rect 4137 -906 4188 -902
rect 4137 -1263 4186 -906
rect 4098 -1272 4186 -1263
rect 4050 -1324 4056 -1272
rect 4108 -1315 4186 -1272
rect 4108 -1324 4114 -1315
rect 3100 -1355 3198 -1354
rect 3100 -1364 3138 -1355
rect 2688 -1407 3138 -1364
rect 3190 -1407 3198 -1355
rect 2688 -1408 3198 -1407
rect 3042 -1886 3048 -1877
rect 3027 -1929 3048 -1886
rect 3100 -1886 3106 -1877
rect 3100 -1920 3615 -1886
rect 3100 -1929 3106 -1920
rect 3027 -5538 3061 -1929
rect 3348 -1998 3400 -1992
rect 3348 -2056 3400 -2050
rect 3357 -2657 3391 -2056
rect 3581 -2270 3615 -1920
rect 3572 -2276 3624 -2270
rect 3572 -2334 3624 -2328
rect 3259 -2691 3759 -2657
rect 3259 -4057 3293 -2691
rect 3379 -2906 3431 -2900
rect 3379 -2964 3431 -2958
rect 3121 -4091 3293 -4057
rect 3121 -5123 3155 -4091
rect 3388 -4159 3422 -2964
rect 3506 -4159 3512 -4150
rect 3388 -4193 3512 -4159
rect 3506 -4202 3512 -4193
rect 3564 -4202 3570 -4150
rect 3186 -5123 3192 -5114
rect 3121 -5157 3192 -5123
rect 3186 -5166 3192 -5157
rect 3244 -5166 3250 -5114
rect 3018 -5544 3070 -5538
rect 3018 -5602 3070 -5596
use preamp  preamp_0
timestamp 1706402911
transform -1 0 4522 0 -1 -374
box 394 136 1494 1340
use th01  th01_0
timestamp 1706270854
transform 1 0 2870 0 -1 -6940
box 316 -1456 1968 6
use th10  th10_0
timestamp 1706270854
transform 1 0 3944 0 -1 -1282
box 270 -794 1168 452
use th11  th11_0
timestamp 1706241174
transform 1 0 2720 0 1 -4710
box 466 -880 1630 468
use th12  th12_0
timestamp 1706270854
transform 1 0 3422 0 1 -1986
box 278 -1078 1572 236
use th14  th14_0
timestamp 1706464016
transform 1 0 2994 0 -1 -3516
box 524 -532 1974 728
use th15  th15_0
timestamp 1706464016
transform -1 0 3478 0 -1 -1688
box 482 -1164 1936 152
<< labels >>
flabel metal1 5118 -628 5218 -528 0 FreeSans 256 180 0 0 Vn
port 17 nsew
flabel metal1 4156 -760 4256 -660 0 FreeSans 256 0 0 0 Vin
port 0 nsew
flabel metal1 4786 -1736 4886 -1636 0 FreeSans 256 0 0 0 Vp
port 1 nsew
flabel metal1 5144 -1192 5244 -1092 0 FreeSans 256 180 0 0 V10
port 10 nsew
flabel metal1 5064 -2424 5164 -2324 0 FreeSans 256 180 0 0 V12
port 12 nsew
flabel metal1 4920 -3600 5020 -3500 0 FreeSans 256 180 0 0 V14
port 14 nsew
flabel metal1 1538 -1162 1638 -1062 0 FreeSans 256 180 0 0 V15
port 15 nsew
flabel metal1 4112 -5022 4212 -4922 0 FreeSans 256 0 0 0 V11
port 11 nsew
flabel metal1 4740 -6440 4840 -6340 0 FreeSans 256 0 0 0 V01
port 2 nsew
<< end >>
