* NGSPICE file created from th08.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_JSJ4VK a_113_n42# a_n239_n216# a_n171_n42# a_n113_n130#
X0 a_113_n42# a_n113_n130# a_n171_n42# a_n239_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.13
C0 a_n171_n42# a_113_n42# 0.0218f
C1 a_n171_n42# a_n113_n130# 0.0154f
C2 a_113_n42# a_n113_n130# 0.0154f
C3 a_113_n42# a_n239_n216# 0.0734f
C4 a_n171_n42# a_n239_n216# 0.0734f
C5 a_n113_n130# a_n239_n216# 0.746f
.ends

.subckt sky130_fd_pr__pfet_01v8_EVXEQ2 a_16_n67# a_n33_n164# a_n74_n67# w_n212_n286#
+ VSUBS
X0 a_16_n67# a_n33_n164# a_n74_n67# w_n212_n286# sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.92 as=0.194 ps=1.92 w=0.67 l=0.16
C0 a_16_n67# a_n33_n164# 0.0198f
C1 a_16_n67# a_n74_n67# 0.107f
C2 a_16_n67# w_n212_n286# 0.0544f
C3 a_n74_n67# a_n33_n164# 0.0198f
C4 w_n212_n286# a_n33_n164# 0.183f
C5 a_n74_n67# w_n212_n286# 0.0184f
C6 a_16_n67# VSUBS 0.0435f
C7 a_n74_n67# VSUBS 0.0673f
C8 a_n33_n164# VSUBS 0.147f
C9 w_n212_n286# VSUBS 0.864f
.ends

.subckt sky130_fd_pr__pfet_01v8_BBE9QE w_n244_n262# a_n106_n43# a_48_n43# a_n48_n140#
+ VSUBS
X0 a_48_n43# a_n48_n140# a_n106_n43# w_n244_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.48
C0 a_n106_n43# a_48_n43# 0.041f
C1 a_n106_n43# a_n48_n140# 0.00893f
C2 a_n106_n43# w_n244_n262# 0.0225f
C3 a_n48_n140# a_48_n43# 0.00893f
C4 w_n244_n262# a_48_n43# 0.0225f
C5 a_n48_n140# w_n244_n262# 0.218f
C6 a_48_n43# VSUBS 0.0495f
C7 a_n106_n43# VSUBS 0.0495f
C8 a_n48_n140# VSUBS 0.203f
C9 w_n244_n262# VSUBS 0.876f
.ends

.subckt sky130_fd_pr__nfet_01v8_NCP4B2 a_n73_n47# a_n141_n221# a_n33_n135# a_15_n47#
X0 a_15_n47# a_n33_n135# a_n73_n47# a_n141_n221# sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.52 as=0.136 ps=1.52 w=0.47 l=0.15
C0 a_15_n47# a_n73_n47# 0.0779f
C1 a_15_n47# a_n33_n135# 0.0213f
C2 a_n73_n47# a_n33_n135# 0.0213f
C3 a_15_n47# a_n141_n221# 0.0686f
C4 a_n73_n47# a_n141_n221# 0.0686f
C5 a_n33_n135# a_n141_n221# 0.317f
.ends

.subckt th08 Vp Vin V08 Vn
XXM0 Vn Vn m1_477_n803# Vin sky130_fd_pr__nfet_01v8_JSJ4VK
XXM1 Vp Vin m1_477_n803# Vp Vn sky130_fd_pr__pfet_01v8_EVXEQ2
XXM2 Vp Vp V08 m1_477_n803# Vn sky130_fd_pr__pfet_01v8_BBE9QE
XXM3 Vn Vn m1_477_n803# V08 sky130_fd_pr__nfet_01v8_NCP4B2
C0 V08 m1_477_n803# 0.108f
C1 m1_477_n803# Vp 0.154f
C2 Vin m1_477_n803# 0.356f
C3 V08 Vp 0.0461f
C4 V08 Vin 0.00163f
C5 Vin Vp 0.0933f
C6 Vp Vn 1.66f
C7 m1_477_n803# Vn 0.656f
C8 V08 Vn 0.271f
C9 Vin Vn 1.02f
.ends

