magic
tech sky130A
magscale 1 2
timestamp 1704962149
<< nwell >>
rect -521 -261 521 261
<< pmos >>
rect -325 -42 325 42
<< pdiff >>
rect -383 30 -325 42
rect -383 -30 -371 30
rect -337 -30 -325 30
rect -383 -42 -325 -30
rect 325 30 383 42
rect 325 -30 337 30
rect 371 -30 383 30
rect 325 -42 383 -30
<< pdiffc >>
rect -371 -30 -337 30
rect 337 -30 371 30
<< nsubdiff >>
rect -485 191 -389 225
rect 389 191 485 225
rect -485 129 -451 191
rect 451 129 485 191
rect -485 -191 -451 -129
rect 451 -191 485 -129
rect -485 -225 -389 -191
rect 389 -225 485 -191
<< nsubdiffcont >>
rect -389 191 389 225
rect -485 -129 -451 129
rect 451 -129 485 129
rect -389 -225 389 -191
<< poly >>
rect -325 123 325 139
rect -325 89 -309 123
rect 309 89 325 123
rect -325 42 325 89
rect -325 -89 325 -42
rect -325 -123 -309 -89
rect 309 -123 325 -89
rect -325 -139 325 -123
<< polycont >>
rect -309 89 309 123
rect -309 -123 309 -89
<< locali >>
rect -485 191 -389 225
rect 389 191 485 225
rect -485 129 -451 191
rect 451 129 485 191
rect -325 89 -309 123
rect 309 89 325 123
rect -371 30 -337 46
rect -371 -46 -337 -30
rect 337 30 371 46
rect 337 -46 371 -30
rect -325 -123 -309 -89
rect 309 -123 325 -89
rect -485 -191 -451 -129
rect 451 -191 485 -129
rect -485 -225 -389 -191
rect 389 -225 485 -191
<< viali >>
rect -309 89 309 123
rect -371 -30 -337 30
rect 337 -30 371 30
rect -309 -123 309 -89
<< metal1 >>
rect -321 123 321 129
rect -321 89 -309 123
rect 309 89 321 123
rect -321 83 321 89
rect -377 30 -331 42
rect -377 -30 -371 30
rect -337 -30 -331 30
rect -377 -42 -331 -30
rect 331 30 377 42
rect 331 -30 337 30
rect 371 -30 377 30
rect 331 -42 377 -30
rect -321 -89 321 -83
rect -321 -123 -309 -89
rect 309 -123 321 -89
rect -321 -129 321 -123
<< properties >>
string FIXED_BBOX -468 -208 468 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 3.25 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
