magic
tech sky130A
magscale 1 2
timestamp 1706628990
<< nwell >>
rect 2878 -1714 3806 -1488
rect 3808 -1708 4222 -1544
rect 4646 -1708 4894 -1528
rect 3808 -1714 4894 -1708
rect 2878 -1754 4894 -1714
rect 2878 -1756 3866 -1754
rect 2878 -1768 3824 -1756
rect 2878 -1840 3806 -1768
rect 4214 -1796 4894 -1754
rect 4214 -1912 4890 -1796
rect 2952 -4424 3304 -4242
rect 2968 -6942 3320 -6592
rect 4637 -6862 5494 -6432
rect 6004 -6834 6106 -6410
rect 6966 -6838 7068 -6312
rect 7312 -6838 8173 -6316
rect 8276 -6824 9203 -6318
rect 8276 -6840 9554 -6824
<< pwell >>
rect 4210 -758 4260 -696
rect 2950 -5580 3358 -5546
rect 1840 -5962 2228 -5872
rect 4824 -5976 5076 -5590
rect 5320 -6092 6119 -5590
rect 6798 -6300 7564 -5796
rect 7647 -6284 8340 -5862
rect 8632 -6084 9308 -5652
<< locali >>
rect 3673 -2476 3770 -2438
<< viali >>
rect 3639 -2476 3673 -2438
rect 3554 -3395 3588 -3361
rect 4896 -4151 4930 -4117
<< metal1 >>
rect 1766 -545 4843 -511
rect 3028 -598 3072 -545
rect 5118 -559 5218 -528
rect 4957 -593 5443 -559
rect 1530 -1108 1536 -1056
rect 1588 -1062 1594 -1056
rect 1588 -1108 1638 -1062
rect 1538 -1162 1638 -1108
rect 1585 -1327 1619 -1162
rect 2945 -1842 2979 -1651
rect 3028 -1714 3065 -598
rect 5118 -628 5218 -593
rect 4156 -698 4256 -660
rect 4156 -702 4308 -698
rect 4156 -754 4209 -702
rect 4261 -754 4308 -702
rect 4156 -758 4308 -754
rect 4156 -760 4256 -758
rect 5409 -769 5443 -593
rect 5228 -894 5234 -842
rect 5286 -894 5292 -842
rect 4982 -1135 5004 -1098
rect 4943 -1169 5004 -1135
rect 5074 -1158 5138 -1098
rect 4982 -1198 5004 -1169
rect 5176 -1232 5276 -1132
rect 4054 -1270 4106 -1264
rect 4054 -1328 4106 -1322
rect 3138 -1355 3190 -1349
rect 3138 -1413 3190 -1407
rect 5340 -1354 5417 -1295
rect 5340 -1391 5420 -1354
rect 5340 -1392 5404 -1391
rect 3022 -1720 3074 -1714
rect 3022 -1778 3074 -1772
rect 1747 -2502 1781 -2325
rect 1700 -2538 1800 -2502
rect 1700 -2590 1714 -2538
rect 1766 -2590 1800 -2538
rect 1700 -2602 1800 -2590
rect 1786 -2956 1823 -2879
rect 1774 -3008 1780 -2956
rect 1832 -3008 1838 -2956
rect 2151 -3012 2203 -3006
rect 2151 -3070 2203 -3064
rect 3331 -3095 3365 -1445
rect 3581 -1591 3615 -1545
rect 4822 -1604 4834 -1598
rect 4814 -1636 4862 -1604
rect 4786 -1669 4886 -1636
rect 5340 -1669 5377 -1392
rect 4217 -1703 5377 -1669
rect 4786 -1736 4886 -1703
rect 4151 -1992 4157 -1940
rect 4209 -1992 4215 -1940
rect 3620 -2324 3626 -2272
rect 3678 -2276 3684 -2272
rect 3678 -2315 3878 -2276
rect 3678 -2324 3684 -2315
rect 5064 -2360 5164 -2324
rect 4956 -2416 5286 -2360
rect 5064 -2424 5164 -2416
rect 3538 -2438 3590 -2432
rect 3633 -2438 3679 -2426
rect 3633 -2447 3639 -2438
rect 3590 -2476 3639 -2447
rect 3673 -2476 3679 -2438
rect 3590 -2481 3679 -2476
rect 3633 -2488 3679 -2481
rect 3538 -2496 3590 -2490
rect 5230 -2772 5286 -2416
rect 5315 -3005 5407 -2971
rect 5315 -3025 5349 -3005
rect 4624 -3059 5349 -3025
rect 3614 -3072 3786 -3059
rect 3331 -3129 3601 -3095
rect 3614 -3116 3788 -3072
rect 3627 -3122 3788 -3116
rect 2145 -3304 2151 -3252
rect 2203 -3304 2209 -3252
rect 3331 -3549 3365 -3129
rect 3521 -3270 3555 -3249
rect 3486 -3322 3492 -3270
rect 3544 -3322 3555 -3270
rect 3501 -3333 3555 -3322
rect 3501 -3343 3595 -3333
rect 3501 -3361 3597 -3343
rect 3501 -3395 3554 -3361
rect 3588 -3395 3597 -3361
rect 3501 -3403 3597 -3395
rect 3548 -3407 3594 -3403
rect 3159 -3583 3365 -3549
rect 4920 -3530 5020 -3500
rect 4920 -3582 4934 -3530
rect 4986 -3582 5020 -3530
rect 2634 -3649 2734 -3600
rect 2994 -3612 3046 -3606
rect 2634 -3683 2853 -3649
rect 2994 -3670 3046 -3664
rect 2634 -3700 2734 -3683
rect 1699 -3841 1837 -3807
rect 1699 -6011 1733 -3841
rect 3159 -3955 3193 -3583
rect 4920 -3600 5020 -3582
rect 5238 -3542 5413 -3499
rect 3269 -3673 3786 -3636
rect 3269 -3739 3306 -3673
rect 4931 -3687 4965 -3600
rect 4781 -3721 4965 -3687
rect 3257 -3791 3263 -3739
rect 3315 -3791 3321 -3739
rect 3015 -3989 3193 -3955
rect 3015 -4400 3049 -3989
rect 4890 -4112 4936 -4105
rect 5238 -4112 5281 -3542
rect 4890 -4117 5281 -4112
rect 4890 -4151 4896 -4117
rect 4930 -4151 5281 -4117
rect 4890 -4155 5281 -4151
rect 4890 -4163 4936 -4155
rect 3082 -4348 3088 -4296
rect 3140 -4305 3146 -4296
rect 3140 -4339 3255 -4305
rect 3140 -4348 3146 -4339
rect 3372 -4370 3424 -4364
rect 3015 -4487 3059 -4400
rect 3372 -4428 3424 -4422
rect 5173 -4487 5207 -4311
rect 1793 -5181 1827 -5093
rect 1793 -5190 1855 -5181
rect 1793 -5215 1921 -5190
rect 1801 -5224 1921 -5215
rect 1801 -5286 1835 -5224
rect 1786 -5386 1886 -5286
rect 1805 -5911 1839 -5386
rect 2933 -5477 2939 -5425
rect 2991 -5477 2997 -5425
rect 2755 -5695 2789 -5583
rect 3025 -5695 3059 -4487
rect 4081 -4521 5207 -4487
rect 3902 -4702 3908 -4693
rect 3195 -4736 3908 -4702
rect 3902 -4745 3908 -4736
rect 3960 -4745 3966 -4693
rect 4112 -5022 4212 -4922
rect 5612 -5276 5664 -5270
rect 4877 -5319 5612 -5285
rect 3874 -5508 3911 -5490
rect 3314 -5537 3366 -5531
rect 3300 -5582 3314 -5545
rect 3863 -5545 3911 -5508
rect 3366 -5582 3954 -5545
rect 3824 -5586 3911 -5582
rect 3314 -5595 3366 -5589
rect 2755 -5729 3059 -5695
rect 2253 -5850 2259 -5798
rect 2311 -5850 2317 -5798
rect 3025 -5817 3059 -5729
rect 3543 -5799 3595 -5793
rect 3025 -5851 3283 -5817
rect 3431 -5842 3543 -5808
rect 3431 -5911 3465 -5842
rect 3543 -5857 3595 -5851
rect 1805 -5945 3465 -5911
rect 1699 -6045 1925 -6011
rect 4877 -6037 4911 -5319
rect 5612 -5334 5664 -5328
rect 5078 -5760 5084 -5708
rect 5136 -5760 5142 -5708
rect 9703 -5751 9737 -5177
rect 5968 -5782 6020 -5776
rect 5916 -5834 5968 -5802
rect 5916 -5840 6020 -5834
rect 5916 -5902 6016 -5840
rect 6198 -5883 6204 -5836
rect 6173 -5888 6204 -5883
rect 6256 -5883 6262 -5836
rect 6256 -5888 6277 -5883
rect 6173 -5917 6277 -5888
rect 7081 -5935 7087 -5883
rect 7139 -5935 7145 -5883
rect 4807 -6071 4911 -6037
rect 6936 -6068 6942 -6016
rect 6994 -6068 7000 -6016
rect 7971 -6075 7977 -6023
rect 8029 -6042 8035 -6023
rect 8029 -6075 8054 -6042
rect 7994 -6076 8054 -6075
rect 8857 -6121 8863 -6069
rect 8915 -6121 8921 -6069
rect 6882 -6244 6982 -6144
rect 8746 -6186 8752 -6178
rect 8698 -6230 8752 -6186
rect 8804 -6230 8810 -6178
rect 8698 -6286 8798 -6230
rect 7761 -6307 7813 -6301
rect 3080 -6454 3086 -6402
rect 3141 -6454 3147 -6402
rect 4740 -6440 4840 -6340
rect 7761 -6365 7813 -6359
rect 9954 -6316 10006 -6310
rect 9954 -6378 10006 -6372
rect 3080 -6455 3209 -6454
rect 3080 -6456 3232 -6455
rect 3080 -6464 3401 -6456
rect 3079 -6498 3401 -6464
rect 3202 -6499 3401 -6498
rect 7732 -6572 7832 -6472
rect 9914 -6610 10014 -6510
rect 6072 -6620 6124 -6614
rect 6072 -6678 6124 -6672
rect 2386 -6980 2486 -6958
rect 2386 -7032 2438 -6980
rect 2490 -7032 2496 -6980
rect 2386 -7060 2486 -7032
<< via1 >>
rect 1536 -1108 1588 -1056
rect 4209 -754 4261 -702
rect 5234 -894 5286 -842
rect 4054 -1322 4106 -1270
rect 3138 -1407 3190 -1355
rect 3022 -1772 3074 -1720
rect 1714 -2590 1766 -2538
rect 1780 -3008 1832 -2956
rect 2151 -3064 2203 -3012
rect 4157 -1992 4209 -1940
rect 3626 -2324 3678 -2272
rect 3538 -2490 3590 -2438
rect 2151 -3304 2203 -3252
rect 3492 -3322 3544 -3270
rect 4934 -3582 4986 -3530
rect 2994 -3664 3046 -3612
rect 3263 -3791 3315 -3739
rect 3088 -4348 3140 -4296
rect 3372 -4422 3424 -4370
rect 2939 -5477 2991 -5425
rect 3908 -4745 3960 -4693
rect 3314 -5589 3366 -5537
rect 2259 -5850 2311 -5798
rect 3543 -5851 3595 -5799
rect 5612 -5328 5664 -5276
rect 5084 -5760 5136 -5708
rect 5968 -5834 6020 -5782
rect 6204 -5888 6256 -5836
rect 7087 -5935 7139 -5883
rect 6942 -6068 6994 -6016
rect 7977 -6075 8029 -6023
rect 8863 -6121 8915 -6069
rect 8752 -6230 8804 -6178
rect 3086 -6454 3141 -6402
rect 7761 -6359 7813 -6307
rect 9954 -6372 10006 -6316
rect 6072 -6672 6124 -6620
rect 2438 -7032 2490 -6980
<< metal2 >>
rect 1452 -376 6610 -332
rect 1452 -2542 1496 -376
rect 1538 -460 5284 -412
rect 1538 -1050 1586 -460
rect 4209 -702 4261 -696
rect 4209 -760 4218 -754
rect 4252 -760 4261 -754
rect 5236 -836 5284 -460
rect 5795 -606 5804 -550
rect 5860 -606 5869 -550
rect 6566 -622 6610 -376
rect 6566 -666 7596 -622
rect 6566 -670 6610 -666
rect 5234 -842 5286 -836
rect 5234 -900 5286 -894
rect 1536 -1056 1588 -1050
rect 1536 -1114 1588 -1108
rect 4048 -1322 4054 -1270
rect 4106 -1279 4112 -1270
rect 4106 -1313 4252 -1279
rect 4106 -1322 4112 -1313
rect 3100 -1355 3198 -1354
rect 3100 -1364 3138 -1355
rect 2688 -1407 3138 -1364
rect 3190 -1407 3198 -1355
rect 2688 -1408 3198 -1407
rect 3016 -1772 3022 -1720
rect 3074 -1729 3080 -1720
rect 3074 -1763 3669 -1729
rect 3074 -1772 3080 -1763
rect 3635 -2266 3669 -1763
rect 4055 -1743 4089 -1322
rect 4055 -1777 4200 -1743
rect 4166 -1934 4200 -1777
rect 5124 -1778 5180 -1769
rect 5124 -1843 5180 -1834
rect 4157 -1940 4209 -1934
rect 4157 -1998 4209 -1992
rect 3626 -2272 3678 -2266
rect 3626 -2330 3678 -2324
rect 3626 -2331 3663 -2330
rect 3481 -2492 3490 -2436
rect 3546 -2438 3555 -2436
rect 3590 -2490 3596 -2438
rect 3546 -2492 3555 -2490
rect 1708 -2542 1714 -2538
rect 1452 -2586 1714 -2542
rect 1708 -2590 1714 -2586
rect 1766 -2590 1772 -2538
rect 1780 -2956 1832 -2950
rect 1780 -3014 1832 -3008
rect 3405 -2961 3766 -2927
rect 1783 -3043 1828 -3014
rect 1768 -3099 1777 -3043
rect 1833 -3099 1842 -3043
rect 2145 -3064 2151 -3012
rect 2203 -3064 2209 -3012
rect 3405 -3023 3439 -2961
rect 2795 -3057 3439 -3023
rect 2160 -3246 2194 -3064
rect 2151 -3252 2203 -3246
rect 2151 -3310 2203 -3304
rect 3030 -3610 3086 -3601
rect 2988 -3664 2994 -3612
rect 3030 -3675 3086 -3666
rect 3263 -3739 3315 -3733
rect 3263 -3797 3315 -3791
rect 3266 -3826 3311 -3797
rect 3251 -3882 3260 -3826
rect 3316 -3882 3325 -3826
rect 3088 -4296 3140 -4290
rect 3077 -4376 3086 -4320
rect 3142 -4376 3151 -4320
rect 3405 -4370 3439 -3057
rect 5258 -3146 5314 -3137
rect 4943 -3191 5258 -3157
rect 3481 -3288 3490 -3232
rect 3546 -3288 3555 -3232
rect 3492 -3328 3544 -3322
rect 4943 -3524 4977 -3191
rect 5258 -3211 5314 -3202
rect 4934 -3530 4986 -3524
rect 4934 -3588 4986 -3582
rect 3366 -4422 3372 -4370
rect 3424 -4413 3439 -4370
rect 3424 -4422 3430 -4413
rect 3908 -4693 3960 -4687
rect 3960 -4736 4255 -4702
rect 3908 -4751 3960 -4745
rect 4221 -4849 4255 -4736
rect 4221 -4883 5123 -4849
rect 5089 -5071 5123 -4883
rect 5089 -5096 5127 -5071
rect 5073 -5152 5082 -5096
rect 5138 -5152 5147 -5096
rect 5606 -5328 5612 -5276
rect 5664 -5288 5670 -5276
rect 5715 -5288 5743 -5224
rect 5664 -5316 5743 -5288
rect 5664 -5328 5670 -5316
rect 5855 -5331 6068 -5288
rect 2929 -5390 2938 -5334
rect 2994 -5390 3003 -5334
rect 5855 -5384 5898 -5331
rect 6466 -5338 6676 -5294
rect 7131 -5311 7419 -5269
rect 9049 -5287 9403 -5245
rect 6466 -5384 6510 -5338
rect 2943 -5419 2988 -5390
rect 4367 -5396 5520 -5384
rect 5854 -5396 5898 -5384
rect 2939 -5425 2991 -5419
rect 2939 -5483 2991 -5477
rect 4367 -5427 5898 -5396
rect 2941 -5538 2984 -5483
rect 3308 -5538 3314 -5537
rect 2941 -5581 3314 -5538
rect 2259 -5798 2311 -5792
rect 2941 -5836 2984 -5581
rect 3308 -5589 3314 -5581
rect 3366 -5589 3372 -5537
rect 2311 -5850 2984 -5836
rect 2259 -5856 2984 -5850
rect 3537 -5851 3543 -5799
rect 3595 -5804 3601 -5799
rect 4367 -5804 4410 -5427
rect 5435 -5439 5898 -5427
rect 6008 -5428 6510 -5384
rect 7131 -5401 7173 -5311
rect 7776 -5336 7954 -5292
rect 7776 -5374 7820 -5336
rect 6008 -5488 6052 -5428
rect 6595 -5443 7173 -5401
rect 7248 -5418 7820 -5374
rect 8577 -5349 8814 -5306
rect 8577 -5376 8620 -5349
rect 6595 -5473 6637 -5443
rect 3595 -5847 4410 -5804
rect 4970 -5532 6052 -5488
rect 6133 -5515 6637 -5473
rect 7248 -5484 7292 -5418
rect 3595 -5851 3601 -5847
rect 2263 -5879 2984 -5856
rect 3076 -6411 3085 -6355
rect 3141 -6411 3150 -6355
rect 3086 -6460 3141 -6454
rect 2438 -6980 2490 -6974
rect 4970 -6984 5014 -5532
rect 6133 -5645 6175 -5515
rect 5073 -5714 5082 -5658
rect 5138 -5714 5147 -5658
rect 5973 -5687 6175 -5645
rect 6946 -5528 7292 -5484
rect 7897 -5419 8620 -5376
rect 9049 -5409 9091 -5287
rect 7897 -5500 7940 -5419
rect 5084 -5766 5136 -5760
rect 5973 -5782 6015 -5687
rect 5962 -5834 5968 -5782
rect 6020 -5834 6026 -5782
rect 6193 -5862 6202 -5806
rect 6258 -5862 6267 -5806
rect 6204 -5894 6256 -5888
rect 6946 -6010 6990 -5528
rect 7829 -5543 7940 -5500
rect 8757 -5451 9091 -5409
rect 7075 -5904 7084 -5848
rect 7140 -5904 7149 -5848
rect 7087 -5941 7139 -5935
rect 6942 -6016 6994 -6010
rect 6942 -6074 6994 -6068
rect 7829 -6304 7872 -5543
rect 7965 -6036 7974 -5980
rect 8030 -6036 8039 -5980
rect 7977 -6081 8029 -6075
rect 8757 -6172 8799 -5451
rect 8851 -6080 8860 -6024
rect 8916 -6080 8925 -6024
rect 8863 -6127 8915 -6121
rect 8752 -6178 8804 -6172
rect 8752 -6236 8804 -6230
rect 7783 -6307 7872 -6304
rect 7755 -6359 7761 -6307
rect 7813 -6355 7872 -6307
rect 10080 -6316 10136 -5238
rect 7813 -6359 7819 -6355
rect 9948 -6372 9954 -6316
rect 10006 -6372 10136 -6316
rect 5448 -6618 5504 -6609
rect 5448 -6683 5504 -6674
rect 6038 -6618 6094 -6609
rect 6124 -6672 6130 -6620
rect 6038 -6683 6094 -6674
rect 2490 -7028 5014 -6984
rect 2438 -7038 2490 -7032
<< via2 >>
rect 5804 -606 5860 -550
rect 5124 -1834 5180 -1778
rect 3490 -2438 3546 -2436
rect 3490 -2490 3538 -2438
rect 3538 -2490 3546 -2438
rect 3490 -2492 3546 -2490
rect 1777 -3099 1833 -3043
rect 3030 -3612 3086 -3610
rect 3030 -3664 3046 -3612
rect 3046 -3664 3086 -3612
rect 3030 -3666 3086 -3664
rect 3260 -3882 3316 -3826
rect 3086 -4348 3088 -4320
rect 3088 -4348 3140 -4320
rect 3140 -4348 3142 -4320
rect 3086 -4376 3142 -4348
rect 3490 -3270 3546 -3232
rect 3490 -3288 3492 -3270
rect 3492 -3288 3544 -3270
rect 3544 -3288 3546 -3270
rect 5258 -3202 5314 -3146
rect 5082 -5152 5138 -5096
rect 2938 -5390 2994 -5334
rect 3085 -6402 3141 -6355
rect 3085 -6411 3086 -6402
rect 3086 -6411 3141 -6402
rect 5082 -5708 5138 -5658
rect 5082 -5714 5084 -5708
rect 5084 -5714 5136 -5708
rect 5136 -5714 5138 -5708
rect 6202 -5836 6258 -5806
rect 6202 -5862 6204 -5836
rect 6204 -5862 6256 -5836
rect 6256 -5862 6258 -5836
rect 7084 -5883 7140 -5848
rect 7084 -5904 7087 -5883
rect 7087 -5904 7139 -5883
rect 7139 -5904 7140 -5883
rect 7974 -6023 8030 -5980
rect 7974 -6036 7977 -6023
rect 7977 -6036 8029 -6023
rect 8029 -6036 8030 -6023
rect 8860 -6069 8916 -6024
rect 8860 -6080 8863 -6069
rect 8863 -6080 8915 -6069
rect 8915 -6080 8916 -6069
rect 5448 -6674 5504 -6618
rect 6038 -6620 6094 -6618
rect 6038 -6672 6072 -6620
rect 6072 -6672 6094 -6620
rect 6038 -6674 6094 -6672
<< metal3 >>
rect 5684 -266 5985 -146
rect 5802 -545 5862 -266
rect 5799 -550 5865 -545
rect 5799 -606 5804 -550
rect 5860 -606 5865 -550
rect 5799 -611 5865 -606
rect 5802 -614 5862 -611
rect 5119 -1776 5185 -1773
rect 3406 -1778 5185 -1776
rect 3406 -1834 5124 -1778
rect 5180 -1834 5185 -1778
rect 3406 -1836 5185 -1834
rect 3406 -2300 3466 -1836
rect 5119 -1839 5185 -1836
rect 10458 -1938 10578 -1756
rect 10444 -2058 10645 -1938
rect 3216 -2360 3466 -2300
rect 1767 -3017 1773 -2953
rect 1837 -3017 1843 -2953
rect 1769 -3043 1839 -3017
rect 1769 -3077 1777 -3043
rect 1772 -3099 1777 -3077
rect 1833 -3081 1839 -3043
rect 1833 -3099 1838 -3081
rect 1772 -3104 1838 -3099
rect 3216 -3376 3276 -2360
rect 3485 -2436 3551 -2431
rect 3485 -2492 3490 -2436
rect 3546 -2492 3551 -2436
rect 3485 -2497 3551 -2492
rect 3488 -3227 3548 -2497
rect 10848 -2630 10968 -2470
rect 10812 -2750 11013 -2630
rect 5253 -3144 5319 -3141
rect 5253 -3146 5396 -3144
rect 5253 -3202 5258 -3146
rect 5314 -3202 5396 -3146
rect 5253 -3204 5396 -3202
rect 5253 -3207 5319 -3204
rect 3485 -3232 3551 -3227
rect 3485 -3288 3490 -3232
rect 3546 -3288 3551 -3232
rect 3485 -3293 3551 -3288
rect 3028 -3436 3276 -3376
rect 3028 -3605 3088 -3436
rect 3025 -3610 3091 -3605
rect 3025 -3666 3030 -3610
rect 3086 -3666 3091 -3610
rect 3025 -3671 3091 -3666
rect 3250 -3800 3256 -3736
rect 3320 -3800 3326 -3736
rect 3252 -3826 3322 -3800
rect 3252 -3860 3260 -3826
rect 3255 -3882 3260 -3860
rect 3316 -3864 3322 -3826
rect 3316 -3882 3321 -3864
rect 3255 -3887 3321 -3882
rect 10608 -4250 10909 -4130
rect 3081 -4320 3147 -4315
rect 3081 -4376 3086 -4320
rect 3142 -4376 3147 -4320
rect 3081 -4381 3147 -4376
rect 2933 -5334 2999 -5329
rect 2933 -5352 2938 -5334
rect 2932 -5390 2938 -5352
rect 2994 -5356 2999 -5334
rect 2994 -5390 3002 -5356
rect 2932 -5416 3002 -5390
rect 2928 -5480 2934 -5416
rect 2998 -5480 3004 -5416
rect 3084 -6253 3144 -4381
rect 10674 -4444 10794 -4250
rect 5077 -5096 5143 -5091
rect 5077 -5152 5082 -5096
rect 5138 -5152 5143 -5096
rect 5077 -5157 5143 -5152
rect 5080 -5653 5140 -5157
rect 5077 -5658 5143 -5653
rect 5077 -5714 5082 -5658
rect 5138 -5714 5143 -5658
rect 5077 -5719 5143 -5714
rect 6200 -5736 8918 -5676
rect 6200 -5801 6260 -5736
rect 6197 -5806 6263 -5801
rect 6197 -5862 6202 -5806
rect 6258 -5862 6263 -5806
rect 7082 -5843 7142 -5736
rect 6197 -5867 6263 -5862
rect 7079 -5848 7145 -5843
rect 7079 -5904 7084 -5848
rect 7140 -5904 7145 -5848
rect 7079 -5909 7145 -5904
rect 7972 -5975 8032 -5736
rect 7969 -5980 8035 -5975
rect 7969 -6036 7974 -5980
rect 8030 -6036 8035 -5980
rect 8858 -6019 8918 -5736
rect 7969 -6041 8035 -6036
rect 8855 -6024 8921 -6019
rect 8855 -6080 8860 -6024
rect 8916 -6080 8921 -6024
rect 8855 -6085 8921 -6080
rect 3083 -6350 3144 -6253
rect 3080 -6355 3146 -6350
rect 3080 -6411 3085 -6355
rect 3141 -6411 3146 -6355
rect 3080 -6416 3146 -6411
rect 5443 -6616 5509 -6613
rect 6033 -6616 6099 -6613
rect 5443 -6618 6099 -6616
rect 5443 -6674 5448 -6618
rect 5504 -6674 6038 -6618
rect 6094 -6674 6099 -6618
rect 5443 -6676 6099 -6674
rect 5443 -6679 5509 -6676
rect 6033 -6679 6099 -6676
<< via3 >>
rect 1773 -3017 1837 -2953
rect 3256 -3800 3320 -3736
rect 2934 -5480 2998 -5416
<< metal4 >>
rect 1775 -2952 1835 -2913
rect 1772 -2953 1838 -2952
rect 1772 -3017 1773 -2953
rect 1837 -3017 1838 -2953
rect 1772 -3018 1838 -3017
rect 1775 -3100 1835 -3018
rect 1774 -3160 3318 -3100
rect 3258 -3735 3318 -3160
rect 3255 -3736 3321 -3735
rect 3255 -3800 3256 -3736
rect 3320 -3800 3321 -3736
rect 3255 -3801 3321 -3800
rect 3258 -4106 3318 -3801
rect 2936 -4166 3318 -4106
rect 2936 -5415 2996 -4166
rect 2933 -5416 2999 -5415
rect 2933 -5480 2934 -5416
rect 2998 -5480 2999 -5416
rect 2933 -5481 2999 -5480
rect 2936 -5484 2996 -5481
use preamp  preamp_0
timestamp 1706402911
transform -1 0 4522 0 -1 -374
box 394 136 1494 1340
use th01  th01_0
timestamp 1706270854
transform 1 0 2870 0 -1 -6940
box 316 -1456 1968 6
use th02  th02_0
timestamp 1706480381
transform -1 0 3306 0 1 -4832
box 378 -1044 1520 426
use th03  th03_0
timestamp 1706270854
transform 0 1 2811 -1 0 -5432
box 516 -1083 1680 238
use th04  th04_0
timestamp 1706270854
transform 1 0 4684 0 -1 -6714
box 374 -1126 1336 148
use th05  th05_0
timestamp 1706270876
transform 1 0 8398 0 -1 -6694
box 474 -1043 1620 148
use th06  th06_0
timestamp 1706231216
transform 1 0 7718 0 -1 -6838
box 200 -976 1084 2
use th07  th07_0
timestamp 1706236611
transform 1 0 6746 0 -1 -6808
box 314 -1014 1088 32
use th08  th08_0
timestamp 1706233216
transform 1 0 5728 0 -1 -6836
box 356 -1052 1272 -2
use th09  th09_0
timestamp 1706479318
transform 1 0 1406 0 -1 -3900
box 368 -754 1692 524
use th10  th10_0
timestamp 1706270854
transform 1 0 3944 0 -1 -1282
box 270 -794 1168 452
use th11  th11_0
timestamp 1706241174
transform 1 0 2720 0 1 -4710
box 466 -880 1630 468
use th12  th12_0
timestamp 1706270854
transform 1 0 3422 0 1 -1986
box 278 -1078 1572 236
use th13  th13_0
timestamp 1706474503
transform -1 0 3736 0 1 -2482
box 438 -680 2042 646
use th14  th14_0
timestamp 1706473616
transform 1 0 2994 0 -1 -3516
box 524 -532 1974 728
use th15  th15_0
timestamp 1706464016
transform -1 0 3478 0 -1 -1688
box 482 -1164 1936 152
use therm  therm_0
timestamp 1706575407
transform 1 0 4303 0 1 -7322
box 771 1832 7058 6890
<< labels >>
flabel metal3 s 10444 -2058 10644 -1938 0 FreeSans 480 0 0 0 b[0]
port 21 nsew signal tristate
flabel metal1 5118 -628 5218 -528 0 FreeSans 256 180 0 0 Vn
port 17 nsew
flabel metal1 9914 -6610 10014 -6510 0 FreeSans 256 0 0 0 V05
port 16 nsew
flabel metal1 8698 -6286 8798 -6186 0 FreeSans 256 0 0 0 V06
port 8 nsew
flabel metal1 7732 -6572 7832 -6472 0 FreeSans 256 0 0 0 V07
port 7 nsew
flabel metal1 6882 -6244 6982 -6144 0 FreeSans 256 0 0 0 V08
port 6 nsew
flabel metal1 5916 -5902 6016 -5802 0 FreeSans 256 0 0 0 V04
port 5 nsew
flabel metal1 2386 -7060 2486 -6960 0 FreeSans 256 90 0 0 V03
port 4 nsew
flabel metal1 1786 -5386 1886 -5286 0 FreeSans 256 180 0 0 V02
port 3 nsew
flabel metal1 2634 -3700 2734 -3600 0 FreeSans 256 0 0 0 V09
port 9 nsew
flabel metal1 1700 -2602 1800 -2502 0 FreeSans 256 180 0 0 V13
port 13 nsew
flabel metal1 4740 -6440 4840 -6340 0 FreeSans 256 0 0 0 V01
port 2 nsew
flabel metal1 4112 -5022 4212 -4922 0 FreeSans 256 0 0 0 V11
port 11 nsew
flabel metal1 1538 -1162 1638 -1062 0 FreeSans 256 180 0 0 V15
port 15 nsew
flabel metal1 4920 -3600 5020 -3500 0 FreeSans 256 180 0 0 V14
port 14 nsew
flabel metal1 5064 -2424 5164 -2324 0 FreeSans 256 180 0 0 V12
port 12 nsew
flabel metal1 4786 -1736 4886 -1636 0 FreeSans 256 0 0 0 Vp
port 1 nsew
flabel metal1 4156 -760 4256 -660 0 FreeSans 256 0 0 0 Vin
port 0 nsew
flabel metal3 s 5684 -266 5984 -146 0 FreeSans 480 0 0 0 b[3]
port 20 nsew signal tristate
flabel metal3 s 10608 -4250 10908 -4130 0 FreeSans 480 0 0 0 b[1]
port 18 nsew signal tristate
rlabel metal3 10905 -4196 10905 -4196 0 b[1]
flabel metal3 s 10812 -2750 11012 -2630 0 FreeSans 480 0 0 0 b[2]
port 19 nsew signal tristate
flabel metal1 5176 -1232 5276 -1132 0 FreeSans 256 0 0 0 V10
port 10 nsew
<< end >>
