/home/cae3/Desktop/ADC/ASIC_ADC/PNR/lef/sky130_scl_9T.lef