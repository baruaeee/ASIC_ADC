* NGSPICE file created from therm_port_resized.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X a_208_47# a_75_199#
+ a_544_297# a_315_47# a_201_297#
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_201_297# A1 0.011f
C1 a_208_47# X 1.91e-19
C2 A2 a_208_47# 0.00102f
C3 A3 VGND 0.0161f
C4 a_75_199# B1 0.102f
C5 a_208_47# VPWR 8.35e-19
C6 a_544_297# X 2.35e-19
C7 a_544_297# VPWR 0.0105f
C8 a_201_297# B1 0.00594f
C9 A1 B1 0.0716f
C10 a_75_199# A3 0.163f
C11 A2 a_315_47# 0.00335f
C12 a_208_47# VGND 0.00302f
C13 a_315_47# VPWR 0.00154f
C14 X VPB 0.0107f
C15 A2 VPB 0.0376f
C16 VPB VPWR 0.0749f
C17 a_544_297# VGND 0.00256f
C18 a_201_297# A3 0.00642f
C19 a_208_47# a_75_199# 0.0159f
C20 C1 X 5.14e-20
C21 a_315_47# VGND 0.00427f
C22 C1 VPWR 0.0146f
C23 VPB VGND 0.00772f
C24 a_75_199# a_544_297# 0.0176f
C25 a_75_199# a_315_47# 0.0202f
C26 C1 VGND 0.0181f
C27 a_544_297# a_201_297# 0.00702f
C28 a_75_199# VPB 0.0486f
C29 A1 a_315_47# 0.00313f
C30 A2 X 3.01e-19
C31 a_201_297# VPB 0.00186f
C32 A1 VPB 0.0306f
C33 a_75_199# C1 0.0628f
C34 a_544_297# B1 1.13e-19
C35 X VPWR 0.0676f
C36 A2 VPWR 0.0174f
C37 a_208_47# A3 3.65e-19
C38 a_201_297# C1 0.00243f
C39 A1 C1 3.21e-19
C40 B1 VPB 0.0292f
C41 X VGND 0.0609f
C42 A2 VGND 0.0119f
C43 VPWR VGND 0.0735f
C44 B1 C1 0.066f
C45 A3 VPB 0.0268f
C46 a_75_199# X 0.0959f
C47 A2 a_75_199# 0.0621f
C48 a_75_199# VPWR 0.109f
C49 a_201_297# X 0.0131f
C50 A2 a_201_297# 0.0112f
C51 A1 X 1.2e-19
C52 A2 A1 0.0689f
C53 a_201_297# VPWR 0.211f
C54 A1 VPWR 0.0151f
C55 a_75_199# VGND 0.362f
C56 B1 X 7.79e-20
C57 a_201_297# VGND 0.00403f
C58 A1 VGND 0.0113f
C59 B1 VPWR 0.0125f
C60 A3 X 0.00317f
C61 A2 A3 0.0747f
C62 A3 VPWR 0.0181f
C63 B1 VGND 0.0171f
C64 a_75_199# a_201_297# 0.16f
C65 a_75_199# A1 0.0696f
C66 C1 VPB 0.0394f
C67 VGND VNB 0.437f
C68 VPWR VNB 0.365f
C69 X VNB 0.0906f
C70 C1 VNB 0.148f
C71 B1 VNB 0.0947f
C72 A1 VNB 0.101f
C73 A2 VNB 0.11f
C74 A3 VNB 0.0908f
C75 VPB VNB 0.782f
C76 a_201_297# VNB 0.00345f
C77 a_75_199# VNB 0.205f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_181_47# a_109_47# a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_27_47# VPWR 0.145f
C1 VGND VPB 0.00604f
C2 a_109_47# VGND 0.00123f
C3 VGND B 0.00714f
C4 C a_27_47# 0.186f
C5 VPB A 0.0426f
C6 a_109_47# A 6.45e-19
C7 A B 0.0869f
C8 VGND VPWR 0.0475f
C9 X a_27_47# 0.087f
C10 a_181_47# a_27_47# 0.00401f
C11 A VPWR 0.0185f
C12 C VGND 0.0703f
C13 VGND X 0.0708f
C14 VGND a_181_47# 0.00261f
C15 VPB B 0.0836f
C16 VGND a_27_47# 0.134f
C17 VPB VPWR 0.0795f
C18 a_109_47# VPWR 3.29e-19
C19 B VPWR 0.128f
C20 a_27_47# A 0.157f
C21 C VPB 0.0347f
C22 C B 0.0746f
C23 X VPB 0.0121f
C24 X B 0.00111f
C25 C VPWR 0.00464f
C26 VGND A 0.0154f
C27 X VPWR 0.0766f
C28 a_181_47# VPWR 3.97e-19
C29 a_27_47# VPB 0.0501f
C30 a_109_47# a_27_47# 0.00517f
C31 a_27_47# B 0.0625f
C32 C X 0.0149f
C33 C a_181_47# 0.00151f
C34 VGND VNB 0.3f
C35 X VNB 0.0923f
C36 C VNB 0.12f
C37 A VNB 0.174f
C38 VPWR VNB 0.274f
C39 B VNB 0.102f
C40 VPB VNB 0.516f
C41 a_27_47# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
C0 VGND VPB 0.0797f
C1 VPWR VPB 0.0625f
C2 VGND VPWR 0.353f
C3 VPWR VNB 0.47f
C4 VGND VNB 0.427f
C5 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VGND VPB 0.116f
C1 VPWR VPB 0.0787f
C2 VGND VPWR 0.546f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_384_47# a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
C0 A1 a_384_47# 0.00884f
C1 VGND a_81_21# 0.173f
C2 X VPB 0.0108f
C3 VPB VPWR 0.068f
C4 VPB A2 0.0373f
C5 X B1 3.04e-20
C6 a_384_47# VGND 0.00366f
C7 B1 VPWR 0.0196f
C8 a_299_297# VPWR 0.202f
C9 a_299_297# A2 0.0468f
C10 VPB a_81_21# 0.0593f
C11 B1 a_81_21# 0.148f
C12 A1 VGND 0.0786f
C13 a_299_297# a_81_21# 0.0821f
C14 a_384_47# a_299_297# 1.48e-19
C15 A1 VPB 0.0264f
C16 X VPWR 0.0847f
C17 A1 B1 0.0817f
C18 VPWR A2 0.0201f
C19 A1 a_299_297# 0.0585f
C20 VPB VGND 0.00713f
C21 X a_81_21# 0.112f
C22 VPWR a_81_21# 0.146f
C23 A2 a_81_21# 7.47e-19
C24 VGND B1 0.0181f
C25 VGND a_299_297# 0.00772f
C26 a_384_47# VPWR 4.08e-19
C27 VPB B1 0.0387f
C28 a_384_47# a_81_21# 0.00138f
C29 VPB a_299_297# 0.0111f
C30 A1 VPWR 0.0209f
C31 A1 A2 0.0921f
C32 B1 a_299_297# 0.00863f
C33 A1 a_81_21# 0.0568f
C34 X VGND 0.0512f
C35 VGND VPWR 0.0579f
C36 VGND A2 0.0495f
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 Y VPB 0.0061f
C1 VPB VGND 0.00649f
C2 VPB VPWR 0.0521f
C3 Y VGND 0.155f
C4 Y VPWR 0.209f
C5 A VPB 0.0742f
C6 VGND VPWR 0.0423f
C7 Y A 0.0894f
C8 A VGND 0.0638f
C9 A VPWR 0.0631f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X a_29_53# a_183_297# a_111_297#
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 VPB a_29_53# 0.0491f
C1 a_29_53# VPWR 0.0833f
C2 X B 6.52e-19
C3 a_111_297# VPWR 5.94e-19
C4 VPB A 0.0377f
C5 A VPWR 0.00936f
C6 C B 0.0802f
C7 VPB VGND 0.00724f
C8 VPWR VGND 0.0459f
C9 X a_29_53# 0.0991f
C10 a_29_53# C 0.0857f
C11 X A 0.00127f
C12 a_183_297# a_29_53# 0.00868f
C13 X VGND 0.036f
C14 C A 0.0343f
C15 VPB VPWR 0.0649f
C16 a_183_297# A 0.00239f
C17 C VGND 0.0161f
C18 a_29_53# B 0.121f
C19 a_183_297# VGND 5.75e-19
C20 B A 0.0787f
C21 VPB X 0.0109f
C22 X VPWR 0.0885f
C23 B VGND 0.0152f
C24 VPB C 0.0396f
C25 C VPWR 0.00457f
C26 a_29_53# a_111_297# 0.005f
C27 a_29_53# A 0.242f
C28 a_183_297# VPWR 8.13e-19
C29 a_111_297# A 0.00223f
C30 a_29_53# VGND 0.217f
C31 a_111_297# VGND 3.96e-19
C32 VPB B 0.0962f
C33 B VPWR 0.147f
C34 A VGND 0.0187f
C35 VGND VNB 0.306f
C36 X VNB 0.0882f
C37 A VNB 0.117f
C38 C VNB 0.16f
C39 B VNB 0.117f
C40 VPWR VNB 0.253f
C41 VPB VNB 0.516f
C42 a_29_53# VNB 0.18f
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 Y VPB 0.0139f
C1 A VGND 0.0486f
C2 B VPB 0.0367f
C3 a_109_297# VPWR 0.00638f
C4 VGND VPWR 0.0314f
C5 Y A 0.0471f
C6 Y VPWR 0.0995f
C7 B A 0.0584f
C8 a_109_297# VGND 0.00128f
C9 B VPWR 0.0148f
C10 VPB A 0.0415f
C11 a_109_297# Y 0.0113f
C12 Y VGND 0.154f
C13 VPB VPWR 0.0449f
C14 B VGND 0.0451f
C15 Y B 0.0877f
C16 VPB VGND 0.00456f
C17 A VPWR 0.0528f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
C0 VPWR VGND 0.903f
C1 VPB VGND 0.161f
C2 VPB VPWR 0.0858f
C3 VPWR VNB 0.867f
C4 VGND VNB 0.761f
C5 VPB VNB 0.605f
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X a_193_297# a_465_47#
+ a_205_47# a_109_297# a_27_47#
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
C0 VPB a_109_297# 0.00421f
C1 X B2 6.77e-20
C2 X B1 9.58e-20
C3 VPB C1 0.0367f
C4 VPWR a_109_297# 0.15f
C5 a_109_297# A1 1.05e-19
C6 VGND B2 0.0174f
C7 B2 a_27_47# 0.0959f
C8 VGND B1 0.0133f
C9 VGND a_205_47# 0.00156f
C10 a_27_47# B1 0.112f
C11 a_27_47# a_205_47# 0.00762f
C12 VPWR C1 0.0139f
C13 C1 A1 1.77e-20
C14 B2 a_193_297# 0.00126f
C15 B1 a_193_297# 0.00869f
C16 VPWR VPB 0.0799f
C17 X a_109_297# 3.99e-19
C18 VPB A1 0.0343f
C19 X C1 5.03e-20
C20 VGND a_109_297# 0.00284f
C21 a_109_297# a_27_47# 0.0961f
C22 VPWR A1 0.0161f
C23 X VPB 0.0113f
C24 VGND C1 0.0196f
C25 A2 C1 9.03e-21
C26 a_109_297# a_193_297# 0.0927f
C27 C1 a_27_47# 0.0792f
C28 B2 B1 0.0784f
C29 VGND VPB 0.00844f
C30 A2 VPB 0.027f
C31 X VPWR 0.0897f
C32 VPB a_27_47# 0.0512f
C33 X A1 2.77e-19
C34 VPWR a_465_47# 5.05e-19
C35 a_465_47# A1 7.06e-19
C36 VPB a_193_297# 0.00774f
C37 VGND VPWR 0.0722f
C38 A2 VPWR 0.0209f
C39 VGND A1 0.0126f
C40 A2 A1 0.0692f
C41 VPWR a_27_47# 0.099f
C42 A1 a_27_47# 0.0984f
C43 B2 a_109_297# 0.0133f
C44 a_109_297# B1 0.00736f
C45 X a_465_47# 1.56e-19
C46 VPWR a_193_297# 0.169f
C47 A1 a_193_297# 0.0109f
C48 B2 C1 0.0726f
C49 X VGND 0.061f
C50 X A2 0.00157f
C51 C1 B1 6.46e-19
C52 X a_27_47# 0.0921f
C53 VGND a_465_47# 0.00257f
C54 a_465_47# a_27_47# 0.013f
C55 B2 VPB 0.0256f
C56 VPB B1 0.0321f
C57 X a_193_297# 0.00367f
C58 VGND A2 0.0168f
C59 VGND a_27_47# 0.395f
C60 A2 a_27_47# 0.153f
C61 VPWR B2 0.00842f
C62 VGND a_193_297# 0.00438f
C63 VPWR B1 0.00982f
C64 A2 a_193_297# 0.00683f
C65 VPWR a_205_47# 1.62e-19
C66 a_109_297# C1 0.00739f
C67 A1 B1 0.0609f
C68 a_27_47# a_193_297# 0.144f
C69 VGND VNB 0.437f
C70 X VNB 0.0919f
C71 VPWR VNB 0.364f
C72 A2 VNB 0.0896f
C73 A1 VNB 0.106f
C74 B1 VNB 0.108f
C75 B2 VNB 0.0887f
C76 C1 VNB 0.139f
C77 VPB VNB 0.782f
C78 a_193_297# VNB 0.0011f
C79 a_109_297# VNB 7.11e-19
C80 a_27_47# VNB 0.216f
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X a_256_47# a_584_47#
+ a_93_21# a_250_297# a_346_47#
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
C0 VGND A1 0.0133f
C1 a_93_21# X 0.0841f
C2 VGND A3 0.00974f
C3 X a_250_297# 5.42e-19
C4 a_93_21# VPWR 0.0907f
C5 VPB a_93_21# 0.0485f
C6 a_346_47# a_93_21# 0.0119f
C7 VPWR a_250_297# 0.313f
C8 VPWR B2 0.0108f
C9 a_93_21# A2 0.0747f
C10 VPB a_250_297# 0.00616f
C11 VPB B2 0.0355f
C12 A2 a_250_297# 0.0129f
C13 A2 B2 1.46e-19
C14 A3 a_256_47# 4.42e-19
C15 a_93_21# B1 0.0774f
C16 a_250_297# B1 0.0125f
C17 B2 B1 0.0823f
C18 a_584_47# VGND 0.00683f
C19 VGND a_256_47# 0.00394f
C20 A1 X 6.03e-20
C21 A1 VPWR 0.016f
C22 VPB A1 0.0296f
C23 a_346_47# A1 0.00465f
C24 X A3 2.45e-19
C25 A1 A2 0.0971f
C26 A3 VPWR 0.0158f
C27 VPB A3 0.0291f
C28 VGND X 0.06f
C29 A1 B1 0.0965f
C30 A3 A2 0.0788f
C31 a_93_21# a_250_297# 0.188f
C32 a_93_21# B2 0.0147f
C33 VGND VPWR 0.076f
C34 VPB VGND 0.00788f
C35 a_250_297# B2 0.0344f
C36 a_346_47# VGND 0.00514f
C37 A3 B1 7.88e-22
C38 VGND A2 0.0114f
C39 VGND B1 0.0344f
C40 a_584_47# VPWR 9.47e-19
C41 a_256_47# VPWR 9.47e-19
C42 a_256_47# A2 0.00256f
C43 a_93_21# A1 0.0641f
C44 A1 a_250_297# 0.0129f
C45 A1 B2 3.14e-19
C46 a_584_47# B1 0.00143f
C47 a_256_47# B1 2.07e-20
C48 a_93_21# A3 0.124f
C49 A3 a_250_297# 0.00602f
C50 A3 B2 9.12e-20
C51 X VPWR 0.0849f
C52 VPB X 0.0108f
C53 X A2 1.19e-19
C54 a_93_21# VGND 0.251f
C55 VGND a_250_297# 0.0072f
C56 VGND B2 0.0469f
C57 VPB VPWR 0.0756f
C58 a_346_47# VPWR 0.00109f
C59 VPWR A2 0.0133f
C60 VPB A2 0.0287f
C61 a_346_47# A2 0.00252f
C62 X B1 3.83e-20
C63 a_584_47# a_93_21# 0.00278f
C64 VPWR B1 0.01f
C65 a_93_21# a_256_47# 0.0114f
C66 VPB B1 0.0276f
C67 a_584_47# a_250_297# 2.43e-19
C68 a_346_47# B1 5.39e-20
C69 A2 B1 1.44e-20
C70 VGND VNB 0.465f
C71 VPWR VNB 0.365f
C72 X VNB 0.0937f
C73 B2 VNB 0.14f
C74 B1 VNB 0.101f
C75 A1 VNB 0.0951f
C76 A2 VNB 0.0921f
C77 A3 VNB 0.0929f
C78 VPB VNB 0.782f
C79 a_250_297# VNB 0.0278f
C80 a_93_21# VNB 0.151f
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X a_277_297# a_205_297# a_27_297#
+ a_109_297#
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 VPWR a_109_297# 9.23e-19
C1 VGND D 0.0517f
C2 VGND a_277_297# 4.65e-19
C3 VGND C 0.0191f
C4 VPWR B 0.193f
C5 D VPB 0.0405f
C6 VPB C 0.0338f
C7 D a_27_297# 0.054f
C8 X a_277_297# 6.43e-20
C9 a_27_297# C 0.158f
C10 a_27_297# a_277_297# 0.00876f
C11 B A 0.0639f
C12 C a_205_297# 0.00261f
C13 VGND a_109_297# 7.58e-19
C14 VPWR A 0.00769f
C15 VGND B 0.0159f
C16 a_109_297# a_27_297# 0.00695f
C17 VGND VPWR 0.0546f
C18 B VPB 0.106f
C19 X B 6.42e-19
C20 B a_27_297# 0.159f
C21 D C 0.0954f
C22 VPWR VPB 0.075f
C23 C a_277_297# 5.54e-19
C24 X VPWR 0.0878f
C25 VPWR a_27_297# 0.084f
C26 VGND A 0.016f
C27 VPWR a_205_297# 5.16e-19
C28 A VPB 0.033f
C29 X A 0.00133f
C30 A a_27_297# 0.163f
C31 a_109_297# C 0.00356f
C32 D B 0.00287f
C33 VGND VPB 0.00796f
C34 VGND X 0.0354f
C35 B C 0.0917f
C36 B a_277_297# 2.29e-19
C37 VGND a_27_297# 0.235f
C38 D VPWR 0.00503f
C39 VPWR C 0.00723f
C40 VPWR a_277_297# 7.48e-19
C41 VGND a_205_297# 3.36e-19
C42 X VPB 0.0109f
C43 VPB a_27_297# 0.0517f
C44 X a_27_297# 0.0991f
C45 D A 2.13e-19
C46 A C 0.028f
C47 a_27_297# a_205_297# 0.00412f
C48 A a_277_297# 2.28e-19
C49 VGND VNB 0.367f
C50 X VNB 0.0883f
C51 A VNB 0.109f
C52 C VNB 0.105f
C53 D VNB 0.175f
C54 B VNB 0.115f
C55 VPWR VNB 0.29f
C56 VPB VNB 0.605f
C57 a_27_297# VNB 0.163f
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
C0 VGND VPWR 1.57f
C1 VGND VPB 0.35f
C2 VPB VPWR 0.137f
C3 VPWR VNB 1.67f
C4 VGND VNB 1.47f
C5 VPB VNB 1.14f
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X a_369_47# a_469_47#
+ a_297_47# a_193_413# a_27_47#
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VGND a_193_413# 0.0915f
C1 VGND a_27_47# 0.103f
C2 VPB VPWR 0.0818f
C3 a_27_47# a_193_413# 0.125f
C4 X VPWR 0.0586f
C5 C a_469_47# 0.00202f
C6 A_N VPWR 0.02f
C7 a_297_47# B 0.00353f
C8 VGND a_469_47# 0.00551f
C9 B a_369_47# 0.00129f
C10 B VPWR 0.0186f
C11 a_193_413# a_469_47# 0.00109f
C12 VPWR D 0.0186f
C13 VPB C 0.0742f
C14 C X 0.00479f
C15 VPB VGND 0.0123f
C16 VGND X 0.0588f
C17 VPB a_193_413# 0.0644f
C18 X a_193_413# 0.108f
C19 C B 0.164f
C20 VGND A_N 0.0205f
C21 VPB a_27_47# 0.092f
C22 VGND B 0.037f
C23 a_193_413# A_N 0.00151f
C24 C D 0.183f
C25 a_193_413# B 0.144f
C26 a_297_47# VPWR 2.82e-19
C27 VGND D 0.0372f
C28 a_27_47# A_N 0.237f
C29 a_369_47# VPWR 6.65e-19
C30 a_27_47# B 0.0794f
C31 a_193_413# D 0.155f
C32 X a_469_47# 0.001f
C33 C a_369_47# 0.00448f
C34 C VPWR 0.0182f
C35 VPB X 0.0108f
C36 a_297_47# VGND 0.00183f
C37 a_469_47# D 0.00183f
C38 VGND a_369_47# 0.00505f
C39 VGND VPWR 0.0727f
C40 a_297_47# a_193_413# 0.00137f
C41 VPB A_N 0.0832f
C42 a_193_413# a_369_47# 0.00181f
C43 a_193_413# VPWR 0.281f
C44 VPB B 0.089f
C45 a_27_47# VPWR 0.106f
C46 VPB D 0.0763f
C47 X D 0.0168f
C48 VGND C 0.0395f
C49 C a_193_413# 0.0389f
C50 a_469_47# VPWR 7.77e-19
C51 VGND VNB 0.456f
C52 X VNB 0.0934f
C53 VPWR VNB 0.368f
C54 D VNB 0.123f
C55 C VNB 0.108f
C56 B VNB 0.12f
C57 A_N VNB 0.198f
C58 VPB VNB 0.782f
C59 a_193_413# VNB 0.136f
C60 a_27_47# VNB 0.224f
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X a_109_93# a_368_53# a_209_311#
+ a_296_53#
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
C0 A_N C 7.6e-19
C1 VPWR X 0.0732f
C2 A_N B 2.03e-19
C3 VPWR VGND 0.0657f
C4 X VPB 0.0119f
C5 B C 0.0671f
C6 VPB VGND 0.00909f
C7 a_109_93# VGND 0.0784f
C8 X a_209_311# 0.0877f
C9 a_209_311# VGND 0.131f
C10 VGND a_368_53# 0.0031f
C11 VPWR a_296_53# 1.15e-19
C12 VPWR A_N 0.0513f
C13 A_N VPB 0.111f
C14 VPWR C 0.005f
C15 a_296_53# a_109_93# 1.84e-19
C16 VPB C 0.0339f
C17 a_296_53# a_209_311# 0.0049f
C18 A_N a_109_93# 0.117f
C19 VPWR B 0.131f
C20 A_N a_209_311# 0.00515f
C21 C a_109_93# 3.91e-20
C22 B VPB 0.0914f
C23 C a_209_311# 0.19f
C24 X VGND 0.0647f
C25 B a_109_93# 0.0802f
C26 B a_209_311# 0.0609f
C27 C a_368_53# 0.00415f
C28 a_296_53# VGND 6.07e-19
C29 VPWR VPB 0.104f
C30 X A_N 1.44e-19
C31 A_N VGND 0.045f
C32 X C 0.0176f
C33 VPWR a_109_93# 0.0984f
C34 C VGND 0.0678f
C35 VPWR a_209_311# 0.155f
C36 VPB a_109_93# 0.0652f
C37 VPB a_209_311# 0.0515f
C38 X B 0.00119f
C39 B VGND 0.00796f
C40 VPWR a_368_53# 4.26e-19
C41 a_109_93# a_209_311# 0.168f
C42 a_209_311# a_368_53# 0.0026f
C43 VGND VNB 0.44f
C44 X VNB 0.0925f
C45 C VNB 0.114f
C46 B VNB 0.101f
C47 VPWR VNB 0.342f
C48 A_N VNB 0.197f
C49 VPB VNB 0.693f
C50 a_209_311# VNB 0.143f
C51 a_109_93# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
C0 a_27_47# A 0.195f
C1 a_27_47# VPWR 0.219f
C2 VGND A 0.0431f
C3 VGND VPWR 0.057f
C4 VPB X 0.0122f
C5 a_27_47# VPB 0.139f
C6 VGND VPB 0.00583f
C7 A VPWR 0.022f
C8 a_27_47# X 0.328f
C9 VGND X 0.216f
C10 A VPB 0.0321f
C11 a_27_47# VGND 0.148f
C12 VPB VPWR 0.0632f
C13 A X 0.014f
C14 X VPWR 0.317f
C15 VGND VNB 0.358f
C16 X VNB 0.067f
C17 VPWR VNB 0.308f
C18 A VNB 0.148f
C19 VPB VNB 0.605f
C20 a_27_47# VNB 0.543f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
C0 a_59_75# VPB 0.0563f
C1 a_59_75# VPWR 0.15f
C2 VPB X 0.0127f
C3 X VPWR 0.111f
C4 VPB VGND 0.008f
C5 B VPB 0.0629f
C6 VGND VPWR 0.0461f
C7 B VPWR 0.0117f
C8 a_59_75# a_145_75# 0.00658f
C9 a_145_75# X 5.76e-19
C10 VPB VPWR 0.0729f
C11 a_145_75# VGND 0.00468f
C12 a_59_75# A 0.0809f
C13 X A 1.68e-19
C14 A VGND 0.0147f
C15 B A 0.0971f
C16 a_59_75# X 0.109f
C17 a_59_75# VGND 0.116f
C18 a_59_75# B 0.143f
C19 X VGND 0.0993f
C20 B X 0.00276f
C21 a_145_75# VPWR 6.31e-19
C22 B VGND 0.0115f
C23 VPB A 0.0806f
C24 A VPWR 0.0362f
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y a_297_297# a_191_297#
+ a_109_297#
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
C0 Y VPB 0.0127f
C1 A VGND 0.0526f
C2 A C 0.00268f
C3 VGND a_191_297# 9.29e-19
C4 Y VPWR 0.0561f
C5 a_191_297# C 0.0195f
C6 VGND a_297_297# 8.1e-19
C7 VPB B 0.0304f
C8 a_109_297# VGND 0.00181f
C9 a_109_297# C 0.0062f
C10 VPWR B 0.0887f
C11 VGND D 0.0456f
C12 C D 0.0523f
C13 A VPB 0.041f
C14 Y B 0.0403f
C15 A VPWR 0.0483f
C16 a_191_297# VPWR 0.0049f
C17 A Y 0.0175f
C18 VPWR a_297_297# 0.00317f
C19 a_109_297# VPWR 0.00576f
C20 Y a_191_297# 0.00142f
C21 VPB D 0.0376f
C22 VGND C 0.0184f
C23 Y a_297_297# 1.24e-19
C24 a_109_297# Y 0.0122f
C25 VPWR D 0.0128f
C26 A B 0.11f
C27 a_191_297# B 0.00223f
C28 Y D 0.108f
C29 B a_297_297# 0.0132f
C30 VGND VPB 0.0048f
C31 VPB C 0.0299f
C32 VGND VPWR 0.0492f
C33 A a_297_297# 3.16e-19
C34 VPWR C 0.0509f
C35 VGND Y 0.151f
C36 Y C 0.125f
C37 VGND B 0.0191f
C38 VPB VPWR 0.0524f
C39 B C 0.173f
C40 VGND VNB 0.322f
C41 VPWR VNB 0.276f
C42 Y VNB 0.0645f
C43 A VNB 0.174f
C44 B VNB 0.0968f
C45 C VNB 0.0911f
C46 D VNB 0.159f
C47 VPB VNB 0.516f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X a_75_212#
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 VPB VPWR 0.0355f
C1 VPB a_75_212# 0.0571f
C2 VPB VGND 0.00507f
C3 A X 8.48e-19
C4 VPB X 0.0128f
C5 VPB A 0.0525f
C6 VPWR VGND 0.0289f
C7 VPWR a_75_212# 0.134f
C8 VGND a_75_212# 0.105f
C9 VPWR X 0.0896f
C10 X VGND 0.0545f
C11 X a_75_212# 0.107f
C12 VPWR A 0.0217f
C13 A VGND 0.0184f
C14 A a_75_212# 0.178f
C15 VGND VNB 0.207f
C16 VPWR VNB 0.176f
C17 X VNB 0.0942f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_75_212# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 VPB X 0.0128f
C1 VPB VGND 0.00505f
C2 VPB a_27_47# 0.0592f
C3 A VPWR 0.0215f
C4 VPB VPWR 0.0355f
C5 VPB A 0.0524f
C6 X VGND 0.0546f
C7 X a_27_47# 0.107f
C8 VGND a_27_47# 0.105f
C9 X VPWR 0.0897f
C10 VPWR VGND 0.029f
C11 VPWR a_27_47# 0.135f
C12 X A 8.48e-19
C13 A VGND 0.0184f
C14 A a_27_47# 0.181f
C15 VGND VNB 0.207f
C16 X VNB 0.0941f
C17 VPWR VNB 0.175f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_27_47# VNB 0.208f
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X a_664_47# a_841_47#
+ a_381_47# a_62_47# a_558_47#
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_558_47# VPB 0.115f
C1 a_664_47# a_841_47# 0.134f
C2 VPWR VPB 0.103f
C3 VPWR a_62_47# 0.149f
C4 VGND VPB 0.008f
C5 VGND a_62_47# 0.144f
C6 X VPB 0.126f
C7 X a_62_47# 0.156f
C8 VPB A 0.105f
C9 a_62_47# A 0.244f
C10 a_558_47# a_841_47# 0.00368f
C11 VPWR a_841_47# 0.0614f
C12 a_558_47# a_664_47# 0.314f
C13 a_841_47# VGND 0.0585f
C14 a_664_47# VPWR 0.131f
C15 a_664_47# VGND 0.125f
C16 VPB a_62_47# 0.0515f
C17 X a_664_47# 6.67e-19
C18 a_558_47# a_381_47# 0.16f
C19 VPWR a_381_47# 0.134f
C20 a_381_47# VGND 0.125f
C21 X a_381_47# 0.318f
C22 a_558_47# VPWR 0.084f
C23 a_381_47# A 5.42e-19
C24 a_558_47# VGND 0.0816f
C25 a_558_47# X 0.0144f
C26 a_841_47# VPB 0.0108f
C27 VPWR VGND 0.0902f
C28 X VPWR 0.108f
C29 a_664_47# VPB 0.043f
C30 X VGND 0.106f
C31 VPWR A 0.0174f
C32 VGND A 0.0176f
C33 X A 0.0142f
C34 a_381_47# VPB 0.0447f
C35 VGND VNB 0.537f
C36 VPWR VNB 0.439f
C37 X VNB 0.163f
C38 A VNB 0.198f
C39 VPB VNB 0.959f
C40 a_841_47# VNB 0.0929f
C41 a_664_47# VNB 0.13f
C42 a_558_47# VNB 0.164f
C43 a_381_47# VNB 0.11f
C44 a_62_47# VNB 0.169f
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y a_129_47# a_47_47# a_285_47#
+ a_377_297#
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VGND A 0.0635f
C1 VGND VPWR 0.0665f
C2 VGND a_47_47# 0.104f
C3 A a_285_47# 0.0353f
C4 a_285_47# a_47_47# 0.0175f
C5 a_285_47# VPWR 0.00255f
C6 B Y 0.00334f
C7 A VPB 0.0822f
C8 a_129_47# a_47_47# 0.00369f
C9 a_129_47# VPWR 9.47e-19
C10 VPB a_47_47# 0.0444f
C11 VPB VPWR 0.0718f
C12 a_47_47# a_377_297# 0.00899f
C13 VPWR a_377_297# 0.00559f
C14 VGND B 0.0389f
C15 B a_285_47# 0.067f
C16 a_129_47# B 0.00236f
C17 B VPB 0.0643f
C18 B a_377_297# 0.00254f
C19 A a_47_47# 0.0307f
C20 A VPWR 0.0349f
C21 a_47_47# VPWR 0.273f
C22 VGND Y 0.0381f
C23 a_285_47# Y 0.0439f
C24 Y VPB 0.00878f
C25 A B 0.236f
C26 B a_47_47# 0.356f
C27 B VPWR 0.0408f
C28 VGND a_285_47# 0.211f
C29 Y a_377_297# 0.00188f
C30 VGND a_129_47# 0.00547f
C31 VGND VPB 0.00568f
C32 a_285_47# VPB 5.53e-19
C33 VGND a_377_297# 0.00125f
C34 A Y 0.00181f
C35 Y a_47_47# 0.143f
C36 Y VPWR 0.107f
C37 VGND VNB 0.4f
C38 Y VNB 0.0783f
C39 VPWR VNB 0.352f
C40 A VNB 0.217f
C41 B VNB 0.212f
C42 VPB VNB 0.693f
C43 a_285_47# VNB 0.0174f
C44 a_47_47# VNB 0.199f
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X a_472_297# a_80_21#
+ a_300_47# a_217_297#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
C0 VPB a_80_21# 0.0661f
C1 a_217_297# VPWR 0.197f
C2 VPB A2 0.0384f
C3 VPWR B1 0.0129f
C4 VPWR a_472_297# 0.00703f
C5 a_217_297# VGND 0.00342f
C6 a_80_21# a_300_47# 0.00997f
C7 X a_217_297# 0.00271f
C8 VGND B1 0.0175f
C9 VGND a_472_297# 0.00188f
C10 a_217_297# A1 0.0124f
C11 X B1 1.18e-19
C12 X a_472_297# 2.6e-19
C13 A1 B1 0.0834f
C14 a_217_297# C1 0.00262f
C15 B1 C1 0.0846f
C16 a_80_21# VPWR 0.119f
C17 a_80_21# VGND 0.293f
C18 X a_80_21# 0.118f
C19 VPWR A2 0.0161f
C20 a_80_21# A1 0.111f
C21 A2 VGND 0.0191f
C22 X A2 6.82e-19
C23 VPB VPWR 0.0754f
C24 a_80_21# C1 0.079f
C25 A2 A1 0.0881f
C26 a_217_297# B1 0.00651f
C27 a_217_297# a_472_297# 0.00517f
C28 VPB VGND 0.00775f
C29 B1 a_472_297# 1.87e-19
C30 X VPB 0.0118f
C31 VPB A1 0.0266f
C32 VPWR a_300_47# 8.53e-19
C33 VPB C1 0.0379f
C34 a_300_47# VGND 0.00536f
C35 X a_300_47# 5.31e-19
C36 a_300_47# A1 5.95e-19
C37 a_217_297# a_80_21# 0.127f
C38 a_80_21# B1 0.0964f
C39 a_80_21# a_472_297# 0.0164f
C40 a_217_297# A2 0.0135f
C41 VPWR VGND 0.0665f
C42 X VPWR 0.0884f
C43 VPWR A1 0.0149f
C44 a_217_297# VPB 0.00494f
C45 VPB B1 0.0267f
C46 X VGND 0.0654f
C47 VGND A1 0.0147f
C48 X A1 3.62e-19
C49 VPWR C1 0.0137f
C50 VGND C1 0.0176f
C51 X C1 7.15e-20
C52 a_80_21# A2 0.128f
C53 VGND VNB 0.385f
C54 VPWR VNB 0.325f
C55 X VNB 0.0899f
C56 C1 VNB 0.144f
C57 B1 VNB 0.0899f
C58 A1 VNB 0.0905f
C59 A2 VNB 0.108f
C60 VPB VNB 0.693f
C61 a_217_297# VNB 0.00117f
C62 a_80_21# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
C0 B C 0.161f
C1 VGND D 0.0898f
C2 VGND VPWR 0.0662f
C3 VGND a_197_47# 0.00387f
C4 D VPB 0.0782f
C5 B a_27_47# 0.13f
C6 VPB VPWR 0.077f
C7 A VPWR 0.044f
C8 a_109_47# VPWR 4.66e-19
C9 a_27_47# X 0.0754f
C10 D a_303_47# 0.00119f
C11 VPWR a_303_47# 4.83e-19
C12 VGND C 0.0408f
C13 C VPB 0.0609f
C14 VGND a_27_47# 0.132f
C15 VPB a_27_47# 0.082f
C16 C a_109_47# 1.72e-20
C17 VGND B 0.0453f
C18 a_27_47# A 0.153f
C19 B VPB 0.0643f
C20 C a_303_47# 0.00527f
C21 a_27_47# a_109_47# 0.00578f
C22 D VPWR 0.0207f
C23 B A 0.0839f
C24 a_197_47# VPWR 5.24e-19
C25 B a_109_47# 0.00153f
C26 a_27_47# a_303_47# 0.00119f
C27 VGND X 0.0903f
C28 VPB X 0.0111f
C29 D C 0.18f
C30 C a_197_47# 0.00123f
C31 C VPWR 0.021f
C32 VGND VPB 0.00852f
C33 D a_27_47# 0.107f
C34 VGND A 0.0151f
C35 a_27_47# a_197_47# 0.00167f
C36 a_27_47# VPWR 0.326f
C37 VGND a_109_47# 0.00223f
C38 VPB A 0.0907f
C39 B a_197_47# 0.00623f
C40 B VPWR 0.0231f
C41 VGND a_303_47# 0.00381f
C42 D X 0.00746f
C43 C a_27_47# 0.0516f
C44 X VPWR 0.0945f
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X a_489_413# a_226_47#
+ a_556_47# a_226_297# a_76_199#
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_226_47# a_489_413# 0.00579f
C1 VPB VPWR 0.0951f
C2 B2 VPWR 0.0161f
C3 B2 a_556_47# 0.00291f
C4 a_489_413# VGND 0.0058f
C5 a_226_297# a_76_199# 0.00354f
C6 a_76_199# VPWR 0.2f
C7 a_76_199# a_556_47# 0.0017f
C8 A2_N VPWR 0.00449f
C9 X VPWR 0.0589f
C10 B1 VGND 0.0471f
C11 a_226_297# A1_N 0.00184f
C12 VPWR A1_N 0.00672f
C13 VPB a_489_413# 0.015f
C14 a_226_47# VGND 0.149f
C15 a_489_413# B2 0.0541f
C16 VPB B1 0.0803f
C17 a_489_413# a_76_199# 0.0473f
C18 B2 B1 0.182f
C19 VPB a_226_47# 0.111f
C20 B1 a_76_199# 0.00185f
C21 a_226_47# B2 0.0975f
C22 a_226_297# VPWR 8.54e-19
C23 a_226_47# a_76_199# 0.188f
C24 VPWR a_556_47# 7.24e-19
C25 A2_N a_226_47# 0.141f
C26 a_226_47# X 0.0108f
C27 VPB VGND 0.0128f
C28 B2 VGND 0.0335f
C29 a_226_47# A1_N 0.0209f
C30 VGND a_76_199# 0.108f
C31 A2_N VGND 0.0174f
C32 VGND X 0.0627f
C33 a_489_413# VPWR 0.143f
C34 VPB B2 0.0645f
C35 VGND A1_N 0.0261f
C36 VPB a_76_199# 0.0817f
C37 VPB A2_N 0.0327f
C38 B1 VPWR 0.0188f
C39 VPB X 0.0113f
C40 B2 a_76_199# 0.0626f
C41 a_226_297# a_226_47# 0.00128f
C42 a_226_47# VPWR 0.0187f
C43 VPB A1_N 0.0339f
C44 A2_N a_76_199# 0.0125f
C45 a_76_199# X 0.0995f
C46 A2_N X 2.55e-19
C47 a_226_297# VGND 5.63e-19
C48 a_76_199# A1_N 0.119f
C49 A2_N A1_N 0.11f
C50 VGND VPWR 0.0743f
C51 VGND a_556_47# 0.00639f
C52 a_489_413# B1 0.0382f
C53 X A1_N 0.00211f
C54 VGND VNB 0.462f
C55 A2_N VNB 0.103f
C56 A1_N VNB 0.111f
C57 VPWR VNB 0.369f
C58 X VNB 0.0975f
C59 B1 VNB 0.206f
C60 B2 VNB 0.106f
C61 VPB VNB 0.782f
C62 a_489_413# VNB 0.0254f
C63 a_226_47# VNB 0.162f
C64 a_76_199# VNB 0.141f
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X a_515_93# a_223_47#
+ a_615_93# a_343_93# a_429_93# a_27_47#
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
C0 B_N C 9.56e-20
C1 VGND C 0.025f
C2 VPB D 0.081f
C3 VPB VPWR 0.106f
C4 B_N a_223_47# 0.0431f
C5 VGND a_223_47# 0.199f
C6 a_27_47# VPWR 0.0897f
C7 a_615_93# D 0.00564f
C8 A_N VPWR 0.0318f
C9 D a_343_93# 0.114f
C10 VGND B_N 0.0427f
C11 a_615_93# VPWR 8.49e-19
C12 a_343_93# a_429_93# 0.00484f
C13 a_343_93# VPWR 0.255f
C14 VPWR a_515_93# 7.86e-19
C15 VPB C 0.0686f
C16 B_N X 4.64e-20
C17 VGND X 0.0609f
C18 VPB a_223_47# 0.0799f
C19 a_615_93# C 0.00407f
C20 a_27_47# a_223_47# 0.267f
C21 C a_343_93# 0.0397f
C22 VPB B_N 0.0646f
C23 VPB VGND 0.0167f
C24 a_223_47# A_N 0.00833f
C25 B_N a_27_47# 0.138f
C26 C a_515_93# 0.00389f
C27 a_223_47# a_343_93# 0.269f
C28 VGND a_27_47# 0.0715f
C29 D VPWR 0.0143f
C30 B_N A_N 0.117f
C31 a_429_93# VPWR 5.19e-19
C32 VGND A_N 0.0146f
C33 B_N a_343_93# 0.00112f
C34 a_223_47# a_515_93# 0.00482f
C35 VGND a_615_93# 0.0044f
C36 VPB X 0.0103f
C37 VGND a_343_93# 0.0548f
C38 VGND a_515_93# 0.00408f
C39 X a_343_93# 0.126f
C40 D C 0.163f
C41 C VPWR 0.012f
C42 VPB a_27_47# 0.154f
C43 D a_223_47# 4.03e-19
C44 VPB A_N 0.0848f
C45 a_223_47# a_429_93# 0.00492f
C46 a_223_47# VPWR 0.114f
C47 VPB a_343_93# 0.0857f
C48 a_27_47# A_N 0.0906f
C49 a_27_47# a_343_93# 0.0406f
C50 D B_N 6.67e-20
C51 VGND D 0.0414f
C52 B_N VPWR 0.0168f
C53 VGND a_429_93# 0.00122f
C54 VGND VPWR 0.0906f
C55 a_615_93# a_343_93# 0.00103f
C56 D X 0.0193f
C57 C a_223_47# 0.151f
C58 a_343_93# a_515_93# 0.00115f
C59 X VPWR 0.0582f
C60 VGND VNB 0.553f
C61 X VNB 0.0908f
C62 VPWR VNB 0.453f
C63 D VNB 0.124f
C64 C VNB 0.107f
C65 B_N VNB 0.134f
C66 A_N VNB 0.144f
C67 VPB VNB 0.959f
C68 a_343_93# VNB 0.172f
C69 a_223_47# VNB 0.141f
C70 a_27_47# VNB 0.259f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 B a_285_297# 0.0553f
C1 a_285_47# VPWR 8.6e-19
C2 a_117_297# X 2.25e-19
C3 B X 0.0149f
C4 a_285_47# a_35_297# 0.00723f
C5 a_285_297# VPB 0.0133f
C6 a_285_47# VGND 0.00552f
C7 B a_117_297# 0.00777f
C8 X VPB 0.0154f
C9 A a_285_297# 0.00749f
C10 B VPB 0.0697f
C11 a_285_297# VPWR 0.246f
C12 A X 0.00166f
C13 a_285_297# a_35_297# 0.025f
C14 VPWR X 0.0537f
C15 a_285_297# VGND 0.00394f
C16 A B 0.221f
C17 X a_35_297# 0.166f
C18 a_117_297# VPWR 0.00852f
C19 X VGND 0.173f
C20 B VPWR 0.0703f
C21 a_117_297# a_35_297# 0.00641f
C22 B a_35_297# 0.203f
C23 a_117_297# VGND 0.00177f
C24 A VPB 0.051f
C25 B VGND 0.0304f
C26 VPWR VPB 0.0689f
C27 VPB a_35_297# 0.0699f
C28 VPB VGND 0.00696f
C29 A VPWR 0.0348f
C30 a_285_47# X 0.00206f
C31 A a_35_297# 0.0633f
C32 A VGND 0.0325f
C33 VPWR a_35_297# 0.096f
C34 VPWR VGND 0.0643f
C35 B a_285_47# 3.98e-19
C36 a_35_297# VGND 0.177f
C37 a_285_297# X 0.0712f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X a_465_297# a_297_297#
+ a_215_297# a_392_297# a_109_53#
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 VPWR A 0.0073f
C1 VPWR X 0.0885f
C2 VPWR a_392_297# 5.29e-19
C3 A a_215_297# 0.157f
C4 D_N a_109_53# 0.0889f
C5 a_215_297# a_392_297# 0.00419f
C6 a_215_297# X 0.0991f
C7 C VPB 0.0337f
C8 A B 0.0666f
C9 C VGND 0.0202f
C10 B X 6.65e-19
C11 a_109_53# VPB 0.0547f
C12 a_109_53# VGND 0.118f
C13 A a_465_297# 5.42e-19
C14 VPWR C 0.00753f
C15 D_N VPB 0.0461f
C16 D_N VGND 0.0531f
C17 C a_215_297# 0.161f
C18 VPWR a_109_53# 0.0418f
C19 C B 0.0893f
C20 a_215_297# a_109_53# 0.0807f
C21 C a_297_297# 0.00375f
C22 VGND VPB 0.0115f
C23 VPWR D_N 0.0412f
C24 a_109_53# B 0.0246f
C25 D_N a_215_297# 3.19e-19
C26 C a_465_297# 6.89e-19
C27 a_109_53# a_297_297# 7.06e-21
C28 A X 0.00127f
C29 VPWR VPB 0.122f
C30 VPWR VGND 0.075f
C31 a_215_297# VPB 0.0508f
C32 a_215_297# VGND 0.237f
C33 VPB B 0.116f
C34 VGND B 0.0161f
C35 VGND a_297_297# 6.5e-19
C36 A C 0.0281f
C37 C a_392_297# 0.00267f
C38 VPWR a_215_297# 0.0871f
C39 VGND a_465_297# 5.02e-19
C40 A a_109_53# 1.19e-19
C41 VPWR B 0.255f
C42 VPWR a_297_297# 8.59e-19
C43 a_215_297# B 0.159f
C44 a_215_297# a_297_297# 0.00659f
C45 VPWR a_465_297# 7.08e-19
C46 a_215_297# a_465_297# 0.00827f
C47 A VPB 0.0325f
C48 A VGND 0.0158f
C49 VPB X 0.011f
C50 C a_109_53# 0.0984f
C51 VGND a_392_297# 3.44e-19
C52 VGND X 0.0359f
C53 VGND VNB 0.469f
C54 X VNB 0.0884f
C55 A VNB 0.108f
C56 C VNB 0.101f
C57 D_N VNB 0.185f
C58 B VNB 0.101f
C59 VPWR VNB 0.399f
C60 VPB VNB 0.782f
C61 a_109_53# VNB 0.159f
C62 a_215_297# VNB 0.142f
.ends

.subckt therm_port_resized VGND VPWR b[0] b[1] b[2] b[3] p[0] p[10] p[11] p[12] p[13]
+ p[14] p[1] p[2] p[3] p[4] p[5] p[6] p[7] p[8] p[9]
X_49_ net7 _02_ _19_ _20_ _21_ VGND VGND VPWR VPWR net17 _49_/a_208_47# _49_/a_75_199#
+ _49_/a_544_297# _49_/a_315_47# _49_/a_201_297# sky130_fd_sc_hd__a311o_1
X_48_ net11 _02_ _07_ VGND VGND VPWR VPWR _21_ _48_/a_181_47# _48_/a_109_47# _48_/a_27_47#
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ net5 _12_ _17_ VGND VGND VPWR VPWR _20_ _47_/a_384_47# _47_/a_81_21# _47_/a_299_297#
+ sky130_fd_sc_hd__a21o_1
X_46_ _04_ VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__inv_2
X_29_ net11 net13 net12 VGND VGND VPWR VPWR _03_ _29_/a_29_53# _29_/a_183_297# _29_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_28_ _00_ _01_ VGND VGND VPWR VPWR _02_ _28_/a_109_297# sky130_fd_sc_hd__nor2_1
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_45_ _02_ _09_ _12_ _13_ _18_ VGND VGND VPWR VPWR net16 _45_/a_193_297# _45_/a_465_47#
+ _45_/a_205_47# _45_/a_109_297# _45_/a_27_47# sky130_fd_sc_hd__a221o_1
X_44_ net14 _14_ _15_ _17_ net2 VGND VGND VPWR VPWR _18_ _44_/a_256_47# _44_/a_584_47#
+ _44_/a_93_21# _44_/a_250_297# _44_/a_346_47# sky130_fd_sc_hd__a32o_1
X_27_ net14 net15 net3 net2 VGND VGND VPWR VPWR _01_ _27_/a_277_297# _27_/a_205_297#
+ _27_/a_27_297# _27_/a_109_297# sky130_fd_sc_hd__or4_1
XFILLER_0_7_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_26_ net5 net4 net6 VGND VGND VPWR VPWR _00_ _26_/a_29_53# _26_/a_183_297# _26_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_43_ _00_ _06_ _10_ _16_ VGND VGND VPWR VPWR _17_ _43_/a_369_47# _43_/a_469_47# _43_/a_297_47#
+ _43_/a_193_413# _43_/a_27_47# sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_42_ net3 net15 net14 VGND VGND VPWR VPWR _16_ _42_/a_109_93# _42_/a_368_53# _42_/a_209_311#
+ _42_/a_296_53# sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_3_Left_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND VPWR VPWR b[0] output16/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_41_ _06_ _10_ VGND VGND VPWR VPWR _15_ _41_/a_145_75# _41_/a_59_75# sky130_fd_sc_hd__and2_1
Xoutput17 net17 VGND VGND VPWR VPWR b[1] output17/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_40_ net15 net3 net2 _00_ VGND VGND VPWR VPWR _14_ _40_/a_297_297# _40_/a_191_297#
+ _40_/a_109_297# sky130_fd_sc_hd__nor4_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput18 net18 VGND VGND VPWR VPWR b[2] output18/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_0_Left_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR b[3] output19/a_27_47# sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 p[0] VGND VGND VPWR VPWR net1 input1/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput2 p[10] VGND VGND VPWR VPWR net2 input2/a_27_47# sky130_fd_sc_hd__buf_1
Xinput3 p[11] VGND VGND VPWR VPWR net3 input3/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 p[12] VGND VGND VPWR VPWR net4 input4/a_75_212# sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 p[13] VGND VGND VPWR VPWR net5 input5/a_664_47# input5/a_841_47# input5/a_381_47#
+ input5/a_62_47# input5/a_558_47# sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_1_Left_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 p[14] VGND VGND VPWR VPWR net6 input6/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 p[1] VGND VGND VPWR VPWR net7 input7/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput10 p[4] VGND VGND VPWR VPWR net10 input10/a_27_47# sky130_fd_sc_hd__buf_1
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 p[2] VGND VGND VPWR VPWR net8 input8/a_27_47# sky130_fd_sc_hd__buf_1
Xinput11 p[5] VGND VGND VPWR VPWR net11 input11/a_27_47# sky130_fd_sc_hd__buf_1
X_39_ net5 net6 VGND VGND VPWR VPWR _13_ _39_/a_129_47# _39_/a_47_47# _39_/a_285_47#
+ _39_/a_377_297# sky130_fd_sc_hd__xnor2_1
Xinput9 p[3] VGND VGND VPWR VPWR net9 input9/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput12 p[6] VGND VGND VPWR VPWR net12 input12/a_27_47# sky130_fd_sc_hd__buf_1
X_55_ _14_ _15_ _20_ _22_ VGND VGND VPWR VPWR net19 _55_/a_472_297# _55_/a_80_21#
+ _55_/a_300_47# _55_/a_217_297# sky130_fd_sc_hd__a211o_1
X_38_ net4 _06_ _10_ _11_ VGND VGND VPWR VPWR _12_ _38_/a_109_47# _38_/a_197_47# _38_/a_303_47#
+ _38_/a_27_47# sky130_fd_sc_hd__and4_1
X_54_ _25_ VGND VGND VPWR VPWR net18 _54_/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput13 p[7] VGND VGND VPWR VPWR net13 input13/a_27_47# sky130_fd_sc_hd__buf_1
X_37_ net14 net15 net3 net2 VGND VGND VPWR VPWR _11_ _37_/a_109_47# _37_/a_197_47#
+ _37_/a_303_47# _37_/a_27_47# sky130_fd_sc_hd__and4_1
Xinput14 p[8] VGND VGND VPWR VPWR net14 input14/a_27_47# sky130_fd_sc_hd__buf_1
X_53_ _21_ _22_ _24_ VGND VGND VPWR VPWR _25_ _53_/a_29_53# _53_/a_183_297# _53_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_36_ net11 net10 net13 net12 VGND VGND VPWR VPWR _10_ _36_/a_109_47# _36_/a_197_47#
+ _36_/a_303_47# _36_/a_27_47# sky130_fd_sc_hd__and4_1
X_52_ _02_ _06_ _23_ _12_ net5 VGND VGND VPWR VPWR _24_ _52_/a_256_47# _52_/a_584_47#
+ _52_/a_93_21# _52_/a_250_297# _52_/a_346_47# sky130_fd_sc_hd__a32o_1
Xinput15 p[9] VGND VGND VPWR VPWR net15 input15/a_27_47# sky130_fd_sc_hd__buf_1
X_35_ _04_ _05_ _07_ _08_ VGND VGND VPWR VPWR _09_ _35_/a_489_413# _35_/a_226_47#
+ _35_/a_556_47# _35_/a_226_297# _35_/a_76_199# sky130_fd_sc_hd__a2bb2o_1
X_51_ _03_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__inv_2
X_34_ net11 net12 VGND VGND VPWR VPWR _08_ _34_/a_129_47# _34_/a_47_47# _34_/a_285_47#
+ _34_/a_377_297# sky130_fd_sc_hd__xnor2_1
X_33_ net13 _06_ net10 VGND VGND VPWR VPWR _07_ _33_/a_109_93# _33_/a_368_53# _33_/a_209_311#
+ _33_/a_296_53# sky130_fd_sc_hd__and3b_1
X_50_ net5 net6 _15_ _11_ VGND VGND VPWR VPWR _22_ _50_/a_515_93# _50_/a_223_47# _50_/a_615_93#
+ _50_/a_343_93# _50_/a_429_93# _50_/a_27_47# sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ net7 net1 net9 net8 VGND VGND VPWR VPWR _06_ _32_/a_109_47# _32_/a_197_47# _32_/a_303_47#
+ _32_/a_27_47# sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_5_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31_ net7 net8 VGND VGND VPWR VPWR _05_ _31_/a_117_297# _31_/a_285_297# _31_/a_285_47#
+ _31_/a_35_297# sky130_fd_sc_hd__xor2_1
X_30_ net9 net10 _03_ net1 VGND VGND VPWR VPWR _04_ _30_/a_465_297# _30_/a_297_297#
+ _30_/a_215_297# _30_/a_392_297# _30_/a_109_53# sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
C0 net9 input8/a_27_47# 3.71e-20
C1 _36_/a_27_47# net1 6.99e-20
C2 _40_/a_109_297# net6 2.53e-20
C3 _36_/a_27_47# net6 5.1e-19
C4 VGND _10_ 1.11f
C5 net14 input5/a_558_47# 0.0325f
C6 net3 input5/a_664_47# 0.00215f
C7 net11 _09_ 0.0262f
C8 _17_ _37_/a_303_47# 1.23e-20
C9 net16 net4 0.155f
C10 _44_/a_250_297# _04_ 5.57e-21
C11 net17 net9 1.26e-20
C12 net1 _27_/a_27_297# 6.05e-21
C13 _11_ _50_/a_27_47# 0.0592f
C14 p[7] VPWR 0.0176f
C15 net15 p[12] 2.99e-19
C16 _50_/a_615_93# _15_ 0.00183f
C17 net7 VPWR 0.78f
C18 net4 _22_ 0.0866f
C19 p[6] b[1] 0.00407f
C20 _53_/a_183_297# _10_ 2.86e-19
C21 input7/a_27_47# input8/a_27_47# 3.2e-20
C22 _31_/a_35_297# VPWR 0.0284f
C23 _34_/a_377_297# VGND -0.00102f
C24 net12 _18_ 2.25e-21
C25 _35_/a_489_413# _03_ 0.0205f
C26 _16_ VPWR 0.126f
C27 net17 input7/a_27_47# 4.99e-20
C28 input5/a_841_47# _02_ 0.00591f
C29 _36_/a_197_47# _06_ 6.18e-19
C30 _35_/a_76_199# net6 4.6e-21
C31 _37_/a_27_47# _44_/a_93_21# 3.19e-19
C32 _17_ _02_ 0.00482f
C33 net10 _39_/a_47_47# 4.72e-22
C34 net3 _55_/a_80_21# 2.35e-19
C35 output19/a_27_47# _44_/a_93_21# 7.25e-20
C36 net1 net9 0.47f
C37 VGND net18 0.255f
C38 _45_/a_27_47# net6 0.021f
C39 _48_/a_27_47# _07_ 0.0524f
C40 _29_/a_29_53# _21_ 0.0775f
C41 VPWR _47_/a_81_21# 0.00889f
C42 _10_ p[12] 0.0994f
C43 net7 net11 1.77e-19
C44 p[8] p[11] 0.00244f
C45 _43_/a_297_47# _00_ 1.26e-19
C46 net13 net5 0.127f
C47 _17_ _42_/a_209_311# 1.22e-19
C48 VGND _38_/a_303_47# 1.78e-19
C49 _43_/a_193_413# net8 1.62e-20
C50 _50_/a_27_47# _02_ 2.09e-19
C51 _13_ net6 0.0106f
C52 net1 input7/a_27_47# 0.0383f
C53 p[13] net5 0.00689f
C54 p[1] net7 0.00514f
C55 p[8] input3/a_27_47# 6.2e-19
C56 _50_/a_429_93# _10_ 0.00167f
C57 _29_/a_111_297# _04_ 9.25e-19
C58 _01_ _32_/a_197_47# 0.00156f
C59 VGND _35_/a_489_413# -8.78e-19
C60 _23_ _07_ 1.27e-19
C61 _43_/a_193_413# input15/a_27_47# 1.62e-20
C62 net14 _27_/a_205_297# 3.63e-19
C63 _33_/a_296_53# VGND -1.43e-19
C64 _26_/a_183_297# _22_ 0.00184f
C65 _12_ _43_/a_27_47# 2.33e-21
C66 p[11] _42_/a_109_93# 1.48e-19
C67 _36_/a_27_47# _20_ 0.00148f
C68 net13 net12 0.363f
C69 _20_ _40_/a_109_297# 2.35e-20
C70 input5/a_381_47# net17 1.37e-20
C71 _49_/a_544_297# _04_ 0.00204f
C72 _36_/a_27_47# b[1] 7.95e-19
C73 _06_ _52_/a_256_47# 0.00207f
C74 _30_/a_215_297# _21_ 1.48e-19
C75 input4/a_75_212# _41_/a_59_75# 0.00153f
C76 _20_ _27_/a_27_297# 3.14e-20
C77 _17_ _55_/a_80_21# 7.64e-21
C78 _26_/a_29_53# net5 0.0237f
C79 net3 net14 0.689f
C80 _43_/a_27_47# _22_ 0.091f
C81 _27_/a_27_297# b[1] 0.00644f
C82 p[2] _02_ 7.38e-19
C83 input3/a_27_47# _42_/a_109_93# 0.00249f
C84 net1 _00_ 9.43e-19
C85 net6 _00_ 0.00178f
C86 input5/a_558_47# p[10] 1.09e-19
C87 p[7] p[4] 7.8e-20
C88 _10_ _29_/a_183_297# 6.24e-20
C89 _33_/a_209_311# _35_/a_226_47# 1.31e-19
C90 output17/a_27_47# _03_ 1.94e-19
C91 p[2] _05_ 3.82e-19
C92 input2/a_27_47# _27_/a_27_297# 1.16e-19
C93 _18_ _43_/a_193_413# 0.0413f
C94 _50_/a_343_93# _11_ 0.0384f
C95 input6/a_27_47# input15/a_27_47# 5.3e-19
C96 _35_/a_76_199# _20_ 3.21e-20
C97 _44_/a_250_297# _42_/a_109_93# 6.38e-19
C98 p[8] input14/a_27_47# 0.0109f
C99 _53_/a_111_297# _02_ 9.57e-20
C100 _35_/a_76_199# b[1] 0.00458f
C101 net6 _52_/a_93_21# 2.33e-19
C102 VGND input5/a_558_47# -0.00123f
C103 net1 input5/a_381_47# 1.27e-19
C104 _12_ VPWR 0.28f
C105 _20_ net9 0.328f
C106 _36_/a_109_47# VPWR -4.66e-19
C107 _40_/a_191_297# VPWR -6.82e-19
C108 VPWR _40_/a_297_297# -5.42e-19
C109 b[3] _41_/a_59_75# 9.66e-22
C110 net1 _32_/a_303_47# 1.45e-19
C111 net9 b[1] 0.0765f
C112 net12 _26_/a_29_53# 6.55e-19
C113 _15_ _37_/a_197_47# 3.02e-19
C114 _28_/a_109_297# _14_ 5.66e-19
C115 net16 VPWR 0.518f
C116 _29_/a_29_53# _30_/a_215_297# 1.72e-19
C117 net10 _50_/a_27_47# 3.78e-21
C118 output17/a_27_47# p[10] 0.117f
C119 input5/a_62_47# _19_ 0.00159f
C120 _53_/a_29_53# net6 2.11e-20
C121 _22_ VPWR 1.4f
C122 _13_ _20_ 7.38e-21
C123 _11_ _02_ 0.0621f
C124 net15 _06_ 0.033f
C125 _27_/a_205_297# _03_ 1.46e-20
C126 net5 _14_ 3.89e-19
C127 p[7] input12/a_27_47# 1.07e-19
C128 _12_ net11 0.00799f
C129 _39_/a_47_47# _03_ 1.47e-19
C130 VGND b[0] 0.181f
C131 input7/a_27_47# b[1] 0.00663f
C132 VGND output17/a_27_47# 0.00231f
C133 _50_/a_343_93# _02_ 6.94e-19
C134 _32_/a_27_47# _10_ 0.00217f
C135 net14 _17_ 0.104f
C136 p[3] _30_/a_109_53# 1.27e-19
C137 net15 _47_/a_299_297# 1.44e-20
C138 net16 net11 4.43e-22
C139 _27_/a_27_297# _15_ 9.85e-20
C140 _18_ net4 0.023f
C141 input2/a_27_47# input7/a_27_47# 1.62e-19
C142 net3 _03_ 4.27e-20
C143 _04_ VPWR 0.456f
C144 _45_/a_193_297# net4 7.41e-19
C145 _45_/a_109_297# net6 7.82e-19
C146 net11 _22_ 6.82e-21
C147 _10_ _06_ 1.14f
C148 input10/a_27_47# p[6] 0.00214f
C149 _19_ _49_/a_75_199# 0.0206f
C150 p[13] p[11] 0.0137f
C151 output18/a_27_47# output16/a_27_47# 7.85e-19
C152 net5 _21_ 0.00784f
C153 net5 net19 0.00124f
C154 _45_/a_205_47# _12_ 7.46e-19
C155 net1 _09_ 5.26e-20
C156 _33_/a_368_53# _05_ 9.2e-19
C157 _20_ _00_ 0.271f
C158 _26_/a_29_53# _24_ 2.11e-20
C159 net6 _09_ 5.43e-20
C160 net7 input8/a_27_47# 1.47e-19
C161 _35_/a_226_47# _07_ 8.96e-19
C162 _36_/a_303_47# VGND 8.14e-19
C163 _47_/a_299_297# _10_ 0.0134f
C164 p[8] p[14] 0.00121f
C165 p[13] input3/a_27_47# 0.00527f
C166 net11 _04_ 0.078f
C167 _15_ net9 0.00113f
C168 _31_/a_35_297# input8/a_27_47# 0.00955f
C169 _34_/a_377_297# _06_ 0.00427f
C170 _34_/a_129_47# net10 0.003f
C171 VGND _27_/a_205_297# -3.36e-19
C172 net3 p[10] 3.61e-19
C173 net7 net17 0.2f
C174 _34_/a_47_47# _02_ 1.09e-19
C175 _05_ _02_ 0.00163f
C176 net2 b[3] 0.00395f
C177 VGND _39_/a_47_47# 0.0665f
C178 net17 _31_/a_35_297# 0.0514f
C179 _05_ _34_/a_47_47# 1.26e-20
C180 p[13] _44_/a_250_297# 4.09e-20
C181 p[1] _04_ 2.46e-21
C182 input5/a_381_47# b[1] 0.0023f
C183 _52_/a_93_21# b[1] 2.82e-19
C184 _42_/a_209_311# _02_ 9.92e-19
C185 net18 _06_ 0.0211f
C186 _13_ _15_ 3.69e-20
C187 input15/a_27_47# p[14] 7.31e-19
C188 _20_ _32_/a_303_47# 1.54e-19
C189 input5/a_664_47# _02_ 0.00187f
C190 net12 _21_ 0.23f
C191 net3 VGND 0.323f
C192 b[2] b[1] 5.48e-19
C193 p[7] net1 7.5e-20
C194 net5 _29_/a_29_53# 8.1e-20
C195 _38_/a_27_47# _25_ 5.76e-19
C196 input5/a_62_47# net2 0.0197f
C197 p[11] p[9] 0.00566f
C198 _35_/a_226_297# net10 2.48e-19
C199 net13 net4 2.48e-19
C200 _53_/a_29_53# b[1] 4.99e-19
C201 net1 net7 0.0712f
C202 _23_ _39_/a_285_47# 1.9e-20
C203 net1 _31_/a_35_297# 0.0111f
C204 _17_ _50_/a_223_47# 5.24e-20
C205 net8 VPWR 0.701f
C206 p[8] VPWR 0.151f
C207 _16_ net6 1.62e-20
C208 _43_/a_193_413# p[9] 1.09e-19
C209 input5/a_664_47# _42_/a_209_311# 0.0124f
C210 p[13] input14/a_27_47# 3.88e-19
C211 _18_ _43_/a_27_47# 0.0201f
C212 _13_ _45_/a_465_47# 0.00134f
C213 _39_/a_47_47# p[12] 3.32e-19
C214 _35_/a_489_413# _06_ 9.22e-19
C215 _33_/a_296_53# _06_ 1.11e-20
C216 _16_ _55_/a_472_297# 3.71e-19
C217 _55_/a_80_21# _02_ 0.164f
C218 _11_ _39_/a_377_297# 2.57e-20
C219 _01_ _49_/a_75_199# 0.009f
C220 _33_/a_368_53# net10 0.00171f
C221 _15_ _00_ 0.207f
C222 input15/a_27_47# VPWR 0.0113f
C223 p[11] _14_ 5.39e-21
C224 net12 _29_/a_29_53# 0.0132f
C225 net1 _47_/a_81_21# 1.58e-21
C226 net6 _47_/a_81_21# 2.14e-19
C227 net5 _30_/a_215_297# 8.27e-21
C228 _50_/a_27_47# _50_/a_223_47# 2.84e-32
C229 net8 net11 1.5e-19
C230 net14 _11_ 5e-19
C231 net10 _02_ 6.74e-19
C232 VGND input5/a_841_47# 0.0942f
C233 _55_/a_300_47# _22_ 2.08e-19
C234 _20_ _09_ 7.11e-19
C235 _43_/a_193_413# _14_ 0.0297f
C236 _42_/a_109_93# VPWR -0.00118f
C237 _26_/a_29_53# net4 0.00412f
C238 _24_ _21_ 0.0388f
C239 _38_/a_27_47# output18/a_27_47# 8.6e-19
C240 input6/a_27_47# p[9] 0.0756f
C241 net10 _34_/a_47_47# 0.0507f
C242 _42_/a_209_311# _55_/a_80_21# 0.0175f
C243 _10_ _39_/a_129_47# 2.51e-19
C244 VGND _17_ 0.312f
C245 _09_ b[1] 0.00408f
C246 _31_/a_285_297# VPWR 0.013f
C247 _49_/a_544_297# net13 3.43e-19
C248 _50_/a_343_93# net14 1.07e-20
C249 _44_/a_93_21# b[3] 7.01e-20
C250 _05_ net10 0.457f
C251 net14 _37_/a_303_47# 0.00112f
C252 _18_ VPWR 0.0721f
C253 _44_/a_250_297# _14_ 4.82e-19
C254 p[11] net19 0.00645f
C255 _44_/a_346_47# _14_ 3.76e-19
C256 input5/a_558_47# _06_ 3.55e-19
C257 _49_/a_201_297# _09_ 1.74e-20
C258 input14/a_27_47# p[9] 8.53e-21
C259 _45_/a_193_297# VPWR -0.00859f
C260 input5/a_62_47# _44_/a_93_21# 5.05e-20
C261 net12 _30_/a_215_297# 0.00676f
C262 VGND _50_/a_27_47# -0.00433f
C263 _43_/a_193_413# net19 3.31e-19
C264 input6/a_27_47# _14_ 3.75e-21
C265 _27_/a_277_297# _04_ 0.00113f
C266 _37_/a_27_47# net15 0.0541f
C267 _48_/a_181_47# VPWR -3.35e-19
C268 input3/a_27_47# net19 0.00105f
C269 net15 output19/a_27_47# 6.88e-19
C270 net14 _02_ 0.00952f
C271 p[7] b[1] 0.00406f
C272 _20_ net7 0.0257f
C273 net3 _29_/a_183_297# 7.38e-21
C274 net7 b[1] 0.0783f
C275 _20_ _31_/a_35_297# 1.69e-19
C276 _35_/a_76_199# _08_ 0.0061f
C277 _16_ _20_ 0.00271f
C278 _44_/a_346_47# net19 0.00124f
C279 net4 _14_ 1.54e-20
C280 _44_/a_250_297# net19 0.00592f
C281 _16_ b[1] 2.21e-19
C282 _31_/a_35_297# b[1] 0.0176f
C283 net9 _08_ 7.71e-21
C284 net9 _30_/a_109_53# 0.0191f
C285 _12_ net6 0.0891f
C286 input2/a_27_47# net7 0.00213f
C287 net3 _42_/a_296_53# 1.81e-19
C288 net14 _42_/a_209_311# 0.0238f
C289 _55_/a_217_297# _14_ 0.0116f
C290 input6/a_27_47# net19 0.00586f
C291 _04_ input8/a_27_47# 2.36e-22
C292 net14 input5/a_664_47# 0.0179f
C293 _49_/a_201_297# net7 0.00419f
C294 _35_/a_226_297# _03_ 0.00101f
C295 _40_/a_191_297# net6 1.16e-20
C296 net6 _40_/a_297_297# 7.47e-22
C297 input2/a_27_47# _31_/a_35_297# 0.00136f
C298 VGND p[2] 0.137f
C299 _48_/a_27_47# p[6] 2.33e-19
C300 _20_ _47_/a_81_21# 0.0457f
C301 net16 net6 8.27e-20
C302 output19/a_27_47# _10_ 3.23e-20
C303 _50_/a_27_47# p[12] 1.34e-19
C304 _49_/a_201_297# _31_/a_35_297# 5.52e-20
C305 net17 _04_ 0.0218f
C306 _48_/a_109_47# VGND 9.44e-19
C307 _50_/a_515_93# _10_ 0.00129f
C308 _11_ _50_/a_223_47# 0.0329f
C309 net13 VPWR 0.599f
C310 net4 net19 2.65e-20
C311 net1 _22_ 0.0129f
C312 _21_ net4 0.00535f
C313 net6 _22_ 0.163f
C314 _53_/a_111_297# VGND -2.89e-19
C315 _31_/a_117_297# VPWR 5.04e-19
C316 net19 input14/a_27_47# 3.63e-19
C317 _27_/a_27_297# _19_ 0.082f
C318 p[13] VPWR 0.197f
C319 _34_/a_129_47# VGND -8.76e-20
C320 _36_/a_303_47# _06_ 5.3e-19
C321 _45_/a_465_47# _09_ 2.77e-19
C322 net8 _27_/a_277_297# 7.99e-20
C323 net14 _55_/a_80_21# 4.7e-19
C324 _39_/a_47_47# _06_ 1.44e-19
C325 p[14] p[9] 0.355f
C326 _35_/a_226_47# _49_/a_75_199# 8.73e-20
C327 net6 _04_ 2.61e-20
C328 net1 _04_ 0.018f
C329 _34_/a_285_47# _02_ 7.14e-19
C330 _03_ _02_ 0.00474f
C331 net13 net11 0.0927f
C332 _26_/a_183_297# _14_ 6.98e-22
C333 net7 _15_ 8.4e-20
C334 VGND _11_ 0.0908f
C335 _03_ _34_/a_47_47# 4.5e-20
C336 VGND _35_/a_226_297# -4.55e-19
C337 net12 net5 0.0674f
C338 net3 _06_ 0.0072f
C339 _30_/a_109_53# _00_ 3.67e-20
C340 _05_ _03_ 0.135f
C341 _16_ _15_ 0.0607f
C342 _50_/a_223_47# _02_ 2.51e-20
C343 _34_/a_285_47# _05_ 7.85e-21
C344 _50_/a_343_93# VGND -4.3e-19
C345 _26_/a_29_53# VPWR 0.0356f
C346 VGND _37_/a_303_47# -1.63e-19
C347 _43_/a_27_47# _14_ 0.00938f
C348 net3 _47_/a_299_297# 2.55e-19
C349 _14_ p[14] 1.66e-20
C350 net8 input8/a_27_47# 0.0181f
C351 _15_ _47_/a_81_21# 0.00332f
C352 net10 p[5] 0.00544f
C353 net2 _37_/a_197_47# 4.74e-20
C354 p[0] p[10] 6.95e-20
C355 _19_ input7/a_27_47# 3.12e-21
C356 net8 net17 0.18f
C357 _33_/a_368_53# VGND 2.38e-19
C358 _12_ _20_ 3.9e-19
C359 VPWR p[9] 0.355f
C360 net16 _54_/a_75_212# 1.69e-21
C361 _20_ _40_/a_297_297# 9.18e-21
C362 _05_ p[10] 6e-20
C363 _26_/a_29_53# net11 1.08e-20
C364 _35_/a_76_199# _52_/a_250_297# 3.4e-21
C365 _12_ b[1] 3.18e-21
C366 _20_ _40_/a_191_297# 2.07e-20
C367 b[0] _39_/a_129_47# 2.6e-20
C368 VGND _02_ 1.63f
C369 _11_ p[12] 4.25e-21
C370 p[0] VGND 0.132f
C371 _42_/a_209_311# p[10] 2.37e-20
C372 net19 p[14] 0.101f
C373 _36_/a_27_47# _23_ 0.00118f
C374 VGND _34_/a_47_47# 0.0892f
C375 _20_ _22_ 0.183f
C376 _33_/a_209_311# _35_/a_489_413# 2.77e-20
C377 _01_ _27_/a_27_297# 8.04e-19
C378 input5/a_841_47# _06_ 1.66e-19
C379 VGND _05_ 0.754f
C380 net2 _40_/a_109_297# 0.0011f
C381 _22_ b[1] 9.74e-20
C382 net13 p[4] 2.34e-20
C383 net5 _24_ 5.83e-20
C384 _17_ _06_ 0.0341f
C385 _31_/a_285_297# input8/a_27_47# 1.04e-19
C386 net17 _42_/a_109_93# 3.1e-21
C387 net1 net8 0.381f
C388 _27_/a_27_297# net2 0.0131f
C389 _14_ VPWR 0.186f
C390 VGND _42_/a_209_311# -0.008f
C391 _10_ _07_ 2.19e-19
C392 _13_ _52_/a_250_297# 5.43e-19
C393 _53_/a_183_297# _02_ 4.14e-19
C394 VGND input5/a_664_47# 0.0134f
C395 net10 _03_ 0.321f
C396 _10_ _43_/a_369_47# 0.00199f
C397 _35_/a_76_199# _01_ 3.08e-21
C398 _33_/a_109_93# _02_ 1.54e-21
C399 _34_/a_285_47# net10 0.0454f
C400 _20_ _04_ 0.0677f
C401 _44_/a_584_47# net2 0.0053f
C402 _44_/a_256_47# VPWR -7.56e-19
C403 _49_/a_201_297# _22_ 2.45e-20
C404 _04_ b[1] 0.0568f
C405 _41_/a_59_75# _00_ 2.43e-20
C406 input15/a_27_47# net6 0.146f
C407 _33_/a_109_93# _05_ 0.0206f
C408 _01_ net9 0.157f
C409 _50_/a_27_47# _06_ 0.0097f
C410 net5 _43_/a_193_413# 1.39e-20
C411 net2 net9 3.64e-20
C412 _34_/a_377_297# _07_ 5.8e-19
C413 _23_ net9 1.21e-19
C414 _09_ _08_ 0.106f
C415 _21_ VPWR 0.869f
C416 net19 VPWR 0.186f
C417 input2/a_27_47# _04_ 4.5e-21
C418 _23_ _45_/a_27_47# 1.74e-19
C419 _30_/a_392_297# net10 3.4e-19
C420 _49_/a_201_297# _04_ 0.0253f
C421 _12_ _15_ 0.00833f
C422 net1 _31_/a_285_297# 5.85e-19
C423 VGND _55_/a_80_21# 0.00281f
C424 net5 _44_/a_250_297# 3.11e-20
C425 net2 input7/a_27_47# 3.24e-19
C426 _18_ net6 0.166f
C427 _13_ _23_ 2.08e-20
C428 net14 _03_ 1.5e-19
C429 _45_/a_193_297# net6 9.84e-20
C430 VGND net10 0.446f
C431 _15_ _22_ 0.0236f
C432 _21_ net11 0.586f
C433 net14 _50_/a_223_47# 5.89e-21
C434 _36_/a_27_47# _25_ 2.34e-20
C435 _52_/a_93_21# _52_/a_250_297# -6.97e-22
C436 _45_/a_465_47# _12_ 0.00211f
C437 _29_/a_29_53# VPWR 0.0299f
C438 net7 _08_ 9.54e-25
C439 _48_/a_109_47# _06_ 9.47e-19
C440 _38_/a_27_47# _10_ 0.0133f
C441 _31_/a_35_297# _30_/a_109_53# 2.89e-20
C442 b[2] _52_/a_250_297# 1.6e-19
C443 _35_/a_489_413# _07_ 0.00429f
C444 _15_ _04_ 3.61e-20
C445 _47_/a_384_47# _10_ 3.53e-19
C446 _53_/a_111_297# _06_ 3.82e-19
C447 net5 net4 0.0447f
C448 net8 _20_ 5.07e-19
C449 net13 net17 5.21e-20
C450 net14 p[10] 1.59e-20
C451 _32_/a_27_47# _11_ 1.65e-20
C452 _34_/a_129_47# _06_ 5.3e-19
C453 _33_/a_109_93# net10 0.0336f
C454 _01_ _00_ 0.00124f
C455 VGND _39_/a_377_297# -6.28e-19
C456 net17 _31_/a_117_297# 0.00149f
C457 net8 b[1] 0.0729f
C458 _19_ _09_ 4.8e-21
C459 net2 _00_ 0.00732f
C460 input9/a_75_212# p[3] 0.016f
C461 net5 _55_/a_217_297# 8.84e-20
C462 input4/a_75_212# _10_ 0.00372f
C463 _32_/a_27_47# _50_/a_343_93# 6.48e-20
C464 _17_ _39_/a_129_47# 1.38e-20
C465 _32_/a_109_47# _02_ 3.98e-19
C466 input2/a_27_47# net8 0.0207f
C467 net15 b[3] 0.00302f
C468 input13/a_27_47# _05_ 3.93e-19
C469 _48_/a_27_47# _53_/a_29_53# 3.14e-21
C470 _29_/a_29_53# net11 0.00514f
C471 net14 VGND 0.441f
C472 _37_/a_27_47# net3 0.094f
C473 net3 output19/a_27_47# 0.00348f
C474 _49_/a_201_297# net8 7.3e-19
C475 _11_ _06_ 0.493f
C476 input5/a_381_47# net2 0.0138f
C477 _01_ _32_/a_303_47# 8.58e-19
C478 _35_/a_226_297# _06_ 1.28e-19
C479 _35_/a_556_47# net10 5.59e-19
C480 _23_ _52_/a_93_21# 0.0166f
C481 _38_/a_27_47# net18 0.00997f
C482 net13 net1 3.51e-19
C483 net12 net4 2.57e-20
C484 _30_/a_215_297# VPWR -0.00548f
C485 net13 net6 0.00188f
C486 _23_ b[2] 2.87e-20
C487 _50_/a_343_93# _06_ 0.0376f
C488 _42_/a_109_93# b[1] 2.38e-19
C489 VGND p[5] 0.115f
C490 _55_/a_300_47# _14_ 8.09e-19
C491 p[13] net1 2.13e-19
C492 _47_/a_299_297# _11_ 0.00738f
C493 _31_/a_285_297# b[1] 0.0101f
C494 input11/a_27_47# VPWR 0.0375f
C495 b[0] output16/a_27_47# 0.014f
C496 _10_ b[3] 6.63e-21
C497 _32_/a_27_47# _02_ 0.00247f
C498 _35_/a_76_199# _35_/a_226_47# -2.84e-32
C499 _09_ _52_/a_250_297# 1.97e-20
C500 _18_ _20_ 0.0151f
C501 net7 _19_ 0.0458f
C502 _50_/a_223_47# _03_ 1.41e-21
C503 _19_ _31_/a_35_297# 1.47e-19
C504 _33_/a_368_53# _06_ 1.7e-19
C505 _32_/a_27_47# _05_ 2.2e-20
C506 _30_/a_215_297# net11 1.04e-19
C507 net12 _29_/a_111_297# 1.21e-19
C508 _35_/a_226_47# net9 1.22e-20
C509 _42_/a_368_53# net19 5.12e-19
C510 input3/a_27_47# p[11] 0.0137f
C511 _30_/a_392_297# _03_ 6.33e-19
C512 _48_/a_27_47# _09_ 0.00541f
C513 net8 _15_ 1.79e-19
C514 _35_/a_226_47# _45_/a_27_47# 5.71e-21
C515 p[10] _03_ 8.74e-20
C516 _06_ _02_ 0.85f
C517 net11 input11/a_27_47# 0.00318f
C518 _43_/a_297_47# _14_ 9.11e-19
C519 _37_/a_27_47# input5/a_841_47# 4.64e-20
C520 _26_/a_29_53# net6 0.0032f
C521 _48_/a_181_47# b[1] 3.46e-19
C522 net15 _49_/a_75_199# 5.13e-20
C523 _06_ _34_/a_47_47# 0.0391f
C524 _37_/a_27_47# _17_ 0.00277f
C525 _10_ _39_/a_285_47# 0.00289f
C526 output19/a_27_47# _17_ 0.00122f
C527 _31_/a_285_47# VPWR -2.91e-19
C528 _21_ input12/a_27_47# 2.32e-19
C529 _05_ _06_ 0.00724f
C530 _50_/a_429_93# net14 6.04e-21
C531 _44_/a_93_21# _00_ 4.54e-20
C532 _13_ _35_/a_226_47# 5.62e-21
C533 input13/a_27_47# net10 8.86e-20
C534 _01_ _09_ 4.69e-21
C535 input15/a_27_47# _15_ 2.15e-20
C536 VGND _03_ 0.119f
C537 _34_/a_285_47# VGND -0.00301f
C538 _24_ net4 8.65e-20
C539 _47_/a_81_21# _41_/a_59_75# 1.5e-19
C540 input3/a_27_47# _44_/a_250_297# 2.07e-19
C541 _42_/a_209_311# _06_ 1.66e-19
C542 net17 _14_ 2.4e-20
C543 _23_ _09_ 0.207f
C544 net6 p[9] 0.14f
C545 input5/a_664_47# _06_ 3.21e-19
C546 VGND _50_/a_223_47# 0.0159f
C547 _15_ _42_/a_109_93# 0.00367f
C548 _28_/a_109_297# VPWR -1.71e-19
C549 _22_ _30_/a_109_53# 3.67e-21
C550 p[11] input14/a_27_47# 3.98e-20
C551 _30_/a_392_297# VGND 3.41e-19
C552 net13 _20_ 5.95e-19
C553 _25_ b[2] 0.0015f
C554 _33_/a_109_93# _03_ 2.78e-19
C555 VGND p[10] 0.177f
C556 net13 b[1] 0.0495f
C557 net5 VPWR 0.613f
C558 _18_ _15_ 0.042f
C559 net17 net19 8.84e-23
C560 _32_/a_27_47# net10 2.76e-20
C561 _53_/a_29_53# _25_ 0.00146f
C562 net6 _14_ 2.11e-19
C563 _31_/a_117_297# b[1] 0.00281f
C564 _01_ net7 0.233f
C565 input3/a_27_47# input14/a_27_47# 5.08e-20
C566 _04_ _30_/a_109_53# 9.19e-21
C567 p[13] b[1] 0.00201f
C568 net9 _30_/a_297_297# 7.53e-19
C569 _55_/a_80_21# _06_ 5.15e-19
C570 net7 net2 0.00234f
C571 p[4] input11/a_27_47# 0.0646f
C572 net14 _42_/a_296_53# 2.18e-19
C573 _01_ _31_/a_35_297# 4.27e-19
C574 _04_ _08_ 5.99e-19
C575 _16_ _01_ 3.24e-19
C576 net13 _49_/a_201_297# 3.31e-19
C577 net3 _37_/a_109_47# 0.00212f
C578 _55_/a_472_297# _14_ 0.00192f
C579 net2 _31_/a_35_297# 0.0635f
C580 _35_/a_226_47# _52_/a_93_21# 4.89e-20
C581 _44_/a_250_297# input14/a_27_47# 8.25e-21
C582 _16_ net2 0.00654f
C583 net10 _06_ 0.184f
C584 _50_/a_615_93# _10_ 8.82e-19
C585 net5 net11 0.0129f
C586 input13/a_27_47# p[5] 3.09e-19
C587 _27_/a_27_297# _27_/a_109_297# -3.68e-20
C588 _10_ p[3] 1.37e-20
C589 _21_ net1 0.0252f
C590 net12 VPWR 0.82f
C591 _26_/a_29_53# _20_ 0.00447f
C592 _01_ _47_/a_81_21# 6.05e-21
C593 _21_ net6 2.92e-20
C594 net6 net19 0.00352f
C595 _53_/a_183_297# VGND -4.34e-19
C596 output18/a_27_47# b[2] 0.0141f
C597 _26_/a_29_53# b[1] 9.93e-21
C598 _12_ _41_/a_59_75# 0.00101f
C599 net2 _47_/a_81_21# 4.95e-19
C600 _33_/a_109_93# VGND -0.0132f
C601 _25_ _09_ 1.49e-19
C602 _53_/a_29_53# output18/a_27_47# 9.46e-19
C603 input9/a_75_212# net9 0.0245f
C604 _39_/a_377_297# _06_ 8.76e-20
C605 net5 _45_/a_205_47# 8.28e-20
C606 net4 _55_/a_217_297# 1.13e-19
C607 VGND p[12] 0.36f
C608 net12 net11 0.356f
C609 _22_ _41_/a_59_75# 6.24e-22
C610 _45_/a_109_297# _35_/a_226_47# 1.59e-21
C611 _37_/a_27_47# _11_ 0.0018f
C612 _29_/a_183_297# _03_ 7.36e-19
C613 VGND _35_/a_556_47# 1.95e-19
C614 _17_ _37_/a_109_47# 8.86e-21
C615 net14 _06_ 1.94e-19
C616 _04_ _19_ 0.356f
C617 _17_ _43_/a_369_47# 5.87e-19
C618 _12_ _52_/a_250_297# 0.0139f
C619 _29_/a_29_53# net1 9.76e-19
C620 _29_/a_29_53# net6 1.4e-20
C621 _50_/a_429_93# VGND 4.71e-19
C622 _26_/a_111_297# VPWR -5.92e-20
C623 net8 _30_/a_109_53# 1.76e-20
C624 _35_/a_226_47# _09_ 0.0599f
C625 _30_/a_215_297# net17 4.69e-20
C626 _20_ _14_ 0.144f
C627 _24_ VPWR 0.0129f
C628 input4/a_75_212# _39_/a_47_47# 3.1e-19
C629 _22_ _52_/a_250_297# 0.0996f
C630 _14_ b[1] 1.1e-19
C631 _16_ _44_/a_93_21# 0.00354f
C632 input5/a_62_47# output17/a_27_47# 1.02e-19
C633 _26_/a_29_53# _15_ 0.00192f
C634 _49_/a_208_47# _09_ 5.43e-21
C635 net15 _37_/a_197_47# 1.78e-19
C636 net15 _43_/a_469_47# 7.41e-19
C637 b[0] _39_/a_285_47# 1.88e-19
C638 p[11] VPWR 0.197f
C639 input6/a_27_47# p[14] 0.0157f
C640 _49_/a_201_297# _14_ 4.76e-21
C641 _34_/a_377_297# p[6] 5.39e-19
C642 _32_/a_27_47# _03_ 1.9e-19
C643 _04_ _52_/a_250_297# 3.98e-21
C644 _12_ net2 1.02e-20
C645 _12_ _23_ 0.00743f
C646 _30_/a_215_297# net1 0.00375f
C647 VGND _29_/a_183_297# 4.41e-19
C648 _21_ _20_ 0.191f
C649 _36_/a_109_47# _23_ 3.44e-19
C650 _30_/a_215_297# net6 3.3e-21
C651 net2 _40_/a_191_297# 0.00143f
C652 _43_/a_193_413# VPWR 0.0063f
C653 net2 _40_/a_297_297# 0.00101f
C654 _20_ net19 1.29e-19
C655 output17/a_27_47# input1/a_75_212# 0.0101f
C656 net19 b[1] 1e-19
C657 input13/a_27_47# VGND 0.0471f
C658 net12 p[4] 5.33e-19
C659 _21_ b[1] 0.00892f
C660 p[7] _35_/a_226_47# 2.82e-19
C661 _15_ p[9] 2.06e-19
C662 _01_ _22_ 0.15f
C663 input3/a_27_47# VPWR 0.0688f
C664 _35_/a_226_47# net7 2.93e-20
C665 net15 _40_/a_109_297# 0.0016f
C666 _37_/a_27_47# _42_/a_209_311# 1.59e-20
C667 net17 _31_/a_285_47# 0.00134f
C668 VGND _32_/a_109_47# 1.05e-19
C669 net2 _22_ 1.93e-20
C670 input2/a_27_47# net19 2.9e-23
C671 net15 _27_/a_27_297# 0.00888f
C672 _06_ _03_ 0.00635f
C673 net3 b[3] 2.43e-20
C674 _44_/a_346_47# VPWR -8.74e-19
C675 _10_ _43_/a_469_47# 0.00124f
C676 _23_ _22_ 0.0187f
C677 _34_/a_285_47# _06_ 0.00598f
C678 _43_/a_27_47# _55_/a_217_297# 2.18e-19
C679 _44_/a_250_297# VPWR 0.0233f
C680 _47_/a_384_47# _17_ 1.1e-20
C681 net8 _19_ 0.0322f
C682 _33_/a_209_311# _34_/a_47_47# 0.017f
C683 _48_/a_109_47# _07_ 3.01e-19
C684 _49_/a_208_47# net7 0.00312f
C685 _01_ _04_ 0.119f
C686 _33_/a_209_311# _05_ 0.0311f
C687 _50_/a_223_47# _06_ 0.0464f
C688 input6/a_27_47# VPWR 0.00162f
C689 _33_/a_109_93# input13/a_27_47# 0.00348f
C690 _15_ _14_ 0.148f
C691 net2 _04_ 0.158f
C692 net3 input5/a_62_47# 0.00164f
C693 _30_/a_465_297# net10 0.00106f
C694 _36_/a_27_47# _10_ 0.00109f
C695 _29_/a_29_53# _20_ 0.0111f
C696 _38_/a_27_47# _50_/a_27_47# 2.37e-20
C697 _29_/a_29_53# b[1] 0.0026f
C698 _32_/a_27_47# VGND 0.0233f
C699 _47_/a_299_297# _50_/a_223_47# 2.74e-20
C700 net15 net9 8.49e-20
C701 net12 input12/a_27_47# 0.0297f
C702 net4 VPWR 1.07f
C703 input15/a_27_47# _41_/a_59_75# 3.96e-20
C704 net5 net17 4.21e-21
C705 VPWR input14/a_27_47# 0.0739f
C706 _19_ _42_/a_109_93# 1.14e-21
C707 _31_/a_285_297# _19_ 1.34e-19
C708 _55_/a_217_297# VPWR -0.00133f
C709 _44_/a_584_47# _10_ 1.14e-20
C710 _21_ _15_ 1.13e-21
C711 _15_ net19 0.166f
C712 VGND _06_ 1.09f
C713 net15 input7/a_27_47# 1.88e-19
C714 _35_/a_76_199# _10_ 7.19e-20
C715 net13 _30_/a_109_53# 1.05e-19
C716 _12_ _25_ 1.23e-20
C717 _52_/a_93_21# _52_/a_256_47# -6.6e-20
C718 _17_ b[3] 7.54e-20
C719 net3 _49_/a_75_199# 2.01e-19
C720 _36_/a_109_47# _25_ 3.76e-21
C721 net13 _08_ 1.82e-19
C722 _10_ net9 0.0438f
C723 _30_/a_215_297# _20_ 6.08e-19
C724 _29_/a_111_297# VPWR -5.85e-19
C725 net16 _25_ 1.16e-19
C726 VGND _47_/a_299_297# -3.63e-19
C727 _38_/a_109_47# _10_ 5.44e-19
C728 net5 net6 0.727f
C729 _45_/a_27_47# _10_ 0.0143f
C730 _30_/a_215_297# b[1] 0.0176f
C731 net5 net1 0.0772f
C732 _12_ _38_/a_197_47# 0.00173f
C733 _53_/a_183_297# _06_ 0.00146f
C734 net12 net17 2.11e-21
C735 _33_/a_109_93# _06_ 6.96e-19
C736 _33_/a_209_311# net10 0.0426f
C737 _25_ _22_ 5.39e-19
C738 _49_/a_544_297# VPWR 0.00504f
C739 _13_ _10_ 0.0621f
C740 net16 _38_/a_197_47# 5.89e-19
C741 input2/a_27_47# _30_/a_215_297# 3.51e-20
C742 input11/a_27_47# b[1] 0.00688f
C743 _01_ net8 0.0802f
C744 _17_ _39_/a_285_47# 7.36e-21
C745 _32_/a_197_47# _02_ 3.78e-19
C746 _07_ _02_ 0.0083f
C747 _49_/a_315_47# _09_ 1.11e-20
C748 net8 net2 0.0525f
C749 _29_/a_111_297# net11 8.27e-19
C750 p[8] net2 0.0177f
C751 _37_/a_27_47# net14 0.0584f
C752 net15 _00_ 0.00147f
C753 _12_ _35_/a_226_47# 8.38e-20
C754 _06_ p[12] 0.0535f
C755 _44_/a_93_21# _04_ 4.47e-21
C756 _07_ _34_/a_47_47# 0.011f
C757 _26_/a_183_297# VPWR -3.03e-19
C758 net14 output19/a_27_47# 0.00142f
C759 p[7] input9/a_75_212# 0.00102f
C760 _05_ _07_ 1.21e-19
C761 _18_ _52_/a_250_297# 1.77e-19
C762 net14 _50_/a_515_93# 1.39e-20
C763 net12 net6 0.00643f
C764 net12 net1 1.17e-19
C765 net15 input5/a_381_47# 7.15e-19
C766 _50_/a_429_93# _06_ 0.00169f
C767 _11_ _38_/a_27_47# 0.071f
C768 net2 input15/a_27_47# 0.00296f
C769 _47_/a_299_297# p[12] 8.13e-21
C770 _35_/a_226_47# _22_ 1.39e-20
C771 _43_/a_27_47# VPWR 0.0186f
C772 _47_/a_384_47# _11_ 7.23e-20
C773 net16 output18/a_27_47# 3.45e-19
C774 VPWR p[14] 0.0354f
C775 _31_/a_285_47# b[1] 8.76e-19
C776 net13 _19_ 4.45e-20
C777 _01_ _31_/a_285_297# 1.92e-19
C778 net2 _42_/a_109_93# 0.00507f
C779 output18/a_27_47# _22_ 7.51e-19
C780 _10_ _00_ 0.301f
C781 _49_/a_315_47# net7 0.00706f
C782 _18_ _01_ 6.1e-20
C783 _35_/a_226_47# _04_ 0.00551f
C784 _20_ _28_/a_109_297# 0.00221f
C785 _30_/a_465_297# _03_ 7.72e-19
C786 _35_/a_489_413# _45_/a_27_47# 3.89e-21
C787 _18_ net2 0.00181f
C788 _10_ _52_/a_93_21# 0.00534f
C789 _26_/a_111_297# net6 1.12e-19
C790 VGND _39_/a_129_47# -0.00126f
C791 _45_/a_193_297# _23_ 4.13e-19
C792 input5/a_558_47# _27_/a_27_297# 1.57e-19
C793 _38_/a_27_47# _02_ 0.00103f
C794 net5 _20_ 0.0651f
C795 input13/a_27_47# _06_ 4.89e-19
C796 net5 b[1] 0.00349f
C797 _24_ net6 0.00121f
C798 _07_ net10 0.0605f
C799 _53_/a_29_53# _10_ 0.00779f
C800 input5/a_558_47# net9 4.42e-19
C801 net18 _52_/a_93_21# 8.21e-21
C802 _21_ _30_/a_109_53# 3.31e-20
C803 p[2] _49_/a_75_199# 1.1e-19
C804 _21_ _08_ 0.00139f
C805 net18 b[2] 0.0131f
C806 net12 _20_ 0.00437f
C807 _30_/a_465_297# VGND 6.42e-19
C808 _43_/a_193_413# net6 2.41e-20
C809 net11 VPWR 0.994f
C810 _45_/a_109_297# _10_ 0.00202f
C811 _33_/a_209_311# _03_ 8.38e-19
C812 net12 b[1] 0.12f
C813 p[9] _41_/a_59_75# 1.02e-19
C814 _32_/a_27_47# _06_ 0.00663f
C815 net13 _01_ 0.00228f
C816 _44_/a_93_21# _42_/a_109_93# 1.25e-19
C817 _53_/a_29_53# net18 0.0118f
C818 p[1] VPWR 0.0793f
C819 input5/a_558_47# input7/a_27_47# 1.22e-20
C820 _28_/a_109_297# _15_ 0.00346f
C821 _52_/a_346_47# _02_ 0.00526f
C822 net13 _23_ 4.11e-19
C823 _10_ _09_ 0.0222f
C824 p[13] _01_ 2.02e-20
C825 net3 _37_/a_197_47# 0.0028f
C826 net14 _37_/a_109_47# 1.71e-19
C827 _37_/a_27_47# VGND -0.0147f
C828 net14 _43_/a_369_47# 6.79e-21
C829 VGND output19/a_27_47# -0.00902f
C830 p[13] net2 0.0246f
C831 _18_ _44_/a_93_21# 0.00485f
C832 _19_ _14_ 2.71e-21
C833 _45_/a_205_47# VPWR -1.62e-19
C834 net15 net7 2.91e-19
C835 _50_/a_515_93# VGND -4.75e-19
C836 net5 _15_ 0.0352f
C837 input6/a_27_47# net6 0.00208f
C838 _49_/a_208_47# net8 1.4e-19
C839 _29_/a_29_53# _30_/a_109_53# 0.0103f
C840 _16_ net15 0.214f
C841 p[2] p[3] 0.0526f
C842 _13_ b[0] 0.00299f
C843 input10/a_27_47# input11/a_27_47# 5.3e-19
C844 _47_/a_299_297# _06_ 0.0174f
C845 p[0] input5/a_62_47# 1.39e-19
C846 _33_/a_209_311# VGND -0.00749f
C847 net3 _40_/a_109_297# 3.14e-19
C848 _39_/a_285_47# _02_ 0.0019f
C849 net4 net6 0.713f
C850 net18 _09_ 1.97e-21
C851 net3 _27_/a_27_297# 0.0166f
C852 net15 _47_/a_81_21# 0.00106f
C853 p[4] VPWR 0.112f
C854 input9/a_75_212# _04_ 7.69e-22
C855 _24_ b[1] 2.68e-19
C856 net7 _10_ 6.22e-20
C857 _16_ _10_ 0.00486f
C858 output19/a_27_47# p[12] 1.78e-19
C859 _27_/a_109_297# _04_ 7.2e-20
C860 net19 _41_/a_59_75# 3.1e-20
C861 p[0] input1/a_75_212# 0.0177f
C862 _45_/a_193_297# _35_/a_226_47# 8.15e-21
C863 _45_/a_27_47# _39_/a_47_47# 1.31e-19
C864 _50_/a_515_93# p[12] 3.12e-21
C865 _17_ _43_/a_469_47# 0.00177f
C866 _17_ _37_/a_197_47# 9.19e-21
C867 p[11] b[1] 2.45e-20
C868 _42_/a_368_53# VPWR -3.03e-19
C869 net2 p[9] 0.00112f
C870 net3 net9 5.09e-20
C871 _49_/a_75_199# _02_ 0.0354f
C872 _43_/a_193_413# _20_ 0.00161f
C873 net8 _30_/a_297_297# 2.42e-21
C874 p[4] net11 0.0557f
C875 _49_/a_315_47# _04_ 7.71e-19
C876 _07_ _03_ 0.0113f
C877 _10_ _47_/a_81_21# 0.0061f
C878 _13_ _39_/a_47_47# 0.00117f
C879 _34_/a_285_47# _07_ 0.00975f
C880 _35_/a_489_413# _09_ 0.0296f
C881 net13 _25_ 0.00297f
C882 _55_/a_300_47# VPWR -4.61e-19
C883 input3/a_27_47# b[1] 2.97e-19
C884 input12/a_27_47# VPWR 0.0646f
C885 _49_/a_544_297# net1 0.00175f
C886 input5/a_381_47# output17/a_27_47# 6.6e-20
C887 _27_/a_277_297# VPWR -3.63e-19
C888 _01_ _14_ 0.0193f
C889 _17_ _40_/a_109_297# 9.67e-19
C890 net2 _14_ 0.0104f
C891 b[0] b[2] 0.183f
C892 VGND output16/a_27_47# 0.0728f
C893 _17_ _27_/a_27_297# 6.78e-22
C894 _48_/a_27_47# _21_ 0.0121f
C895 _43_/a_297_47# VPWR -2.11e-19
C896 _36_/a_27_47# _50_/a_27_47# 6.08e-19
C897 net13 _35_/a_226_47# 0.00709f
C898 net15 _12_ 8.14e-21
C899 _39_/a_47_47# _00_ 1.85e-20
C900 net11 input12/a_27_47# 0.00246f
C901 _01_ _21_ 7.94e-19
C902 _01_ net19 4.9e-19
C903 _43_/a_27_47# net6 9.07e-20
C904 net6 p[14] 0.00245f
C905 input8/a_27_47# VPWR 0.0863f
C906 input5/a_841_47# net9 2.7e-19
C907 VGND _32_/a_197_47# 8.12e-20
C908 VGND _07_ 0.195f
C909 VGND _37_/a_109_47# -7.9e-19
C910 net15 _40_/a_191_297# 8.41e-19
C911 net15 _40_/a_297_297# 4.08e-19
C912 VGND _43_/a_369_47# -8.43e-19
C913 _20_ net4 3.01e-20
C914 _05_ p[3] 8.47e-21
C915 _21_ _23_ 0.0217f
C916 _17_ net9 2.89e-23
C917 p[11] _15_ 0.00178f
C918 net2 net19 0.599f
C919 net17 VPWR 0.037f
C920 net3 _00_ 2.12e-19
C921 _17_ _45_/a_27_47# 1.16e-20
C922 net14 b[3] 9.2e-19
C923 p[1] _27_/a_277_297# 1.22e-21
C924 net15 _22_ 2.74e-19
C925 _20_ _55_/a_217_297# 0.0013f
C926 _43_/a_193_413# _15_ 4.86e-19
C927 _52_/a_93_21# _39_/a_47_47# 1.44e-20
C928 net12 input10/a_27_47# 0.00115f
C929 _33_/a_209_311# input13/a_27_47# 5.85e-20
C930 input3/a_27_47# _15_ 7.53e-19
C931 _12_ _10_ 0.19f
C932 net5 _30_/a_109_53# 5.84e-22
C933 _33_/a_109_93# _07_ 3.2e-19
C934 net14 input5/a_62_47# 5.28e-20
C935 net3 input5/a_381_47# 0.0299f
C936 _45_/a_27_47# _50_/a_27_47# 0.109f
C937 _44_/a_250_297# _15_ 0.00517f
C938 net16 _10_ 0.0338f
C939 net15 _04_ 0.0569f
C940 _29_/a_29_53# _01_ 8.33e-20
C941 net11 net17 3.19e-20
C942 net1 VPWR 1.17f
C943 net6 VPWR 0.999f
C944 input5/a_558_47# net7 0.00358f
C945 input6/a_27_47# _15_ 5.75e-19
C946 _44_/a_93_21# _14_ 0.04f
C947 _13_ _50_/a_27_47# 0.00169f
C948 _10_ _22_ 0.0904f
C949 p[1] input8/a_27_47# 5.13e-20
C950 p[1] net17 6.79e-20
C951 _49_/a_544_297# b[1] 8.23e-19
C952 _35_/a_556_47# _07_ 0.00128f
C953 _55_/a_472_297# VPWR 0.00488f
C954 _37_/a_27_47# _06_ 2.5e-20
C955 p[6] _34_/a_47_47# 4.27e-19
C956 p[4] input12/a_27_47# 8.26e-19
C957 _44_/a_256_47# _44_/a_93_21# -6.6e-20
C958 output19/a_27_47# _06_ 1.53e-19
C959 _12_ net18 8.24e-19
C960 net13 _30_/a_297_297# 3.27e-20
C961 net12 _30_/a_109_53# 4.25e-20
C962 net12 _08_ 0.0269f
C963 _50_/a_515_93# _06_ 0.00244f
C964 _17_ _00_ 0.0851f
C965 VGND _38_/a_27_47# 0.00766f
C966 _10_ _04_ 9.24e-20
C967 net10 p[3] 8.3e-19
C968 net14 _49_/a_75_199# 3.67e-19
C969 _15_ net4 0.00427f
C970 p[2] net9 1.4e-20
C971 net1 net11 1.13e-19
C972 VGND _47_/a_384_47# -2.05e-19
C973 net11 net6 1.08e-19
C974 net16 net18 0.00585f
C975 net7 output17/a_27_47# 0.0018f
C976 _11_ _40_/a_109_297# 0.00522f
C977 _12_ _38_/a_303_47# 0.00153f
C978 _39_/a_47_47# _09_ 7.7e-21
C979 _44_/a_93_21# net19 0.0074f
C980 _15_ _55_/a_217_297# 0.0474f
C981 _20_ _43_/a_27_47# 0.0124f
C982 net18 _22_ 1.68e-19
C983 _21_ _25_ 0.00164f
C984 p[1] net1 0.029f
C985 _33_/a_209_311# _06_ 0.0187f
C986 input4/a_75_212# VGND 0.0529f
C987 _50_/a_27_47# _00_ 0.00197f
C988 net16 _38_/a_303_47# 6.47e-19
C989 p[2] input7/a_27_47# 0.0023f
C990 _34_/a_377_297# _04_ 1.7e-20
C991 net5 _19_ 6.41e-21
C992 _45_/a_205_47# net6 2.59e-20
C993 _35_/a_76_199# _11_ 6.99e-22
C994 net5 _41_/a_59_75# 2.41e-19
C995 net15 net8 0.2f
C996 p[8] net15 1.73e-20
C997 net14 _50_/a_615_93# 1.69e-20
C998 net13 input9/a_75_212# 4.4e-19
C999 net13 _36_/a_197_47# 1.06e-19
C1000 VGND _52_/a_346_47# -0.00175f
C1001 _11_ net9 5.39e-19
C1002 _21_ _35_/a_226_47# 9.87e-19
C1003 _54_/a_75_212# VPWR 0.0475f
C1004 _36_/a_27_47# _02_ 9.37e-20
C1005 _11_ _45_/a_27_47# 0.0703f
C1006 _20_ VPWR 0.34f
C1007 VGND b[3] 0.127f
C1008 net10 p[6] 0.0023f
C1009 _27_/a_27_297# _02_ 0.00179f
C1010 VPWR b[1] 1.05f
C1011 _26_/a_183_297# _15_ 4.63e-36
C1012 _50_/a_343_93# net9 6.64e-19
C1013 net15 input15/a_27_47# 0.00325f
C1014 _01_ _31_/a_285_47# 3.36e-19
C1015 _36_/a_27_47# _05_ 3.67e-21
C1016 _45_/a_109_297# _17_ 4.29e-22
C1017 _21_ output18/a_27_47# 0.00103f
C1018 input4/a_75_212# p[12] 0.02f
C1019 net3 net7 7.45e-20
C1020 _03_ _49_/a_75_199# 0.0849f
C1021 net5 _52_/a_250_297# 0.018f
C1022 _13_ _11_ 0.164f
C1023 net8 _10_ 5.86e-19
C1024 input2/a_27_47# VPWR 0.00832f
C1025 net15 _42_/a_109_93# 4.62e-19
C1026 _16_ net3 1.77e-19
C1027 VGND input5/a_62_47# 0.0489f
C1028 _49_/a_201_297# VPWR 0.0175f
C1029 _50_/a_343_93# _13_ 5.63e-20
C1030 _27_/a_27_297# _42_/a_209_311# 4.7e-20
C1031 _54_/a_75_212# net11 0.00956f
C1032 _15_ _43_/a_27_47# 8.96e-20
C1033 _35_/a_76_199# _02_ 5.73e-19
C1034 _15_ p[14] 5.32e-19
C1035 _20_ net11 0.00128f
C1036 VGND _39_/a_285_47# -0.0046f
C1037 input5/a_664_47# _27_/a_27_297# 0.0116f
C1038 input15/a_27_47# _10_ 4.5e-19
C1039 net9 _02_ 0.00611f
C1040 net11 b[1] 0.0777f
C1041 _35_/a_76_199# _05_ 0.00238f
C1042 _38_/a_109_47# _02_ 1.63e-19
C1043 _29_/a_29_53# _35_/a_226_47# 2.64e-19
C1044 _18_ net15 0.0382f
C1045 net3 _47_/a_81_21# 6.66e-19
C1046 _45_/a_27_47# _02_ 0.00449f
C1047 VGND input1/a_75_212# 0.0581f
C1048 net9 _34_/a_47_47# 1.41e-20
C1049 b[3] p[12] 7.54e-20
C1050 net5 _01_ 0.0779f
C1051 _07_ _06_ 0.185f
C1052 _05_ net9 0.124f
C1053 _12_ b[0] 2.61e-20
C1054 net1 input12/a_27_47# 7.44e-20
C1055 _45_/a_27_47# _05_ 9.34e-23
C1056 _43_/a_369_47# _06_ -2.02e-19
C1057 _50_/a_27_47# _09_ 1.3e-19
C1058 p[1] b[1] 0.00409f
C1059 _49_/a_201_297# net11 1.42e-19
C1060 _11_ _00_ 0.238f
C1061 net5 _23_ 0.0052f
C1062 net5 net2 0.0616f
C1063 _13_ _02_ 0.0676f
C1064 p[3] _03_ 0.00347f
C1065 p[0] input7/a_27_47# 5.13e-20
C1066 VGND _49_/a_75_199# 5.87e-20
C1067 net12 _48_/a_27_47# 0.0126f
C1068 net16 b[0] 0.0306f
C1069 input2/a_27_47# p[1] 0.0118f
C1070 input5/a_558_47# _04_ 1.25e-20
C1071 input5/a_841_47# net7 0.00193f
C1072 input5/a_664_47# net9 5.29e-19
C1073 _50_/a_343_93# _00_ 0.102f
C1074 _13_ _05_ 2.57e-20
C1075 _18_ _10_ 0.133f
C1076 _15_ VPWR 0.912f
C1077 p[6] p[5] 0.0563f
C1078 _16_ input5/a_841_47# 8.62e-19
C1079 _45_/a_193_297# _10_ 0.0047f
C1080 _43_/a_297_47# net6 8.23e-22
C1081 _36_/a_27_47# net10 0.0364f
C1082 _16_ _17_ 0.242f
C1083 net12 _01_ 1.67e-21
C1084 input5/a_664_47# input7/a_27_47# 1.08e-21
C1085 net1 input8/a_27_47# 0.0347f
C1086 _52_/a_584_47# _02_ 0.00389f
C1087 net12 _23_ 2.28e-21
C1088 _43_/a_193_413# _19_ 4.85e-21
C1089 _53_/a_29_53# _11_ 2.33e-20
C1090 net1 net17 2.89e-19
C1091 net14 _43_/a_469_47# 1.44e-20
C1092 net14 _37_/a_197_47# 7e-19
C1093 p[4] b[1] 0.00668f
C1094 output17/a_27_47# _04_ 0.027f
C1095 _17_ _47_/a_81_21# 0.0456f
C1096 _02_ _00_ 0.0269f
C1097 _45_/a_465_47# VPWR -5.05e-19
C1098 net13 net15 8.84e-19
C1099 _35_/a_76_199# net10 0.0226f
C1100 _50_/a_615_93# VGND -5.19e-19
C1101 _12_ _39_/a_47_47# 0.0317f
C1102 _24_ _52_/a_250_297# 3.03e-19
C1103 VGND p[3] 0.17f
C1104 _53_/a_111_297# _09_ 3.4e-19
C1105 net16 _39_/a_47_47# 7.7e-20
C1106 p[13] net15 1.46e-19
C1107 input9/a_75_212# _21_ 1.17e-21
C1108 _05_ _00_ 5.03e-22
C1109 net9 net10 0.111f
C1110 net3 _12_ 3.09e-20
C1111 _52_/a_93_21# _02_ 0.0962f
C1112 _38_/a_27_47# _06_ 0.0172f
C1113 _42_/a_368_53# b[1] 5.32e-20
C1114 _34_/a_285_47# p[6] 8.62e-20
C1115 net3 _40_/a_191_297# 1.89e-19
C1116 net3 _40_/a_297_297# 2.54e-19
C1117 _45_/a_109_297# _11_ 0.00168f
C1118 b[2] _02_ 2.81e-19
C1119 net14 _27_/a_27_297# 0.0118f
C1120 net5 _44_/a_93_21# 3.61e-20
C1121 _32_/a_303_47# _02_ 1.15e-20
C1122 net13 _10_ 0.00151f
C1123 _05_ _52_/a_93_21# 1.12e-20
C1124 net5 _25_ 6.42e-19
C1125 _55_/a_300_47# b[1] 1.1e-19
C1126 net3 _22_ 9.39e-20
C1127 _13_ net10 4.52e-21
C1128 input4/a_75_212# _06_ 0.00205f
C1129 net7 p[2] 0.00156f
C1130 input5/a_558_47# net8 0.00357f
C1131 _53_/a_29_53# _02_ 0.0388f
C1132 _11_ _09_ 0.0665f
C1133 input12/a_27_47# b[1] 0.00658f
C1134 _27_/a_205_297# _04_ 6.42e-19
C1135 input5/a_381_47# _42_/a_209_311# 3.88e-19
C1136 _35_/a_226_297# _09_ 4.98e-19
C1137 net14 _44_/a_584_47# 7.2e-19
C1138 _26_/a_29_53# net15 9.06e-21
C1139 _27_/a_277_297# b[1] 1.24e-19
C1140 p[2] _31_/a_35_297# 0.00264f
C1141 _53_/a_29_53# _34_/a_47_47# 5.88e-22
C1142 _24_ _23_ 0.012f
C1143 _30_/a_215_297# _30_/a_297_297# -8.88e-34
C1144 _29_/a_29_53# input9/a_75_212# 9.7e-21
C1145 net4 _41_/a_59_75# 1.76e-19
C1146 net3 _04_ 0.113f
C1147 net14 net9 7.12e-20
C1148 input10/a_27_47# VPWR 0.00986f
C1149 _55_/a_80_21# _00_ 5.5e-19
C1150 _52_/a_346_47# _06_ 0.0031f
C1151 net15 p[9] 0.00295f
C1152 VGND p[6] 0.128f
C1153 net2 p[11] 0.00557f
C1154 _45_/a_109_297# _02_ 8.44e-19
C1155 input5/a_558_47# _42_/a_109_93# 1.75e-19
C1156 net8 output17/a_27_47# 0.0043f
C1157 net12 _25_ 4.46e-20
C1158 _43_/a_193_413# _01_ 8.16e-19
C1159 _12_ _17_ 0.0109f
C1160 _26_/a_29_53# _10_ 0.0265f
C1161 b[3] _06_ 9.96e-21
C1162 input8/a_27_47# b[1] 0.00172f
C1163 _45_/a_109_297# _05_ 2.79e-22
C1164 _43_/a_193_413# net2 1.52e-19
C1165 _17_ _40_/a_191_297# 4.35e-19
C1166 net14 input7/a_27_47# 3.48e-19
C1167 _20_ net17 4e-20
C1168 net17 b[1] 0.0287f
C1169 input3/a_27_47# net2 0.0229f
C1170 _09_ _02_ 0.297f
C1171 net4 _52_/a_250_297# 0.00136f
C1172 _16_ _11_ 4.42e-20
C1173 input10/a_27_47# net11 0.112f
C1174 _17_ _22_ 0.00334f
C1175 _49_/a_201_297# input8/a_27_47# 2.46e-21
C1176 _52_/a_93_21# net10 7.84e-20
C1177 _05_ _09_ 0.0683f
C1178 _44_/a_346_47# net2 1.64e-19
C1179 net15 _14_ 0.0538f
C1180 _55_/a_300_47# _15_ 1.42e-20
C1181 _10_ p[9] 0.00225f
C1182 _30_/a_215_297# input9/a_75_212# 6.24e-21
C1183 _27_/a_27_297# _03_ 2.68e-19
C1184 input2/a_27_47# net17 0.0398f
C1185 net2 _44_/a_250_297# 0.0188f
C1186 _12_ _50_/a_27_47# 0.00354f
C1187 _36_/a_27_47# _50_/a_223_47# 1.27e-20
C1188 _39_/a_285_47# _06_ 1.23e-20
C1189 output17/a_27_47# _42_/a_109_93# 8.6e-21
C1190 net13 _35_/a_489_413# 7.36e-20
C1191 VPWR _30_/a_109_53# 9.49e-19
C1192 VPWR _08_ -0.0171f
C1193 net12 _35_/a_226_47# 8.29e-19
C1194 net16 _50_/a_27_47# 2.35e-20
C1195 net13 _33_/a_296_53# 3.71e-20
C1196 _11_ _47_/a_81_21# 0.0454f
C1197 _20_ net6 9.69e-20
C1198 input6/a_27_47# net2 0.0047f
C1199 _53_/a_29_53# net10 7.88e-22
C1200 _26_/a_29_53# net18 2.57e-21
C1201 VGND _37_/a_197_47# -4.58e-19
C1202 net1 _20_ 0.363f
C1203 input13/a_27_47# p[3] 0.00101f
C1204 net1 b[1] 0.0593f
C1205 _35_/a_76_199# _03_ 0.0733f
C1206 _17_ _04_ 4.34e-19
C1207 _22_ _50_/a_27_47# 0.0276f
C1208 net14 _00_ 4.11e-20
C1209 _50_/a_343_93# _47_/a_81_21# 0.00282f
C1210 _20_ _55_/a_472_297# 0.00212f
C1211 _27_/a_27_297# p[10] 1.63e-19
C1212 net7 _02_ 0.445f
C1213 net9 _03_ 0.149f
C1214 _10_ _14_ 0.0571f
C1215 net15 net19 0.0501f
C1216 p[0] net7 1.36e-19
C1217 input2/a_27_47# net1 4.81e-19
C1218 _31_/a_35_297# _02_ 0.00316f
C1219 net3 net8 9.23e-19
C1220 _45_/a_27_47# _03_ 2.06e-20
C1221 p[8] net3 2.13e-19
C1222 _49_/a_201_297# net1 0.00304f
C1223 _01_ _55_/a_217_297# 0.00112f
C1224 net11 _08_ 8.83e-19
C1225 net2 input14/a_27_47# 0.0235f
C1226 _16_ _02_ 0.00564f
C1227 _36_/a_27_47# VGND 0.0209f
C1228 net7 _05_ 0.0129f
C1229 net14 input5/a_381_47# 0.00479f
C1230 VGND _40_/a_109_297# -0.00181f
C1231 p[14] _41_/a_59_75# 5.13e-20
C1232 _33_/a_209_311# _07_ 0.00859f
C1233 _04_ _50_/a_27_47# 2.07e-21
C1234 net9 _50_/a_223_47# 2e-19
C1235 VGND _27_/a_27_297# -0.0157f
C1236 _05_ _31_/a_35_297# 0.00649f
C1237 _13_ _03_ 1.74e-20
C1238 _43_/a_193_413# _44_/a_93_21# 0.0161f
C1239 net3 input15/a_27_47# 8.74e-20
C1240 _30_/a_392_297# net9 9.92e-19
C1241 input10/a_27_47# p[4] 0.0215f
C1242 _47_/a_81_21# _02_ 1.59e-20
C1243 input5/a_664_47# net7 0.00199f
C1244 _16_ _42_/a_209_311# 0.00129f
C1245 net10 _09_ 0.037f
C1246 _44_/a_584_47# VGND -0.00145f
C1247 _21_ _10_ 0.00421f
C1248 _13_ _50_/a_223_47# 8.2e-20
C1249 _10_ net19 0.00224f
C1250 p[13] input5/a_558_47# 0.00156f
C1251 net3 _42_/a_109_93# 0.0435f
C1252 _35_/a_76_199# VGND -0.0034f
C1253 _18_ _39_/a_47_47# 1.23e-19
C1254 _49_/a_544_297# _01_ 0.00109f
C1255 _19_ VPWR 0.0335f
C1256 _44_/a_93_21# _44_/a_250_297# -6.97e-22
C1257 _44_/a_346_47# _44_/a_93_21# -5.12e-20
C1258 _50_/a_615_93# _06_ 0.00264f
C1259 _45_/a_193_297# _39_/a_47_47# 1.4e-20
C1260 _53_/a_111_297# _22_ 4.7e-20
C1261 net12 _30_/a_297_297# 7.14e-21
C1262 input13/a_27_47# p[6] 1.07e-19
C1263 VGND net9 0.372f
C1264 VGND _38_/a_109_47# 2.3e-19
C1265 p[3] _06_ 1.59e-20
C1266 _34_/a_377_297# _21_ 2.37e-19
C1267 _18_ net3 7.34e-20
C1268 VGND _45_/a_27_47# -0.029f
C1269 _15_ net6 0.17f
C1270 VPWR _41_/a_59_75# 0.0179f
C1271 p[2] _04_ 1.9e-20
C1272 net8 input5/a_841_47# 0.025f
C1273 _12_ _11_ 0.195f
C1274 input6/a_27_47# _44_/a_93_21# 8.53e-19
C1275 net7 _55_/a_80_21# 0.00163f
C1276 net8 _17_ 4.52e-20
C1277 _03_ _00_ 2.31e-20
C1278 _11_ _40_/a_297_297# 9.94e-19
C1279 _12_ _35_/a_226_297# 3.35e-20
C1280 net5 _36_/a_197_47# 0.00254f
C1281 _31_/a_35_297# _55_/a_80_21# 5.9e-21
C1282 _11_ _40_/a_191_297# 0.00207f
C1283 _15_ _55_/a_472_297# 0.00626f
C1284 input10/a_27_47# input12/a_27_47# 0.0154f
C1285 _54_/a_75_212# b[1] 0.0023f
C1286 _33_/a_109_93# _35_/a_76_199# 3.08e-19
C1287 _16_ _55_/a_80_21# 0.0143f
C1288 _50_/a_343_93# _12_ 5.63e-20
C1289 _21_ net18 0.00215f
C1290 net16 _11_ 0.172f
C1291 _13_ VGND 0.363f
C1292 VGND input7/a_27_47# 0.0574f
C1293 p[7] net10 5.17e-19
C1294 p[13] output17/a_27_47# 0.00118f
C1295 net11 _19_ 6.27e-21
C1296 _29_/a_29_53# _10_ 5.17e-19
C1297 _01_ _43_/a_27_47# 9.77e-20
C1298 _20_ b[1] 0.00465f
C1299 _50_/a_223_47# _00_ 0.00738f
C1300 net7 net10 1.65e-36
C1301 _33_/a_109_93# net9 0.00211f
C1302 _11_ _22_ 0.15f
C1303 _17_ input15/a_27_47# 6.14e-19
C1304 net10 _31_/a_35_297# 3.95e-20
C1305 _52_/a_93_21# _03_ 0.00985f
C1306 net2 _43_/a_27_47# 0.01f
C1307 VPWR _52_/a_250_297# 0.019f
C1308 _45_/a_465_47# net6 6.06e-20
C1309 net2 p[14] 1.38e-19
C1310 p[1] _19_ 2.91e-20
C1311 _50_/a_343_93# _22_ 0.0597f
C1312 input2/a_27_47# b[1] 0.014f
C1313 _49_/a_201_297# _20_ 5.24e-21
C1314 _17_ _42_/a_109_93# 7.83e-20
C1315 _49_/a_201_297# b[1] 0.0025f
C1316 net12 _36_/a_197_47# 4.67e-20
C1317 net13 _36_/a_303_47# 5.5e-20
C1318 _38_/a_197_47# net4 7.64e-19
C1319 VGND _52_/a_584_47# -0.00112f
C1320 _48_/a_27_47# VPWR 0.0158f
C1321 _12_ _02_ 0.265f
C1322 _21_ _35_/a_489_413# 0.0448f
C1323 _35_/a_226_297# _04_ 4.51e-19
C1324 _18_ _17_ 0.271f
C1325 net16 _02_ 8.94e-19
C1326 output19/a_27_47# b[3] 0.028f
C1327 VGND _00_ 0.139f
C1328 p[6] _06_ 2.49e-19
C1329 _30_/a_215_297# _10_ 5.66e-20
C1330 net11 _52_/a_250_297# 1.2e-19
C1331 _12_ _05_ 2.52e-19
C1332 net13 net3 3.25e-21
C1333 _01_ VPWR 0.521f
C1334 net14 net7 2.23e-19
C1335 _22_ _02_ 0.552f
C1336 net2 VPWR 0.955f
C1337 _23_ VPWR -0.00374f
C1338 p[13] net3 3.64e-19
C1339 net8 p[2] 0.00801f
C1340 VGND input5/a_381_47# -0.0034f
C1341 _22_ _34_/a_47_47# 3.9e-21
C1342 _48_/a_27_47# net11 0.0179f
C1343 _16_ net14 0.00266f
C1344 VGND _52_/a_93_21# -0.0175f
C1345 _05_ _22_ 3.33e-21
C1346 _20_ _15_ 0.691f
C1347 _18_ _50_/a_27_47# 0.0665f
C1348 VGND b[2] 0.0779f
C1349 p[7] p[5] 2.65e-19
C1350 VGND _32_/a_303_47# -4.83e-19
C1351 _38_/a_27_47# output16/a_27_47# 9.02e-19
C1352 _15_ b[1] 1.19e-19
C1353 _42_/a_209_311# _22_ 1.72e-19
C1354 _04_ _02_ 0.0541f
C1355 _09_ _03_ 0.326f
C1356 input5/a_558_47# net19 2.24e-20
C1357 _01_ net11 3.82e-20
C1358 _53_/a_29_53# VGND -0.0168f
C1359 _04_ _34_/a_47_47# 1.17e-20
C1360 _29_/a_183_297# net9 3.51e-19
C1361 net17 _30_/a_109_53# 4.18e-20
C1362 _05_ _04_ 0.0352f
C1363 _23_ net11 0.0461f
C1364 input2/a_27_47# _15_ 3.18e-20
C1365 _44_/a_93_21# p[14] 2.82e-20
C1366 input13/a_27_47# net9 2.42e-19
C1367 _32_/a_27_47# _36_/a_27_47# 0.011f
C1368 _33_/a_109_93# _52_/a_93_21# 2.89e-21
C1369 _26_/a_29_53# net3 2.83e-21
C1370 p[2] _31_/a_285_297# 0.00155f
C1371 net9 _32_/a_109_47# 6.44e-19
C1372 _42_/a_209_311# _04_ 9.84e-22
C1373 p[1] net2 6.12e-20
C1374 input5/a_664_47# _04_ 6.73e-21
C1375 _11_ net8 1.81e-20
C1376 p[8] _11_ 5.85e-20
C1377 net5 net15 0.0226f
C1378 _12_ net10 7.82e-20
C1379 _45_/a_109_297# VGND -0.00179f
C1380 p[13] input5/a_841_47# 1.59e-19
C1381 _36_/a_27_47# _06_ 0.05f
C1382 _55_/a_80_21# _22_ 0.00926f
C1383 _40_/a_109_297# _06_ 0.00175f
C1384 _50_/a_343_93# net8 7.25e-19
C1385 net3 p[9] 1.63e-19
C1386 _28_/a_109_297# _10_ 4.34e-19
C1387 net1 _30_/a_109_53# 0.0297f
C1388 net7 _03_ 0.078f
C1389 _11_ input15/a_27_47# 4.4e-19
C1390 _31_/a_35_297# _03_ 0.00749f
C1391 VGND _09_ 0.396f
C1392 _32_/a_27_47# net9 0.0136f
C1393 net13 _50_/a_27_47# 7.27e-21
C1394 _44_/a_93_21# VPWR 0.005f
C1395 _25_ VPWR 0.0829f
C1396 net5 _10_ 0.199f
C1397 _12_ _39_/a_377_297# 6.77e-19
C1398 _35_/a_76_199# _06_ 0.00425f
C1399 net8 _02_ 0.334f
C1400 net3 _14_ 0.0295f
C1401 net17 _19_ 0.0211f
C1402 _53_/a_183_297# _09_ 4.18e-19
C1403 net7 p[10] 0.00479f
C1404 input10/a_27_47# _54_/a_75_212# 1.17e-22
C1405 net9 _06_ 0.0505f
C1406 _04_ net10 0.121f
C1407 _38_/a_197_47# VPWR -5.24e-19
C1408 _31_/a_35_297# p[10] 2.39e-19
C1409 _33_/a_109_93# _09_ 7.36e-20
C1410 _44_/a_256_47# net3 0.00101f
C1411 _45_/a_27_47# _06_ 0.0021f
C1412 _18_ _11_ 0.484f
C1413 net8 _05_ 0.0146f
C1414 _45_/a_193_297# _11_ 0.0292f
C1415 p[7] VGND 0.195f
C1416 input10/a_27_47# b[1] 0.00691f
C1417 net8 _42_/a_209_311# 7.7e-21
C1418 net11 _25_ 0.0262f
C1419 _50_/a_343_93# _18_ 0.0276f
C1420 VGND net7 0.419f
C1421 net12 _10_ 0.00257f
C1422 _13_ _06_ 0.00187f
C1423 _17_ p[9] 1.03e-20
C1424 VGND _31_/a_35_297# -0.00829f
C1425 input5/a_664_47# net8 0.0116f
C1426 _35_/a_226_47# VPWR 0.00159f
C1427 net14 _22_ 2.23e-19
C1428 _26_/a_29_53# _50_/a_27_47# 5.56e-19
C1429 net3 net19 0.611f
C1430 _01_ _55_/a_300_47# 0.00113f
C1431 _16_ VGND -0.00582f
C1432 _35_/a_556_47# _09_ 0.00122f
C1433 net1 _19_ 2.86e-19
C1434 output18/a_27_47# VPWR 0.0689f
C1435 _31_/a_285_297# _02_ 5.86e-20
C1436 _32_/a_27_47# _00_ 0.00228f
C1437 net6 _41_/a_59_75# 0.0373f
C1438 net12 _34_/a_377_297# 0.00251f
C1439 _49_/a_208_47# VPWR -5.93e-19
C1440 VGND _47_/a_81_21# -0.0112f
C1441 _31_/a_285_297# _05_ 6.12e-19
C1442 net14 _04_ 0.0863f
C1443 _17_ _14_ 0.489f
C1444 _18_ _02_ 2.96e-20
C1445 _35_/a_226_47# net11 3.21e-19
C1446 _52_/a_584_47# _06_ 0.00218f
C1447 _20_ _30_/a_109_53# 8.12e-19
C1448 _45_/a_193_297# _02_ 0.00988f
C1449 net8 _55_/a_80_21# 1.84e-21
C1450 _30_/a_109_53# b[1] 0.00655f
C1451 _08_ b[1] 0.0127f
C1452 net11 output18/a_27_47# 6.84e-20
C1453 _26_/a_111_297# _10_ 7.13e-20
C1454 _06_ _00_ 0.1f
C1455 _29_/a_29_53# net3 1.68e-20
C1456 _07_ _49_/a_75_199# 4.05e-21
C1457 _45_/a_193_297# _05_ 4.84e-22
C1458 net15 p[11] 3.03e-20
C1459 input2/a_27_47# _30_/a_109_53# 1.54e-20
C1460 _01_ input8/a_27_47# 1.43e-19
C1461 net13 _35_/a_226_297# 6.88e-19
C1462 _48_/a_181_47# _02_ 3.9e-19
C1463 _18_ _42_/a_209_311# 3.21e-19
C1464 net8 net10 2.05e-21
C1465 net15 _43_/a_193_413# 0.00169f
C1466 _12_ _03_ 2.76e-20
C1467 net6 _52_/a_250_297# 0.00133f
C1468 _18_ input5/a_664_47# 1.09e-20
C1469 _01_ net17 0.0988f
C1470 _21_ input5/a_841_47# 1.59e-21
C1471 _24_ _10_ 0.00484f
C1472 _29_/a_183_297# _09_ 4.51e-20
C1473 net15 input3/a_27_47# 6.19e-20
C1474 _47_/a_299_297# _00_ 7.59e-21
C1475 _17_ net19 0.0269f
C1476 _52_/a_93_21# _06_ 0.0584f
C1477 input13/a_27_47# _09_ 1.27e-21
C1478 net2 net17 0.261f
C1479 input5/a_381_47# _06_ 1.6e-19
C1480 _12_ _50_/a_223_47# 0.00327f
C1481 _06_ b[2] 0.0116f
C1482 VPWR _30_/a_297_297# -5.22e-19
C1483 _22_ _03_ 2.55e-20
C1484 net12 _35_/a_489_413# 3.97e-20
C1485 net15 _44_/a_250_297# 8.86e-20
C1486 net16 _50_/a_223_47# 4.77e-21
C1487 net13 _33_/a_368_53# 2.1e-20
C1488 net12 _33_/a_296_53# 1.23e-20
C1489 _53_/a_29_53# _06_ 0.0709f
C1490 net5 input5/a_558_47# 0.0597f
C1491 _21_ _50_/a_27_47# 3.38e-21
C1492 _43_/a_193_413# _10_ 0.0174f
C1493 _22_ _50_/a_223_47# 0.031f
C1494 net15 input6/a_27_47# 0.00115f
C1495 _01_ net1 0.0509f
C1496 _26_/a_29_53# _11_ 1.09e-19
C1497 _18_ _55_/a_80_21# 1.44e-20
C1498 _31_/a_285_297# net10 1.68e-19
C1499 net13 _02_ 0.00154f
C1500 _24_ net18 5.57e-21
C1501 _20_ _19_ 0.00734f
C1502 net14 net8 0.0516f
C1503 net1 net2 1.64e-19
C1504 _04_ _03_ 0.586f
C1505 _23_ net6 2.13e-19
C1506 net2 net6 0.00139f
C1507 net13 _34_/a_47_47# 1.68e-19
C1508 p[8] net14 0.0091f
C1509 _26_/a_29_53# _50_/a_343_93# 2.61e-19
C1510 _12_ VGND 0.816f
C1511 p[13] _02_ 7.32e-20
C1512 p[7] input13/a_27_47# 0.0162f
C1513 _19_ b[1] 0.00967f
C1514 _01_ _55_/a_472_297# 6.28e-19
C1515 net13 _05_ 0.192f
C1516 p[13] p[0] 1.88e-19
C1517 _36_/a_109_47# VGND 3.56e-19
C1518 net15 net4 8.68e-19
C1519 VGND _40_/a_191_297# -9.29e-19
C1520 VGND _40_/a_297_297# -5.1e-19
C1521 _04_ _50_/a_223_47# 7.89e-22
C1522 _44_/a_346_47# _10_ 9.13e-21
C1523 _18_ net10 1.47e-21
C1524 _20_ _41_/a_59_75# 1.78e-20
C1525 _45_/a_109_297# _06_ 0.0023f
C1526 _11_ p[9] 1.01e-19
C1527 net16 VGND 0.144f
C1528 input2/a_27_47# _19_ 5.26e-20
C1529 net5 b[0] 3.39e-19
C1530 input9/a_75_212# VPWR 0.0641f
C1531 net5 output17/a_27_47# 5.01e-20
C1532 _36_/a_197_47# VPWR -5.24e-19
C1533 input6/a_27_47# _10_ 4.57e-20
C1534 _30_/a_465_297# net9 0.00138f
C1535 net15 _55_/a_217_297# 7.79e-19
C1536 VGND _22_ 0.0404f
C1537 _27_/a_109_297# VPWR -2.45e-19
C1538 _04_ p[10] 8.48e-21
C1539 _29_/a_29_53# _50_/a_27_47# 1.44e-20
C1540 _06_ _09_ 0.0965f
C1541 p[13] input5/a_664_47# 7.57e-19
C1542 _26_/a_29_53# _02_ 0.0466f
C1543 net14 _42_/a_109_93# 0.00351f
C1544 _33_/a_109_93# _12_ 9.75e-20
C1545 _10_ net4 0.183f
C1546 _49_/a_315_47# VPWR 3.4e-19
C1547 _39_/a_129_47# _00_ 1.63e-20
C1548 _11_ _14_ 0.0415f
C1549 _53_/a_183_297# _22_ 3.71e-20
C1550 _53_/a_111_297# _21_ 4.38e-19
C1551 VGND _04_ 0.135f
C1552 VPWR _41_/a_145_75# -2.46e-19
C1553 _12_ p[12] 6.43e-20
C1554 input9/a_75_212# net11 1.1e-20
C1555 _32_/a_27_47# net7 0.00559f
C1556 _33_/a_109_93# _22_ 1.34e-22
C1557 _18_ net14 0.0147f
C1558 _07_ p[6] 1.27e-19
C1559 net5 _36_/a_303_47# 0.00256f
C1560 _10_ _55_/a_217_297# 1.43e-19
C1561 _50_/a_343_93# _14_ 9.76e-19
C1562 _32_/a_27_47# _31_/a_35_297# 9.17e-20
C1563 _48_/a_27_47# b[1] 0.00666f
C1564 p[7] _06_ 0.00863f
C1565 _33_/a_209_311# _35_/a_76_199# 9.95e-21
C1566 _15_ _19_ 1.46e-20
C1567 net5 _39_/a_47_47# 0.0389f
C1568 net8 _03_ 0.0287f
C1569 net13 net10 0.375f
C1570 _22_ p[12] 2.13e-21
C1571 net7 _06_ 0.00447f
C1572 _11_ net19 2.19e-19
C1573 _21_ _11_ 9.98e-20
C1574 _44_/a_93_21# net6 1.08e-20
C1575 _33_/a_209_311# net9 4.33e-20
C1576 _33_/a_109_93# _04_ 0.0299f
C1577 _42_/a_209_311# p[9] 5.51e-21
C1578 _01_ _20_ 0.161f
C1579 _15_ _41_/a_59_75# 0.0139f
C1580 _01_ b[1] 0.00233f
C1581 _32_/a_27_47# _47_/a_81_21# 5.06e-21
C1582 _16_ _06_ 0.00162f
C1583 net5 net3 0.0365f
C1584 VPWR _52_/a_256_47# -9.47e-19
C1585 _20_ net2 8.83e-19
C1586 _23_ b[1] 7.65e-19
C1587 net2 b[1] 0.0389f
C1588 _14_ _02_ 0.0316f
C1589 net12 _36_/a_303_47# 1.37e-19
C1590 net15 p[14] 0.00137f
C1591 _38_/a_303_47# net4 5.95e-19
C1592 net8 p[10] 0.00463f
C1593 _01_ _49_/a_201_297# 0.0105f
C1594 input2/a_27_47# net2 0.024f
C1595 _26_/a_183_297# _10_ 5.74e-19
C1596 _06_ _47_/a_81_21# 0.0388f
C1597 _31_/a_285_297# _03_ 0.00677f
C1598 _42_/a_209_311# _14_ 0.00142f
C1599 _37_/a_27_47# _00_ 6.15e-20
C1600 _26_/a_29_53# net10 3.48e-22
C1601 net1 _35_/a_226_47# 1.3e-20
C1602 net13 net14 2.21e-21
C1603 VGND net8 0.405f
C1604 p[8] VGND 0.0828f
C1605 net19 _02_ 0.0474f
C1606 _18_ _03_ 7.25e-23
C1607 _21_ _02_ 0.397f
C1608 _43_/a_27_47# _10_ 0.0279f
C1609 _10_ p[14] 1.53e-19
C1610 p[13] net14 1.89e-19
C1611 _45_/a_193_297# _03_ 2.57e-20
C1612 _21_ _34_/a_47_47# 8.93e-19
C1613 _21_ _05_ 0.0104f
C1614 _42_/a_109_93# p[10] 1.82e-21
C1615 net5 input5/a_841_47# 0.0221f
C1616 _18_ _50_/a_223_47# 0.0367f
C1617 net15 VPWR 0.61f
C1618 net13 p[5] 1.05e-19
C1619 net5 _17_ 0.00408f
C1620 VGND input15/a_27_47# 0.0156f
C1621 _42_/a_209_311# net19 0.0766f
C1622 _01_ _15_ 0.007f
C1623 input3/a_27_47# output17/a_27_47# 3.15e-19
C1624 input5/a_664_47# net19 1.38e-21
C1625 _21_ input5/a_664_47# 9.42e-22
C1626 _55_/a_80_21# _14_ 0.0175f
C1627 _29_/a_183_297# _04_ 0.0015f
C1628 _35_/a_76_199# _07_ 0.00226f
C1629 VGND _42_/a_109_93# -0.0045f
C1630 net2 _15_ 9.8e-19
C1631 _13_ output16/a_27_47# 4.58e-19
C1632 _26_/a_29_53# net14 1.33e-20
C1633 _54_/a_75_212# _25_ 0.0247f
C1634 VGND _31_/a_285_297# -0.00136f
C1635 _07_ net9 1.39e-20
C1636 _29_/a_29_53# _02_ 6.76e-21
C1637 net5 _50_/a_27_47# 0.0169f
C1638 net9 _32_/a_197_47# 6.06e-19
C1639 _25_ b[1] 0.0015f
C1640 _45_/a_27_47# _07_ 1.02e-20
C1641 _10_ VPWR 0.577f
C1642 _18_ VGND 0.0166f
C1643 _32_/a_27_47# _22_ 1.76e-19
C1644 _29_/a_29_53# _05_ 3.79e-20
C1645 _12_ _06_ 0.136f
C1646 _45_/a_193_297# VGND -0.00241f
C1647 net14 p[9] 1.05e-19
C1648 net15 p[1] 6.22e-20
C1649 _36_/a_109_47# _06_ 0.00168f
C1650 _13_ _07_ 3.22e-23
C1651 _40_/a_191_297# _06_ 5.84e-19
C1652 _06_ _40_/a_297_297# 1.64e-19
C1653 _55_/a_80_21# net19 0.00423f
C1654 input15/a_27_47# p[12] 5.48e-19
C1655 net1 _30_/a_297_297# 7.34e-20
C1656 net13 _03_ 0.271f
C1657 net16 _06_ 0.0511f
C1658 _34_/a_377_297# VPWR -0.00192f
C1659 net13 _34_/a_285_47# 4.11e-20
C1660 _31_/a_117_297# _03_ 5.32e-19
C1661 input9/a_75_212# input8/a_27_47# 3.09e-20
C1662 _48_/a_181_47# VGND 3.03e-19
C1663 net3 p[11] 0.00296f
C1664 _12_ _47_/a_299_297# 0.00805f
C1665 b[0] net4 0.0024f
C1666 _21_ net10 0.0275f
C1667 net11 _10_ 0.0109f
C1668 _22_ _06_ 0.124f
C1669 _32_/a_27_47# _04_ 1.43e-19
C1670 _20_ _35_/a_226_47# 5.19e-20
C1671 net12 _50_/a_27_47# 7.99e-21
C1672 net3 _43_/a_193_413# 5.65e-20
C1673 net18 VPWR 0.104f
C1674 _30_/a_215_297# _02_ 3.58e-21
C1675 _35_/a_226_47# b[1] 0.00334f
C1676 _54_/a_75_212# output18/a_27_47# 2.28e-19
C1677 net13 _30_/a_392_297# 6.64e-20
C1678 net3 input3/a_27_47# 0.03f
C1679 net14 _14_ 0.184f
C1680 _18_ p[12] 4.76e-21
C1681 output18/a_27_47# b[1] 9.26e-19
C1682 _30_/a_215_297# _05_ 0.0453f
C1683 _33_/a_209_311# _09_ 3.79e-20
C1684 _04_ _06_ 0.0132f
C1685 _44_/a_346_47# net3 8.04e-19
C1686 _44_/a_256_47# net14 0.00379f
C1687 _38_/a_303_47# VPWR -4.83e-19
C1688 _49_/a_201_297# _35_/a_226_47# 1.66e-20
C1689 net3 _44_/a_250_297# 0.0088f
C1690 _45_/a_205_47# _10_ 6.19e-20
C1691 p[13] p[10] 0.00177f
C1692 _49_/a_208_47# b[1] 2.93e-19
C1693 _26_/a_29_53# _03_ 7.93e-21
C1694 _44_/a_93_21# _15_ 0.0168f
C1695 input9/a_75_212# net1 0.002f
C1696 _11_ _28_/a_109_297# 6.29e-19
C1697 _36_/a_197_47# net6 6.94e-20
C1698 net11 net18 0.00221f
C1699 net13 VGND 0.142f
C1700 net3 input6/a_27_47# 2.52e-19
C1701 net8 _32_/a_109_47# 0.0011f
C1702 _29_/a_29_53# net10 1.77e-19
C1703 _35_/a_489_413# VPWR -0.00725f
C1704 _26_/a_29_53# _50_/a_223_47# 0.00124f
C1705 net4 _39_/a_47_47# 0.0202f
C1706 net14 _21_ 7.17e-21
C1707 VGND _31_/a_117_297# -0.00177f
C1708 _16_ _37_/a_27_47# 2.07e-19
C1709 net14 net19 0.148f
C1710 _33_/a_296_53# VPWR -1.15e-19
C1711 p[13] VGND 0.0912f
C1712 _13_ _38_/a_27_47# 4.58e-19
C1713 net5 _11_ 0.207f
C1714 net3 net4 9.28e-21
C1715 input4/a_75_212# _45_/a_27_47# 2.18e-20
C1716 p[7] _33_/a_209_311# 9.77e-20
C1717 net15 _55_/a_300_47# 1.09e-19
C1718 _48_/a_27_47# _08_ 2.58e-19
C1719 net3 input14/a_27_47# 9.36e-19
C1720 _43_/a_193_413# _17_ 0.0503f
C1721 _50_/a_343_93# net5 0.00124f
C1722 net13 _33_/a_109_93# 0.0254f
C1723 _31_/a_285_47# _05_ 5.61e-19
C1724 net3 _55_/a_217_297# 5.78e-20
C1725 _32_/a_27_47# net8 0.0275f
C1726 _44_/a_584_47# b[3] 1.26e-19
C1727 _30_/a_297_297# b[1] 3.14e-19
C1728 net15 _27_/a_277_297# 1.93e-19
C1729 _12_ _39_/a_129_47# 0.00175f
C1730 _26_/a_29_53# VGND 0.0381f
C1731 _44_/a_346_47# _17_ 7.2e-19
C1732 _30_/a_215_297# net10 0.0512f
C1733 _17_ _44_/a_250_297# 0.0336f
C1734 _29_/a_29_53# net14 1.61e-20
C1735 input5/a_558_47# VPWR 0.0083f
C1736 net12 _11_ 3.82e-21
C1737 net8 _06_ 0.00282f
C1738 _23_ _08_ 1.81e-19
C1739 net5 _02_ 0.233f
C1740 input6/a_27_47# _17_ 7.13e-22
C1741 _47_/a_384_47# _00_ 5.15e-20
C1742 VGND p[9] 0.0725f
C1743 _17_ net4 7.52e-21
C1744 input5/a_62_47# net9 3.12e-19
C1745 _21_ _03_ 0.0818f
C1746 _07_ _09_ 0.0416f
C1747 _24_ _53_/a_111_297# 9.08e-21
C1748 input15/a_27_47# _06_ 4.73e-19
C1749 net15 net17 5.19e-19
C1750 net5 _42_/a_209_311# 3.27e-21
C1751 _34_/a_285_47# _21_ 6.94e-20
C1752 net12 _33_/a_368_53# 2.63e-19
C1753 b[0] VPWR 0.142f
C1754 input9/a_75_212# b[1] 0.00598f
C1755 _27_/a_27_297# _49_/a_75_199# 0.011f
C1756 _32_/a_27_47# _18_ 1.18e-20
C1757 output17/a_27_47# VPWR 0.0268f
C1758 net5 input5/a_664_47# 0.0536f
C1759 input10/a_27_47# _25_ 2.03e-20
C1760 _43_/a_297_47# _10_ 0.00118f
C1761 _21_ _50_/a_223_47# 2.91e-21
C1762 _42_/a_109_93# _06_ 5.53e-20
C1763 _27_/a_109_297# b[1] 8.35e-20
C1764 net12 _02_ 2.28e-19
C1765 VGND _14_ 0.226f
C1766 p[1] input5/a_558_47# 1.61e-21
C1767 _31_/a_285_297# _06_ 1.01e-20
C1768 _53_/a_29_53# _38_/a_27_47# 1.29e-19
C1769 net12 _34_/a_47_47# 0.0385f
C1770 _28_/a_109_297# _55_/a_80_21# 2.05e-20
C1771 net3 p[14] 0.00446f
C1772 net4 _50_/a_27_47# 0.0239f
C1773 _44_/a_256_47# VGND -0.00184f
C1774 _13_ _39_/a_285_47# 0.00451f
C1775 p[10] net19 1.26e-21
C1776 net13 input13/a_27_47# 0.00139f
C1777 net12 _05_ 0.0414f
C1778 _24_ _11_ 7.29e-20
C1779 _18_ _06_ 0.54f
C1780 p[9] p[12] 1.4e-19
C1781 _49_/a_315_47# b[1] 5.66e-19
C1782 net15 net1 7.44e-20
C1783 _01_ _19_ 0.031f
C1784 _45_/a_193_297# _06_ 0.00201f
C1785 net15 net6 0.0664f
C1786 net2 _19_ 0.101f
C1787 net9 _49_/a_75_199# 0.00382f
C1788 _29_/a_29_53# _03_ 0.0414f
C1789 net5 _55_/a_80_21# 2.78e-19
C1790 input1/a_75_212# input7/a_27_47# 3.2e-20
C1791 _36_/a_303_47# VPWR -4.83e-19
C1792 _52_/a_93_21# _52_/a_346_47# -5.12e-20
C1793 _21_ VGND 0.295f
C1794 VGND net19 0.133f
C1795 input11/a_27_47# p[5] 0.0433f
C1796 _27_/a_205_297# VPWR 1.05e-19
C1797 _48_/a_181_47# _06_ 6.4e-19
C1798 _39_/a_47_47# VPWR 0.0668f
C1799 _29_/a_29_53# _50_/a_223_47# 1.45e-20
C1800 _33_/a_209_311# _12_ 2.88e-20
C1801 _43_/a_193_413# _11_ 5.45e-19
C1802 net5 net10 0.0316f
C1803 _10_ net6 0.0965f
C1804 net1 _10_ 4.34e-19
C1805 net3 VPWR 0.351f
C1806 _38_/a_27_47# _09_ 0.00195f
C1807 b[1] _52_/a_256_47# 8.49e-20
C1808 _39_/a_285_47# _00_ 1.47e-21
C1809 _36_/a_303_47# net11 7.63e-20
C1810 _24_ _02_ 0.0232f
C1811 _33_/a_109_93# _21_ 1.62e-20
C1812 _10_ _55_/a_472_297# 7.35e-21
C1813 _24_ _34_/a_47_47# 6.84e-21
C1814 _17_ _43_/a_27_47# 0.00131f
C1815 _53_/a_111_297# net4 2.09e-19
C1816 _23_ _52_/a_250_297# 3.17e-19
C1817 _17_ p[14] 5.46e-21
C1818 _32_/a_27_47# p[13] 6.49e-20
C1819 net9 p[3] 0.0375f
C1820 _30_/a_215_297# _03_ 0.0393f
C1821 net5 _39_/a_377_297# 0.00234f
C1822 _29_/a_29_53# VGND 0.0544f
C1823 _35_/a_226_47# _08_ 0.00117f
C1824 net19 p[12] 6.8e-20
C1825 net13 _06_ 0.0758f
C1826 net12 net10 0.539f
C1827 _33_/a_209_311# _04_ 0.00133f
C1828 _21_ _35_/a_556_47# 2.69e-19
C1829 net5 net14 0.0263f
C1830 _43_/a_193_413# _02_ 9.4e-21
C1831 _11_ net4 0.0858f
C1832 _01_ net2 2.72e-19
C1833 _42_/a_209_311# p[11] 2.58e-19
C1834 _11_ input14/a_27_47# 1.42e-19
C1835 net15 _20_ 0.0021f
C1836 input5/a_841_47# VPWR 0.0775f
C1837 net15 b[1] 0.00314f
C1838 _17_ VPWR 0.306f
C1839 _50_/a_343_93# net4 0.00124f
C1840 net16 output16/a_27_47# 0.0101f
C1841 input3/a_27_47# _42_/a_209_311# 1.56e-19
C1842 _31_/a_285_47# _03_ 8.54e-19
C1843 _30_/a_215_297# VGND 0.00687f
C1844 input2/a_27_47# net15 1.61e-19
C1845 _26_/a_29_53# _06_ 0.0135f
C1846 net15 _49_/a_201_297# 1.41e-19
C1847 _12_ _07_ 2.94e-23
C1848 _37_/a_27_47# p[8] 9.82e-21
C1849 _37_/a_27_47# net8 6.66e-21
C1850 VGND input11/a_27_47# 0.0274f
C1851 p[8] output19/a_27_47# 0.00805f
C1852 _20_ _10_ 0.179f
C1853 _50_/a_27_47# VPWR -0.00335f
C1854 input5/a_558_47# net17 2.88e-21
C1855 _10_ b[1] 2.37e-20
C1856 p[11] _55_/a_80_21# 6.43e-20
C1857 net4 _02_ 0.00376f
C1858 _06_ p[9] 0.00205f
C1859 _37_/a_27_47# input15/a_27_47# 3.27e-19
C1860 _07_ _22_ 1.19e-20
C1861 net12 p[5] 0.00294f
C1862 _33_/a_109_93# _30_/a_215_297# 0.00104f
C1863 _42_/a_296_53# net19 2.71e-19
C1864 _43_/a_193_413# _55_/a_80_21# 2.54e-19
C1865 _55_/a_217_297# _02_ 6.01e-19
C1866 net5 _03_ 1.04e-19
C1867 _34_/a_377_297# b[1] 0.00115f
C1868 _49_/a_208_47# _19_ 7.12e-20
C1869 _37_/a_27_47# _42_/a_109_93# 2.55e-20
C1870 output19/a_27_47# _42_/a_109_93# 1.56e-20
C1871 net3 _42_/a_368_53# 3.82e-19
C1872 VGND _31_/a_285_47# 8.88e-34
C1873 _54_/a_75_212# net18 0.0143f
C1874 net11 _50_/a_27_47# 6.05e-21
C1875 input5/a_558_47# net1 1.1e-19
C1876 _09_ _49_/a_75_199# 2.93e-19
C1877 net5 _50_/a_223_47# 0.00202f
C1878 net15 _15_ 0.156f
C1879 net17 output17/a_27_47# 0.0149f
C1880 input5/a_62_47# net7 2.04e-19
C1881 _07_ _04_ 9.74e-20
C1882 _14_ _06_ 0.0556f
C1883 p[2] VPWR 0.102f
C1884 net18 b[1] 0.00134f
C1885 _11_ _43_/a_27_47# 4.27e-19
C1886 _35_/a_226_47# _52_/a_250_297# 2.63e-20
C1887 _37_/a_27_47# _18_ 3.31e-20
C1888 _32_/a_27_47# _21_ 8.95e-19
C1889 net2 _44_/a_93_21# 0.0273f
C1890 net5 p[10] 5.12e-21
C1891 _36_/a_27_47# _35_/a_76_199# 3.22e-19
C1892 _23_ _25_ 0.00465f
C1893 VGND _28_/a_109_297# -9.87e-19
C1894 net3 _27_/a_277_297# 2.71e-19
C1895 _53_/a_111_297# VPWR 1.11e-34
C1896 net12 _34_/a_285_47# 8.07e-20
C1897 net12 _03_ 0.0268f
C1898 _12_ _38_/a_27_47# 0.0527f
C1899 net7 input1/a_75_212# 3.77e-19
C1900 _34_/a_129_47# VPWR -9.47e-19
C1901 _36_/a_27_47# net9 0.00493f
C1902 _12_ _47_/a_384_47# 9.51e-20
C1903 net14 p[11] 1.9e-19
C1904 net4 _55_/a_80_21# 1.06e-19
C1905 b[0] net6 2.52e-19
C1906 _15_ _10_ 0.479f
C1907 net1 output17/a_27_47# 8.12e-19
C1908 _21_ _06_ 0.143f
C1909 net16 _38_/a_27_47# 0.114f
C1910 net19 _06_ 0.00522f
C1911 net5 VGND 1.2f
C1912 net14 _43_/a_193_413# 1.11e-19
C1913 _35_/a_489_413# b[1] 0.00104f
C1914 net7 _49_/a_75_199# 0.09f
C1915 _48_/a_109_47# net11 1.74e-19
C1916 net14 input3/a_27_47# 3.47e-19
C1917 _55_/a_217_297# _55_/a_80_21# 1.42e-32
C1918 _38_/a_27_47# _22_ 2.86e-19
C1919 input4/a_75_212# _12_ 2.09e-20
C1920 _33_/a_296_53# b[1] 2.69e-20
C1921 net12 _30_/a_392_297# 2.19e-20
C1922 net13 _30_/a_465_297# 6.36e-20
C1923 _31_/a_35_297# _49_/a_75_199# 6.24e-19
C1924 net4 net10 8.28e-22
C1925 p[1] p[2] 0.0525f
C1926 _35_/a_226_297# VPWR -8.54e-19
C1927 _43_/a_27_47# _02_ 1.88e-21
C1928 _11_ VPWR 0.352f
C1929 _23_ _35_/a_226_47# 4.21e-19
C1930 net3 net17 3.72e-19
C1931 _27_/a_27_297# input7/a_27_47# 0.00119f
C1932 _35_/a_76_199# _45_/a_27_47# 2.04e-21
C1933 _34_/a_129_47# net11 0.00242f
C1934 net14 _44_/a_250_297# 4.24e-20
C1935 _44_/a_346_47# net14 0.00464f
C1936 _50_/a_343_93# VPWR -0.0126f
C1937 _45_/a_465_47# _10_ 3.32e-19
C1938 _49_/a_208_47# _01_ 2.13e-19
C1939 _36_/a_303_47# net6 1.25e-19
C1940 net12 VGND 0.344f
C1941 _37_/a_303_47# VPWR -3.13e-19
C1942 net8 _32_/a_197_47# 3.39e-20
C1943 _12_ _52_/a_346_47# 3.8e-19
C1944 _13_ _35_/a_76_199# 3.01e-21
C1945 _42_/a_209_311# p[14] 3.45e-22
C1946 net14 input6/a_27_47# 7.05e-19
C1947 _24_ _03_ 9.46e-20
C1948 _29_/a_29_53# _06_ 0.00111f
C1949 net4 _39_/a_377_297# 8.88e-19
C1950 net6 _39_/a_47_47# 0.0249f
C1951 _33_/a_368_53# VPWR -4.26e-19
C1952 p[7] p[3] 0.0366f
C1953 net5 p[12] 4.99e-20
C1954 input5/a_558_47# b[1] 0.00214f
C1955 net3 net1 4.25e-20
C1956 _27_/a_109_297# _19_ 7.54e-21
C1957 net14 net4 2.21e-21
C1958 _13_ _45_/a_27_47# 0.0703f
C1959 net3 net6 0.00152f
C1960 net14 input14/a_27_47# 0.0232f
C1961 _43_/a_297_47# _17_ 5.72e-20
C1962 VPWR _02_ 0.332f
C1963 p[0] VPWR 0.0834f
C1964 net12 _33_/a_109_93# 0.0435f
C1965 input2/a_27_47# input5/a_558_47# 2.04e-20
C1966 net13 _33_/a_209_311# 0.0227f
C1967 VPWR _34_/a_47_47# 0.0372f
C1968 _05_ VPWR 0.118f
C1969 net14 _55_/a_217_297# 2.1e-19
C1970 _49_/a_315_47# _19_ 1.33e-19
C1971 _26_/a_111_297# VGND -2.75e-19
C1972 _43_/a_27_47# _55_/a_80_21# 1.56e-19
C1973 _12_ _39_/a_285_47# 0.0221f
C1974 input5/a_381_47# _27_/a_27_297# 1.47e-19
C1975 _42_/a_209_311# VPWR -0.00753f
C1976 _30_/a_215_297# _06_ 2.03e-20
C1977 output17/a_27_47# b[1] 0.0373f
C1978 input5/a_664_47# VPWR 0.00488f
C1979 net11 _02_ 0.0327f
C1980 net16 _39_/a_285_47# 1.29e-19
C1981 _18_ _43_/a_369_47# 1.49e-19
C1982 net9 _00_ 0.00501f
C1983 _24_ VGND -0.00863f
C1984 p[11] p[10] 0.0074f
C1985 net11 _34_/a_47_47# 0.0309f
C1986 _45_/a_27_47# _00_ 4.84e-20
C1987 _37_/a_27_47# p[9] 0.0117f
C1988 input2/a_27_47# output17/a_27_47# 0.107f
C1989 net11 _05_ 2.76e-19
C1990 _35_/a_76_199# _52_/a_93_21# 6.83e-21
C1991 output19/a_27_47# p[9] 0.0832f
C1992 p[7] p[6] 0.0717f
C1993 p[1] p[0] 0.053f
C1994 net1 input5/a_841_47# 1.33e-19
C1995 _48_/a_181_47# _07_ 5.93e-19
C1996 output18/a_27_47# _25_ 0.072f
C1997 input5/a_62_47# _04_ 0.00345f
C1998 input5/a_381_47# net9 3.4e-19
C1999 VGND p[11] 0.148f
C2000 _17_ net6 3.12e-19
C2001 _13_ _00_ 3.77e-20
C2002 input5/a_558_47# _15_ 0.00166f
C2003 _45_/a_27_47# _52_/a_93_21# 1.18e-19
C2004 _32_/a_303_47# net9 0.00218f
C2005 net5 _32_/a_109_47# 5.69e-21
C2006 _55_/a_80_21# VPWR 0.0289f
C2007 _43_/a_193_413# VGND -0.0147f
C2008 input10/a_27_47# net18 4.16e-20
C2009 _22_ _49_/a_75_199# 9.85e-21
C2010 input3/a_27_47# VGND 0.0414f
C2011 _20_ _39_/a_47_47# 2.3e-20
C2012 _27_/a_205_297# b[1] 1.41e-19
C2013 output19/a_27_47# _14_ 1.43e-19
C2014 _37_/a_27_47# _14_ 0.00137f
C2015 _10_ _08_ 1.51e-19
C2016 _13_ _52_/a_93_21# 1.31e-19
C2017 p[1] input5/a_664_47# 1.21e-20
C2018 net10 VPWR 0.375f
C2019 net14 _43_/a_27_47# 4.87e-20
C2020 net4 _50_/a_223_47# 0.0107f
C2021 net6 _50_/a_27_47# 0.0428f
C2022 net14 p[14] 6.11e-20
C2023 p[2] input8/a_27_47# 0.0163f
C2024 net2 _27_/a_109_297# 7.24e-20
C2025 _44_/a_346_47# VGND -0.00198f
C2026 VGND _44_/a_250_297# -0.00591f
C2027 net3 _20_ 4.07e-19
C2028 input4/a_75_212# input15/a_27_47# 1.1e-21
C2029 net12 input13/a_27_47# 0.0163f
C2030 net3 b[1] 0.00334f
C2031 _13_ _53_/a_29_53# 9.05e-19
C2032 _01_ _49_/a_315_47# 1.82e-19
C2033 net13 _07_ 0.00686f
C2034 _04_ _49_/a_75_199# 0.0782f
C2035 _32_/a_27_47# net5 0.0961f
C2036 input6/a_27_47# VGND -0.00259f
C2037 _29_/a_111_297# _03_ 7.48e-19
C2038 _37_/a_27_47# net19 0.0105f
C2039 net15 _19_ 0.00628f
C2040 output19/a_27_47# net19 0.0273f
C2041 p[8] b[3] 0.00229f
C2042 _35_/a_76_199# _09_ 0.047f
C2043 net11 net10 0.592f
C2044 net5 _06_ 0.41f
C2045 _49_/a_544_297# _03_ 0.00568f
C2046 net15 _41_/a_59_75# 1.16e-20
C2047 VGND net4 0.564f
C2048 net9 _09_ 2.62e-19
C2049 VGND input14/a_27_47# 0.0389f
C2050 input4/a_75_212# _18_ 4.36e-19
C2051 net1 p[2] 0.0269f
C2052 net14 VPWR 0.182f
C2053 _45_/a_27_47# _09_ 0.00823f
C2054 input15/a_27_47# b[3] 0.00109f
C2055 net8 input5/a_62_47# 2.05e-19
C2056 p[8] input5/a_62_47# 1.22e-19
C2057 _55_/a_300_47# _02_ 0.00371f
C2058 VGND _55_/a_217_297# -0.00342f
C2059 net12 _32_/a_27_47# 1.52e-19
C2060 net5 _47_/a_299_297# 0.00198f
C2061 net7 _27_/a_27_297# 1.22e-19
C2062 _15_ _27_/a_205_297# 5.5e-20
C2063 _04_ p[3] 2.34e-21
C2064 _16_ _27_/a_27_297# 3.74e-22
C2065 input12/a_27_47# _02_ 1.88e-19
C2066 _23_ _52_/a_256_47# 6.66e-19
C2067 _13_ _09_ 0.0927f
C2068 input5/a_841_47# b[1] 7.07e-19
C2069 _20_ _17_ 0.102f
C2070 _52_/a_93_21# b[2] 1.63e-19
C2071 input6/a_27_47# p[12] 2.78e-19
C2072 input12/a_27_47# _34_/a_47_47# 2.17e-19
C2073 _29_/a_111_297# VGND -1.9e-19
C2074 p[5] VPWR 0.0923f
C2075 net12 _06_ 0.284f
C2076 _35_/a_489_413# _08_ 5.56e-19
C2077 _10_ _41_/a_59_75# 0.0172f
C2078 _35_/a_76_199# net7 1.79e-20
C2079 net14 net11 9.95e-19
C2080 net3 _15_ 0.224f
C2081 _36_/a_197_47# _25_ 2.37e-21
C2082 _53_/a_29_53# _52_/a_93_21# 0.00116f
C2083 p[7] net9 8.26e-19
C2084 _53_/a_29_53# b[2] 6.22e-19
C2085 net4 p[12] 0.00758f
C2086 net7 net9 0.00233f
C2087 _45_/a_109_297# _00_ 4.86e-20
C2088 net8 _49_/a_75_199# 0.00214f
C2089 _49_/a_544_297# VGND -0.00256f
C2090 _11_ net6 0.0257f
C2091 p[4] net10 0.00268f
C2092 net14 p[1] 0.0025f
C2093 input8/a_27_47# _02_ 5.08e-20
C2094 net11 p[5] 0.0598f
C2095 _26_/a_183_297# VGND 2.42e-19
C2096 _50_/a_343_93# net6 0.00214f
C2097 _50_/a_429_93# net4 4.16e-19
C2098 net17 _02_ 0.0608f
C2099 _09_ _00_ 9.35e-21
C2100 _10_ _52_/a_250_297# 0.00368f
C2101 _05_ input8/a_27_47# 1.58e-19
C2102 net15 _01_ 0.0314f
C2103 net7 input7/a_27_47# 0.00318f
C2104 net17 _05_ 0.0111f
C2105 VPWR _03_ 0.835f
C2106 net15 net2 0.324f
C2107 _26_/a_111_297# _06_ 9e-19
C2108 _43_/a_369_47# _14_ 0.00135f
C2109 net9 _47_/a_81_21# 3.49e-19
C2110 _34_/a_285_47# VPWR -0.00233f
C2111 _48_/a_27_47# _10_ 4.55e-19
C2112 _52_/a_93_21# _09_ 0.0227f
C2113 VGND p[14] 0.366f
C2114 VGND _43_/a_27_47# -0.0153f
C2115 _42_/a_209_311# net17 1.04e-21
C2116 _09_ b[2] 4.28e-20
C2117 _50_/a_223_47# VPWR -0.00601f
C2118 _24_ _06_ 0.113f
C2119 net8 p[3] 0.0015f
C2120 _17_ _15_ 0.0752f
C2121 p[2] b[1] 0.00188f
C2122 net1 _02_ 0.00251f
C2123 net5 _39_/a_129_47# 0.00344f
C2124 net6 _02_ 0.00427f
C2125 p[0] net1 0.00473f
C2126 net10 input12/a_27_47# 0.00182f
C2127 _33_/a_209_311# _30_/a_215_297# 1.56e-19
C2128 _01_ _10_ 2.22e-19
C2129 _48_/a_109_47# b[1] 9.32e-20
C2130 _21_ _07_ 0.133f
C2131 _37_/a_109_47# net19 1.16e-20
C2132 _53_/a_29_53# _09_ 0.00642f
C2133 _34_/a_285_47# net11 -7.11e-33
C2134 p[10] VPWR 0.234f
C2135 net1 _05_ 0.151f
C2136 net11 _03_ 0.0952f
C2137 _55_/a_472_297# _02_ 1.25e-19
C2138 net2 _10_ 3.15e-19
C2139 _23_ _10_ 0.00192f
C2140 net7 _00_ 8.12e-21
C2141 _36_/a_27_47# _12_ 0.00178f
C2142 _49_/a_201_297# p[2] 4.58e-20
C2143 _16_ _00_ 0.00613f
C2144 _34_/a_129_47# b[1] 3.51e-19
C2145 net14 _42_/a_368_53# 7.39e-19
C2146 _42_/a_209_311# net6 1.32e-20
C2147 _43_/a_193_413# _06_ 0.0138f
C2148 _15_ _50_/a_27_47# 5.65e-19
C2149 p[4] p[5] 0.249f
C2150 input5/a_664_47# net1 2.41e-19
C2151 p[14] p[12] 0.00101f
C2152 VGND VPWR -0.454f
C2153 input5/a_381_47# net7 4.91e-19
C2154 _36_/a_27_47# _22_ 2.82e-20
C2155 _54_/a_75_212# _11_ 3.22e-20
C2156 p[13] input5/a_62_47# 0.0201f
C2157 _47_/a_81_21# _00_ 0.0258f
C2158 _11_ _20_ 0.268f
C2159 net17 net10 8.67e-21
C2160 _35_/a_76_199# _12_ 6.84e-20
C2161 _35_/a_226_297# b[1] 1.03e-19
C2162 _23_ net18 -4.05e-24
C2163 net14 _27_/a_277_297# 5.1e-19
C2164 _29_/a_29_53# _07_ 1.19e-20
C2165 _50_/a_343_93# _20_ 0.00826f
C2166 net15 _44_/a_93_21# 0.00573f
C2167 _12_ net9 4.39e-22
C2168 _12_ _38_/a_109_47# 0.00179f
C2169 p[1] p[10] 1.8e-20
C2170 _36_/a_27_47# _04_ 0.00169f
C2171 _33_/a_109_93# VPWR -0.00817f
C2172 VGND net11 0.475f
C2173 _12_ _45_/a_27_47# 0.0867f
C2174 input6/a_27_47# _06_ 2.85e-19
C2175 net1 _55_/a_80_21# 1.8e-19
C2176 _35_/a_76_199# _22_ 6.58e-21
C2177 p[13] input1/a_75_212# 4.16e-19
C2178 _27_/a_27_297# _04_ 0.0526f
C2179 _37_/a_27_47# net5 1.13e-20
C2180 net16 _45_/a_27_47# 8.68e-19
C2181 net16 _38_/a_109_47# 4.17e-19
C2182 net13 _49_/a_75_199# 3.2e-19
C2183 net14 _43_/a_297_47# 1.09e-21
C2184 b[3] p[9] 0.107f
C2185 input12/a_27_47# p[5] 0.00359f
C2186 net9 _22_ 0.0023f
C2187 _13_ _12_ 0.462f
C2188 VPWR p[12] 0.0376f
C2189 p[1] VGND 0.137f
C2190 net12 _30_/a_465_297# 8.01e-20
C2191 net1 net10 0.00388f
C2192 _33_/a_368_53# b[1] 4.19e-19
C2193 _21_ _38_/a_27_47# 3.87e-19
C2194 net6 net10 1.35e-20
C2195 net4 _06_ 0.281f
C2196 output17/a_27_47# _19_ 7.69e-19
C2197 _54_/a_75_212# _02_ 6.6e-20
C2198 _45_/a_27_47# _22_ 0.0131f
C2199 _35_/a_556_47# VPWR -7.24e-19
C2200 _44_/a_93_21# _10_ 2.48e-19
C2201 _20_ _02_ 0.1f
C2202 _13_ net16 0.0198f
C2203 _35_/a_76_199# _04_ 0.0269f
C2204 _45_/a_205_47# VGND -2.47e-19
C2205 p[7] _09_ 9.25e-21
C2206 _02_ b[1] 0.00718f
C2207 net14 net17 5.43e-19
C2208 _33_/a_109_93# net11 5.14e-19
C2209 _50_/a_429_93# VPWR -3.61e-19
C2210 _55_/a_217_297# _06_ 3.46e-19
C2211 _10_ _25_ 0.0109f
C2212 p[0] b[1] 0.00128f
C2213 _47_/a_299_297# net4 3.28e-19
C2214 _13_ _22_ 0.00309f
C2215 _34_/a_47_47# b[1] 0.0197f
C2216 _20_ _05_ 6.79e-19
C2217 net9 _04_ 0.0213f
C2218 net7 _09_ 0.00258f
C2219 _05_ b[1] 0.0316f
C2220 _20_ _42_/a_209_311# 1.66e-20
C2221 _29_/a_111_297# _06_ 6.74e-20
C2222 _11_ _15_ 0.113f
C2223 _38_/a_197_47# _10_ 6.29e-19
C2224 net6 _39_/a_377_297# 0.00143f
C2225 _42_/a_209_311# b[1] 5.21e-19
C2226 input2/a_27_47# _05_ 1.83e-19
C2227 net13 p[3] 9.49e-19
C2228 _12_ _00_ 0.00396f
C2229 _13_ _04_ 1.17e-21
C2230 input5/a_664_47# b[1] 0.00195f
C2231 VGND p[4] 0.366f
C2232 _27_/a_277_297# _03_ 2.1e-20
C2233 _50_/a_343_93# _15_ 0.0098f
C2234 net14 net6 2.82e-21
C2235 net14 net1 6.64e-20
C2236 _01_ input5/a_558_47# 3.97e-20
C2237 _52_/a_584_47# _22_ 6.24e-19
C2238 input2/a_27_47# _42_/a_209_311# 1e-22
C2239 _35_/a_226_47# _10_ 1.25e-19
C2240 _25_ net18 0.0594f
C2241 net12 _33_/a_209_311# 0.0769f
C2242 input5/a_558_47# net2 5.99e-21
C2243 _36_/a_27_47# net8 1.52e-19
C2244 input2/a_27_47# input5/a_664_47# 4.47e-21
C2245 _29_/a_183_297# VPWR -8.13e-19
C2246 _12_ _52_/a_93_21# 0.0157f
C2247 b[3] net19 0.054f
C2248 net8 _27_/a_27_297# 0.0108f
C2249 _32_/a_27_47# _43_/a_27_47# 2.01e-20
C2250 _22_ _00_ 0.477f
C2251 input13/a_27_47# VPWR 0.0696f
C2252 VGND _42_/a_368_53# -4.05e-19
C2253 net3 _19_ 0.0129f
C2254 _26_/a_183_297# _06_ 3.16e-19
C2255 _12_ b[2] 3.89e-20
C2256 _20_ _55_/a_80_21# 0.0291f
C2257 net7 _31_/a_35_297# 0.0384f
C2258 _16_ net7 7.5e-20
C2259 _04_ _52_/a_584_47# 2.5e-19
C2260 _42_/a_296_53# VPWR -6.37e-20
C2261 _32_/a_109_47# VPWR 0.00124f
C2262 _55_/a_80_21# b[1] 6.03e-19
C2263 _15_ _02_ 0.101f
C2264 _52_/a_93_21# _22_ 0.0347f
C2265 net5 output16/a_27_47# 4.14e-19
C2266 _53_/a_29_53# _12_ 3.46e-20
C2267 net17 _03_ 5.1e-19
C2268 VGND _55_/a_300_47# -0.00109f
C2269 _54_/a_75_212# net10 7.43e-19
C2270 _43_/a_27_47# _06_ 0.0329f
C2271 _18_ _43_/a_469_47# 1.59e-19
C2272 _04_ _00_ 1.98e-20
C2273 _06_ p[14] 1.04e-19
C2274 _20_ net10 3.23e-19
C2275 _14_ _49_/a_75_199# 6.79e-20
C2276 _53_/a_29_53# net16 2.04e-20
C2277 _22_ b[2] 0.0043f
C2278 net2 output17/a_27_47# 0.0285f
C2279 net11 _29_/a_183_297# 3.64e-19
C2280 VGND input12/a_27_47# 0.0405f
C2281 net10 b[1] 0.117f
C2282 VGND _27_/a_277_297# -4.65e-19
C2283 net8 net9 0.0605f
C2284 _27_/a_27_297# _42_/a_109_93# 1.35e-20
C2285 _53_/a_29_53# _22_ 0.00749f
C2286 output18/a_27_47# net18 0.0106f
C2287 _04_ _52_/a_93_21# 2.35e-19
C2288 _42_/a_209_311# _15_ 0.0521f
C2289 input2/a_27_47# net10 1.17e-20
C2290 input5/a_664_47# _15_ 9.15e-22
C2291 _32_/a_27_47# VPWR 0.0395f
C2292 _45_/a_109_297# _12_ 0.00587f
C2293 _36_/a_27_47# _18_ 5.46e-20
C2294 net5 _32_/a_197_47# 5.61e-21
C2295 _37_/a_27_47# _43_/a_193_413# 0.0102f
C2296 _43_/a_297_47# VGND -1.33e-19
C2297 net8 input7/a_27_47# 2.03e-21
C2298 net17 p[10] 0.179f
C2299 net1 _03_ 0.298f
C2300 net6 _03_ 2.9e-20
C2301 net16 _45_/a_109_297# 5.1e-20
C2302 _21_ _49_/a_75_199# 6.64e-19
C2303 _10_ _30_/a_297_297# 1.25e-20
C2304 _17_ _19_ 8.82e-21
C2305 _12_ _09_ 0.00526f
C2306 input3/a_27_47# output19/a_27_47# 4.77e-21
C2307 VGND input8/a_27_47# 0.0573f
C2308 net6 _50_/a_223_47# 0.0194f
C2309 _45_/a_109_297# _22_ 0.0426f
C2310 _06_ VPWR 1.4f
C2311 input5/a_558_47# _44_/a_93_21# 2.71e-19
C2312 net14 _20_ 8.01e-20
C2313 VGND net17 0.212f
C2314 _18_ _35_/a_76_199# 6.82e-21
C2315 _23_ _39_/a_47_47# 5.24e-21
C2316 net16 _09_ 0.00707f
C2317 _17_ _41_/a_59_75# 0.00149f
C2318 net14 b[1] 0.00256f
C2319 _15_ _55_/a_80_21# 0.107f
C2320 output19/a_27_47# _44_/a_250_297# 6.42e-20
C2321 net3 _01_ 1.16e-19
C2322 net12 _07_ 0.18f
C2323 _47_/a_299_297# VPWR 0.0643f
C2324 _18_ net9 1.51e-19
C2325 _22_ _09_ 0.0279f
C2326 _37_/a_27_47# input6/a_27_47# 9.35e-19
C2327 net1 p[10] 1.22e-19
C2328 _34_/a_129_47# _08_ 3.29e-19
C2329 net3 net2 0.519f
C2330 _18_ _45_/a_27_47# 0.00347f
C2331 input6/a_27_47# output19/a_27_47# 0.107f
C2332 input2/a_27_47# net14 0.0102f
C2333 input13/a_27_47# p[4] 7.37e-20
C2334 net14 _49_/a_201_297# 1.52e-19
C2335 net8 _00_ 3.23e-19
C2336 net11 _06_ 0.546f
C2337 _50_/a_27_47# _41_/a_59_75# 9.59e-22
C2338 p[5] b[1] 0.00702f
C2339 _29_/a_29_53# _49_/a_75_199# 1.28e-19
C2340 _21_ p[3] 5.54e-21
C2341 VGND net1 0.512f
C2342 _13_ _18_ 0.019f
C2343 VGND net6 0.472f
C2344 input9/a_75_212# _10_ 5.49e-21
C2345 _36_/a_197_47# _10_ 1.54e-19
C2346 net13 _36_/a_27_47# 0.0488f
C2347 _04_ _09_ 0.0904f
C2348 net8 input5/a_381_47# 7.48e-19
C2349 net5 _38_/a_27_47# 1.76e-19
C2350 output19/a_27_47# input14/a_27_47# 0.0101f
C2351 VGND _55_/a_472_297# -0.00188f
C2352 net5 _47_/a_384_47# 0.00129f
C2353 net8 _32_/a_303_47# 2.22e-34
C2354 net7 _22_ 2.73e-20
C2355 _54_/a_75_212# _03_ 5.45e-21
C2356 _16_ _22_ 3.8e-19
C2357 _12_ _47_/a_81_21# 0.00158f
C2358 input4/a_75_212# net5 0.0104f
C2359 _01_ _17_ 1.46e-20
C2360 net13 _35_/a_76_199# 0.0337f
C2361 net14 _15_ 0.225f
C2362 _24_ _07_ 5.67e-19
C2363 _10_ _41_/a_145_75# 5.18e-19
C2364 _33_/a_368_53# _08_ 5.04e-19
C2365 _20_ _03_ 0.0794f
C2366 _03_ b[1] 0.0738f
C2367 _36_/a_303_47# _25_ 2.03e-21
C2368 _17_ net2 0.181f
C2369 _18_ _00_ 0.157f
C2370 _34_/a_285_47# b[1] 0.00368f
C2371 input5/a_381_47# _42_/a_109_93# 0.00763f
C2372 _29_/a_29_53# p[3] 2.51e-19
C2373 net13 net9 0.035f
C2374 net6 p[12] 0.0941f
C2375 _30_/a_109_53# _02_ 5.03e-22
C2376 _26_/a_29_53# _36_/a_27_47# 1.6e-19
C2377 net7 _04_ 0.0602f
C2378 _20_ _50_/a_223_47# 1.71e-19
C2379 _45_/a_193_297# _00_ 4.38e-20
C2380 _04_ _31_/a_35_297# 1.89e-20
C2381 _08_ _02_ 2.26e-20
C2382 _22_ _47_/a_81_21# 7.25e-19
C2383 input2/a_27_47# _03_ 2.71e-19
C2384 p[13] net9 1.72e-19
C2385 _49_/a_201_297# _03_ 0.00842f
C2386 net5 _52_/a_346_47# 7.03e-19
C2387 _34_/a_47_47# _08_ 0.00123f
C2388 net3 _44_/a_93_21# 0.0102f
C2389 _21_ p[6] 0.00203f
C2390 _05_ _08_ 0.00897f
C2391 _05_ _30_/a_109_53# 0.033f
C2392 _39_/a_129_47# VPWR -9.47e-19
C2393 _18_ _52_/a_93_21# 1.97e-19
C2394 _10_ _52_/a_256_47# 1.65e-19
C2395 net13 _13_ 4e-21
C2396 _50_/a_429_93# net6 6.18e-19
C2397 _30_/a_392_297# b[1] 3.99e-19
C2398 _43_/a_193_413# _43_/a_369_47# -1.25e-19
C2399 _45_/a_193_297# _52_/a_93_21# 6.01e-19
C2400 p[10] b[1] 0.103f
C2401 _43_/a_469_47# _14_ 0.00259f
C2402 input10/a_27_47# net10 0.00321f
C2403 _54_/a_75_212# VGND 0.053f
C2404 _11_ _41_/a_59_75# 8.7e-19
C2405 _30_/a_215_297# p[3] 1.73e-19
C2406 _37_/a_27_47# p[14] 1.37e-19
C2407 output19/a_27_47# p[14] 0.0943f
C2408 VGND _20_ 0.471f
C2409 input2/a_27_47# p[10] 0.00905f
C2410 _26_/a_29_53# net9 0.00343f
C2411 net4 output16/a_27_47# 0.00706f
C2412 net5 input5/a_62_47# 0.00329f
C2413 _55_/a_300_47# _06_ 2.5e-20
C2414 VGND b[1] 0.557f
C2415 _50_/a_343_93# _41_/a_59_75# 6.13e-22
C2416 input12/a_27_47# _06_ 5.3e-22
C2417 net5 _39_/a_285_47# 0.05f
C2418 _30_/a_465_297# VPWR -4.57e-19
C2419 _01_ p[2] 0.00164f
C2420 _40_/a_109_297# _14_ -1.78e-33
C2421 input2/a_27_47# VGND -0.0137f
C2422 _15_ _03_ 7.39e-20
C2423 VGND _49_/a_201_297# -0.00403f
C2424 _27_/a_27_297# _14_ 1.66e-21
C2425 input13/a_27_47# net1 1.9e-19
C2426 _19_ _02_ 0.213f
C2427 _15_ _50_/a_223_47# 0.00698f
C2428 _17_ _44_/a_93_21# 0.0646f
C2429 net16 _12_ 0.131f
C2430 net15 _10_ 0.0101f
C2431 _33_/a_109_93# b[1] 0.00411f
C2432 net8 net7 0.295f
C2433 _43_/a_297_47# _06_ 4.81e-20
C2434 net8 _31_/a_35_297# 0.0408f
C2435 _16_ net8 0.00624f
C2436 net13 _52_/a_93_21# 7.21e-19
C2437 net10 _30_/a_109_53# 5.6e-20
C2438 net10 _08_ 0.194f
C2439 _37_/a_27_47# VPWR -0.0178f
C2440 _18_ _09_ 7.01e-21
C2441 _12_ _22_ 0.196f
C2442 output19/a_27_47# VPWR 0.0228f
C2443 _36_/a_27_47# _21_ 0.0276f
C2444 _45_/a_193_297# _09_ 0.00961f
C2445 _50_/a_515_93# VPWR -5.03e-19
C2446 p[13] input5/a_381_47# 0.00146f
C2447 _27_/a_27_297# net19 1.98e-19
C2448 _26_/a_29_53# _52_/a_584_47# 7.45e-20
C2449 net16 _22_ 0.00606f
C2450 input5/a_664_47# _19_ 2.19e-21
C2451 _35_/a_556_47# b[1] 3.23e-19
C2452 net8 _47_/a_81_21# 2.08e-21
C2453 _16_ input15/a_27_47# 7.13e-19
C2454 _12_ _04_ 1.42e-19
C2455 _26_/a_29_53# _00_ 0.0466f
C2456 input10/a_27_47# p[5] 0.0181f
C2457 _32_/a_27_47# net1 0.0211f
C2458 _11_ net2 0.234f
C2459 VGND _15_ 0.149f
C2460 _11_ _23_ 2e-20
C2461 _33_/a_209_311# VPWR -0.0131f
C2462 _36_/a_109_47# _04_ 2.39e-19
C2463 _02_ _52_/a_250_297# 0.0128f
C2464 _13_ _14_ 1.47e-20
C2465 net7 _31_/a_285_297# 0.00227f
C2466 _35_/a_76_199# _21_ 0.0175f
C2467 _50_/a_343_93# _01_ 0.0131f
C2468 _50_/a_343_93# net2 1.25e-20
C2469 _05_ _52_/a_250_297# 8.86e-22
C2470 _04_ _22_ 1.76e-20
C2471 _18_ net7 2.58e-20
C2472 _21_ net9 0.0282f
C2473 _48_/a_27_47# _02_ 0.00435f
C2474 net2 _37_/a_303_47# 4.41e-19
C2475 net1 _06_ 0.0115f
C2476 _36_/a_27_47# _29_/a_29_53# 6.92e-20
C2477 _21_ _45_/a_27_47# 1.18e-20
C2478 net6 _06_ 0.307f
C2479 _48_/a_27_47# _34_/a_47_47# 4.45e-21
C2480 _16_ _18_ 0.144f
C2481 _33_/a_209_311# net11 2.49e-19
C2482 _45_/a_465_47# VGND -8.14e-19
C2483 _38_/a_27_47# net4 0.0119f
C2484 _47_/a_299_297# net6 3.63e-19
C2485 _13_ _21_ 1.69e-19
C2486 net13 _09_ 0.0379f
C2487 _01_ _02_ 0.106f
C2488 _18_ _47_/a_81_21# 7.96e-20
C2489 _23_ _02_ 0.0648f
C2490 input3/a_27_47# b[3] 1.4e-19
C2491 _15_ p[12] 0.0163f
C2492 input13/a_27_47# b[1] 0.00624f
C2493 input5/a_62_47# p[11] 0.00153f
C2494 _01_ _05_ 5.03e-19
C2495 _29_/a_29_53# _35_/a_76_199# 9.88e-19
C2496 _14_ _00_ 0.133f
C2497 _38_/a_303_47# _10_ 7.36e-19
C2498 input4/a_75_212# net4 0.0189f
C2499 _42_/a_296_53# b[1] 2.38e-20
C2500 net2 _05_ 4.03e-20
C2501 _44_/a_250_297# b[3] 3.33e-19
C2502 _01_ _42_/a_209_311# 1.58e-19
C2503 _29_/a_29_53# net9 0.0205f
C2504 VPWR output16/a_27_47# 0.122f
C2505 _36_/a_27_47# _30_/a_215_297# 7.13e-20
C2506 _50_/a_429_93# _15_ 6.82e-19
C2507 input3/a_27_47# input5/a_62_47# 0.00179f
C2508 input5/a_381_47# _14_ 5.68e-20
C2509 net2 _42_/a_209_311# 5.1e-19
C2510 net3 _27_/a_109_297# 5.45e-19
C2511 _35_/a_489_413# _10_ 3.41e-19
C2512 input6/a_27_47# b[3] 0.00217f
C2513 p[7] net13 0.00514f
C2514 input5/a_664_47# net2 8.11e-20
C2515 _11_ _44_/a_93_21# 4.78e-20
C2516 _21_ _00_ 9.26e-20
C2517 input5/a_62_47# _44_/a_250_297# 2.45e-20
C2518 net14 _19_ 0.0512f
C2519 net10 _52_/a_250_297# 2.86e-21
C2520 net13 net7 1.72e-19
C2521 _11_ _25_ 7.05e-19
C2522 net15 input5/a_558_47# 0.00672f
C2523 _32_/a_27_47# _20_ 0.0069f
C2524 net7 _31_/a_117_297# 0.00472f
C2525 net8 _22_ 3.3e-20
C2526 _03_ _30_/a_109_53# 0.0189f
C2527 _32_/a_27_47# b[1] 6.39e-19
C2528 _03_ _08_ 0.0144f
C2529 _34_/a_285_47# _08_ 0.00414f
C2530 _07_ VPWR 0.0728f
C2531 net13 _31_/a_35_297# 1.86e-20
C2532 input10/a_27_47# VGND 0.00285f
C2533 p[13] net7 1.91e-19
C2534 _32_/a_197_47# VPWR 0.00146f
C2535 _43_/a_369_47# VPWR -3.75e-19
C2536 _37_/a_109_47# VPWR -4.38e-19
C2537 _48_/a_27_47# net10 0.00377f
C2538 b[3] input14/a_27_47# 0.00296f
C2539 input5/a_381_47# net19 0.00173f
C2540 _54_/a_75_212# _06_ 0.00727f
C2541 _01_ _55_/a_80_21# 0.0121f
C2542 _21_ _52_/a_93_21# 9.4e-19
C2543 _30_/a_215_297# net9 0.0456f
C2544 _20_ _06_ 0.133f
C2545 _21_ b[2] 2.14e-19
C2546 _06_ b[1] 0.0885f
C2547 net8 _04_ 0.02f
C2548 net12 p[6] 0.0256f
C2549 _42_/a_296_53# _15_ 1.28e-19
C2550 _53_/a_29_53# _21_ 0.00959f
C2551 net2 net10 2.05e-20
C2552 _42_/a_109_93# _22_ 1.21e-19
C2553 net11 _07_ 0.0206f
C2554 _47_/a_299_297# _20_ 0.002f
C2555 net4 _39_/a_285_47# 9.71e-19
C2556 _18_ _12_ 0.0115f
C2557 net6 _39_/a_129_47# 6.91e-19
C2558 _23_ net10 0.00216f
C2559 _25_ _02_ 0.0156f
C2560 _45_/a_193_297# _12_ 0.0103f
C2561 _18_ net16 8.17e-21
C2562 _25_ _34_/a_47_47# 1.08e-19
C2563 VGND _30_/a_109_53# -0.0072f
C2564 net16 _45_/a_193_297# 0.00187f
C2565 VGND _08_ 0.161f
C2566 _18_ _22_ 0.0211f
C2567 _42_/a_209_311# _44_/a_93_21# 2.21e-19
C2568 _04_ _42_/a_109_93# 5.77e-22
C2569 _45_/a_193_297# _22_ 0.0234f
C2570 input5/a_664_47# _44_/a_93_21# 1.88e-20
C2571 _19_ _03_ 0.0019f
C2572 _32_/a_27_47# _15_ 1.19e-19
C2573 _36_/a_27_47# net5 0.0163f
C2574 _38_/a_27_47# VPWR -0.0142f
C2575 net14 _01_ 8.29e-19
C2576 net5 _27_/a_27_297# 3.48e-19
C2577 _47_/a_384_47# VPWR -1.45e-19
C2578 _35_/a_226_47# _02_ 2.21e-19
C2579 net15 _39_/a_47_47# 9.44e-22
C2580 _18_ _04_ 1.94e-21
C2581 _21_ _09_ 0.263f
C2582 net14 net2 0.151f
C2583 output18/a_27_47# _02_ 4.13e-19
C2584 b[3] p[14] 0.0976f
C2585 _28_/a_109_297# net9 3.7e-19
C2586 _35_/a_226_47# _05_ 0.0134f
C2587 _15_ _06_ 0.22f
C2588 net7 _14_ 0.00251f
C2589 net3 net15 0.394f
C2590 input4/a_75_212# VPWR 0.06f
C2591 _19_ p[10] 9.65e-20
C2592 _33_/a_209_311# net17 7.03e-21
C2593 _49_/a_208_47# _02_ 0.00193f
C2594 net13 _12_ 0.00632f
C2595 _16_ _14_ 0.0584f
C2596 _37_/a_27_47# net6 4.3e-20
C2597 net5 _35_/a_76_199# 3.38e-19
C2598 _36_/a_303_47# _10_ 4.09e-19
C2599 _38_/a_27_47# net11 1.68e-20
C2600 output19/a_27_47# net6 0.00112f
C2601 input9/a_75_212# p[2] 5.13e-20
C2602 net12 _36_/a_27_47# 0.0177f
C2603 net13 _36_/a_109_47# 0.00126f
C2604 _47_/a_299_297# _15_ 0.0103f
C2605 net5 net9 0.0368f
C2606 _35_/a_556_47# _08_ 7.71e-19
C2607 _50_/a_515_93# net6 4.7e-19
C2608 _10_ _39_/a_47_47# 0.00824f
C2609 net5 _45_/a_27_47# 0.0288f
C2610 VGND _19_ 0.379f
C2611 net13 _22_ 4.63e-20
C2612 _25_ net10 2.66e-19
C2613 _14_ _47_/a_81_21# 6.24e-20
C2614 _20_ _39_/a_129_47# 1.71e-20
C2615 _52_/a_346_47# VPWR -0.00109f
C2616 _29_/a_29_53# _09_ 0.00488f
C2617 _21_ net7 3e-19
C2618 _48_/a_27_47# _34_/a_285_47# 6.66e-20
C2619 net3 _10_ 3.89e-19
C2620 _13_ net5 0.0381f
C2621 VGND _41_/a_59_75# 0.0138f
C2622 _49_/a_315_47# p[2] 6.65e-20
C2623 _16_ net19 0.206f
C2624 b[3] VPWR 0.129f
C2625 net12 _35_/a_76_199# 0.0132f
C2626 net8 _31_/a_285_297# 0.0215f
C2627 _26_/a_29_53# _12_ 0.00243f
C2628 _01_ _03_ 2.85e-19
C2629 net12 net9 0.0596f
C2630 net13 _04_ 0.569f
C2631 net15 input5/a_841_47# 0.00585f
C2632 input5/a_62_47# VPWR 0.0601f
C2633 _18_ net8 1.15e-21
C2634 net2 _03_ 1.89e-19
C2635 net15 _17_ 0.195f
C2636 _23_ _03_ 0.0564f
C2637 _35_/a_226_47# net10 0.018f
C2638 net5 _52_/a_584_47# 0.0022f
C2639 net14 _44_/a_93_21# 0.0646f
C2640 VGND _52_/a_250_297# -0.00314f
C2641 _39_/a_285_47# VPWR -9.53e-19
C2642 _26_/a_29_53# _22_ 0.09f
C2643 _30_/a_465_297# b[1] 4.8e-19
C2644 _29_/a_29_53# net7 6.01e-19
C2645 net5 _00_ 0.00954f
C2646 _18_ input15/a_27_47# 8.27e-21
C2647 _48_/a_27_47# VGND 0.0548f
C2648 p[12] _41_/a_59_75# 0.0547f
C2649 input1/a_75_212# VPWR 0.0786f
C2650 net2 p[10] 0.0334f
C2651 _17_ _10_ 0.0233f
C2652 net5 input5/a_381_47# 0.0546f
C2653 _26_/a_29_53# _04_ 2.3e-21
C2654 _33_/a_109_93# _52_/a_250_297# 5.17e-22
C2655 net6 output16/a_27_47# 1.5e-19
C2656 net5 _52_/a_93_21# 0.0124f
C2657 VPWR _49_/a_75_199# 0.0154f
C2658 _01_ VGND 0.0939f
C2659 _12_ _14_ 1.98e-20
C2660 net5 b[2] 7.33e-20
C2661 net5 _32_/a_303_47# 7.18e-21
C2662 _14_ _40_/a_297_297# 1.58e-19
C2663 _40_/a_191_297# _14_ 2.4e-19
C2664 VGND net2 0.848f
C2665 VGND _23_ 0.16f
C2666 p[12] _52_/a_250_297# 1.84e-20
C2667 input9/a_75_212# _05_ 1.24e-21
C2668 _32_/a_27_47# _30_/a_109_53# 1.51e-19
C2669 _24_ _45_/a_27_47# 4.57e-19
C2670 _10_ _50_/a_27_47# 0.0154f
C2671 net13 net8 7.51e-20
C2672 _30_/a_215_297# _31_/a_35_297# 6.37e-19
C2673 net1 _07_ 6.08e-22
C2674 _14_ _22_ 0.00449f
C2675 _33_/a_209_311# b[1] 0.0129f
C2676 _49_/a_315_47# _02_ 0.00134f
C2677 net1 _32_/a_197_47# 0.00142f
C2678 net6 _43_/a_369_47# 3.62e-21
C2679 _13_ _24_ 2.47e-19
C2680 p[1] input1/a_75_212# 0.0023f
C2681 _06_ _30_/a_109_53# 1.96e-19
C2682 net8 _31_/a_117_297# 5.91e-19
C2683 net11 _49_/a_75_199# 4.49e-19
C2684 net10 _30_/a_297_297# 1.68e-19
C2685 p[13] net8 0.00353f
C2686 _06_ _08_ 0.0343f
C2687 p[13] p[8] 0.00255f
C2688 _12_ _21_ 7.99e-20
C2689 _25_ _03_ 0.00422f
C2690 _50_/a_615_93# VPWR -5.34e-19
C2691 net16 _21_ 1.89e-19
C2692 net5 _45_/a_109_297# 0.0184f
C2693 p[3] VPWR 0.0867f
C2694 _04_ _14_ 2.04e-21
C2695 _36_/a_27_47# net4 0.0103f
C2696 net3 input5/a_558_47# 0.0137f
C2697 _22_ net19 2.17e-19
C2698 _21_ _22_ 0.00314f
C2699 _26_/a_111_297# _00_ 3.7e-19
C2700 _13_ _43_/a_193_413# 5.58e-21
C2701 _37_/a_27_47# _15_ 1.11e-19
C2702 net5 _09_ 5.18e-19
C2703 net13 _31_/a_285_297# 3.85e-20
C2704 _02_ _52_/a_256_47# 0.00344f
C2705 net7 _31_/a_285_47# 0.00132f
C2706 _50_/a_515_93# _15_ 0.00147f
C2707 net15 _11_ 0.145f
C2708 b[0] _39_/a_47_47# 2.04e-19
C2709 _35_/a_226_47# _03_ 0.028f
C2710 _53_/a_111_297# _10_ 2.06e-19
C2711 net13 _18_ 1.06e-20
C2712 _04_ net19 2.07e-20
C2713 input9/a_75_212# net10 0.00699f
C2714 _21_ _04_ 0.39f
C2715 p[8] p[9] 0.00347f
C2716 VGND _44_/a_93_21# -0.0223f
C2717 net3 output17/a_27_47# 0.00248f
C2718 net4 net9 1.99e-22
C2719 net15 _37_/a_303_47# 0.00118f
C2720 _24_ _52_/a_93_21# 0.0211f
C2721 VGND _25_ 0.199f
C2722 p[1] p[3] 7.76e-20
C2723 _38_/a_109_47# net4 7.32e-19
C2724 _45_/a_27_47# net4 0.024f
C2725 _49_/a_208_47# _03_ 3.86e-19
C2726 _29_/a_29_53# _22_ 2.24e-21
C2727 net12 _09_ 0.0374f
C2728 _16_ _28_/a_109_297# 1.26e-19
C2729 _24_ b[2] 1.85e-19
C2730 _43_/a_193_413# _00_ 0.00721f
C2731 _11_ _10_ 0.176f
C2732 input15/a_27_47# p[9] 0.0192f
C2733 p[6] VPWR 0.0732f
C2734 _20_ _07_ 1.28e-21
C2735 net5 net7 0.195f
C2736 _53_/a_29_53# _24_ 0.0835f
C2737 VGND _38_/a_197_47# 2.29e-19
C2738 _06_ _41_/a_59_75# 0.0429f
C2739 net5 _31_/a_35_297# 2.04e-21
C2740 input5/a_558_47# _17_ 2.13e-21
C2741 _16_ net5 1.99e-20
C2742 _13_ net4 0.212f
C2743 input4/a_75_212# net6 0.0273f
C2744 _07_ b[1] 0.0417f
C2745 net15 _02_ 0.0806f
C2746 _50_/a_343_93# _10_ 0.0284f
C2747 net8 _14_ 4.23e-19
C2748 _26_/a_29_53# _18_ 5.26e-20
C2749 _01_ _32_/a_109_47# 0.00129f
C2750 _29_/a_111_297# net9 8.06e-21
C2751 _29_/a_29_53# _04_ 0.0408f
C2752 _44_/a_250_297# _00_ 6.39e-20
C2753 VGND _35_/a_226_47# -0.0111f
C2754 _47_/a_299_297# _41_/a_59_75# 0.00146f
C2755 net14 _27_/a_109_297# 1.32e-19
C2756 net3 _27_/a_205_297# 4.37e-19
C2757 net3 _39_/a_47_47# 1.66e-20
C2758 net5 _47_/a_81_21# 4.59e-19
C2759 net11 p[6] 0.0099f
C2760 p[7] net12 0.0313f
C2761 input15/a_27_47# _14_ 9.48e-21
C2762 VGND output18/a_27_47# 0.0581f
C2763 _30_/a_215_297# _22_ 2.46e-21
C2764 net10 _52_/a_256_47# 8.13e-20
C2765 net15 _42_/a_209_311# 0.0157f
C2766 _06_ _52_/a_250_297# 0.0058f
C2767 net12 net7 1.57e-19
C2768 net15 input5/a_664_47# 0.0216f
C2769 _03_ _30_/a_297_297# 0.00117f
C2770 _49_/a_208_47# VGND -0.00164f
C2771 _10_ _02_ 0.0537f
C2772 net8 net19 1.15e-19
C2773 _21_ net8 0.00656f
C2774 p[8] net19 1.25e-19
C2775 _42_/a_109_93# _14_ 0.00141f
C2776 _37_/a_197_47# VPWR -3.27e-19
C2777 net6 b[3] 0.00152f
C2778 _32_/a_27_47# _01_ 0.0266f
C2779 _33_/a_109_93# _35_/a_226_47# 4.9e-19
C2780 _48_/a_27_47# _06_ 0.0251f
C2781 _43_/a_469_47# VPWR -2.75e-19
C2782 _24_ _09_ 0.0202f
C2783 net4 _00_ 0.0166f
C2784 _10_ _05_ 9.25e-21
C2785 _30_/a_215_297# _04_ 0.00225f
C2786 input15/a_27_47# net19 0.00236f
C2787 input8/a_27_47# _49_/a_75_199# 1.99e-20
C2788 net1 input5/a_62_47# 7.59e-20
C2789 _18_ _14_ 0.243f
C2790 net4 _52_/a_93_21# 7.93e-20
C2791 _54_/a_75_212# _38_/a_27_47# 2.67e-19
C2792 _36_/a_27_47# VPWR -0.00832f
C2793 _01_ _06_ 0.00157f
C2794 net17 _49_/a_75_199# 0.00127f
C2795 _40_/a_109_297# VPWR -4.23e-19
C2796 net15 _55_/a_80_21# 0.00759f
C2797 net6 _39_/a_285_47# 1.53e-19
C2798 net13 _26_/a_29_53# 2.23e-20
C2799 net2 _06_ 0.0108f
C2800 _47_/a_384_47# _20_ 1.72e-19
C2801 _23_ _06_ 0.218f
C2802 _42_/a_109_93# net19 0.0448f
C2803 _27_/a_27_297# VPWR 0.0329f
C2804 net18 _02_ 8.53e-20
C2805 _17_ _39_/a_47_47# 1.47e-20
C2806 _13_ _43_/a_27_47# 1.66e-20
C2807 _53_/a_29_53# net4 3.26e-19
C2808 input9/a_75_212# _03_ 9.32e-20
C2809 net1 input1/a_75_212# 0.00208f
C2810 p[4] p[6] 0.0051f
C2811 VGND _30_/a_297_297# -5.13e-19
C2812 _47_/a_299_297# net2 1.18e-19
C2813 _44_/a_584_47# VPWR -2.28e-19
C2814 _27_/a_109_297# _03_ 1.97e-20
C2815 _18_ net19 4.89e-20
C2816 _35_/a_76_199# VPWR -0.00947f
C2817 net3 _17_ 0.0698f
C2818 _36_/a_27_47# net11 0.0707f
C2819 _10_ _55_/a_80_21# 5.49e-19
C2820 net5 _12_ 0.983f
C2821 net1 _49_/a_75_199# 0.00799f
C2822 _36_/a_109_47# net5 0.00144f
C2823 _27_/a_27_297# net11 1.58e-20
C2824 _26_/a_183_297# _00_ 4.53e-19
C2825 net9 VPWR 0.496f
C2826 p[3] input8/a_27_47# 0.0023f
C2827 _49_/a_315_47# _03_ 9.22e-19
C2828 _45_/a_27_47# VPWR -0.00418f
C2829 _45_/a_109_297# net4 6.43e-20
C2830 _38_/a_109_47# VPWR -4.66e-19
C2831 net5 net16 0.00476f
C2832 _35_/a_489_413# _02_ 3.86e-19
C2833 _10_ net10 4.45e-19
C2834 _33_/a_209_311# _08_ 0.0122f
C2835 _16_ p[11] 4e-20
C2836 _52_/a_346_47# b[1] 6.37e-20
C2837 _43_/a_193_413# net7 3.49e-19
C2838 net5 _22_ 0.405f
C2839 p[1] _27_/a_27_297# 2.35e-19
C2840 _30_/a_215_297# net8 8.14e-21
C2841 _43_/a_27_47# _00_ 0.0431f
C2842 _16_ _43_/a_193_413# 0.0261f
C2843 input13/a_27_47# _35_/a_226_47# 3.94e-20
C2844 _35_/a_76_199# net11 4e-19
C2845 net14 net15 1.07f
C2846 net4 _09_ 0.00262f
C2847 _13_ VPWR 0.0804f
C2848 input7/a_27_47# VPWR 0.0768f
C2849 _33_/a_296_53# _05_ 4.53e-19
C2850 p[6] input12/a_27_47# 0.017f
C2851 input9/a_75_212# VGND 0.063f
C2852 net12 _12_ 7.94e-21
C2853 _36_/a_197_47# VGND -3.75e-19
C2854 VGND _27_/a_109_297# -6.15e-19
C2855 net11 net9 0.136f
C2856 _34_/a_377_297# net10 1.62e-19
C2857 net5 _04_ 0.00476f
C2858 _50_/a_615_93# net6 1.43e-19
C2859 _45_/a_27_47# net11 3.64e-20
C2860 _47_/a_384_47# _15_ 0.00112f
C2861 _16_ _44_/a_250_297# 3.25e-19
C2862 _10_ _39_/a_377_297# 7.42e-19
C2863 net1 p[3] 6.54e-19
C2864 input5/a_62_47# b[1] 0.0024f
C2865 net18 net10 3.35e-20
C2866 _25_ _06_ 0.144f
C2867 net13 _21_ 0.13f
C2868 net12 _22_ 5.73e-20
C2869 _29_/a_111_297# _09_ 5.79e-20
C2870 _13_ net11 2.34e-19
C2871 _52_/a_584_47# VPWR -9.47e-19
C2872 _49_/a_315_47# VGND -0.0034f
C2873 net14 _10_ 2.4e-19
C2874 VGND _41_/a_145_75# 3.75e-19
C2875 _26_/a_29_53# _14_ 3.67e-19
C2876 VPWR _00_ 0.416f
C2877 _38_/a_197_47# _06_ 4.32e-19
C2878 net8 _31_/a_285_47# 0.00129f
C2879 p[1] input7/a_27_47# 0.0168f
C2880 input1/a_75_212# b[1] 0.0074f
C2881 _49_/a_544_297# _09_ 2.56e-20
C2882 net12 _04_ 0.267f
C2883 _16_ net4 2.73e-20
C2884 _17_ _50_/a_27_47# 3.93e-20
C2885 input5/a_558_47# _42_/a_209_311# 7.85e-20
C2886 net7 _55_/a_217_297# 1.04e-19
C2887 _13_ _45_/a_205_47# 7.51e-20
C2888 input5/a_381_47# VPWR 8.33e-19
C2889 _20_ _49_/a_75_199# 0.0233f
C2890 _35_/a_226_47# _06_ 0.00487f
C2891 _35_/a_489_413# net10 0.00225f
C2892 _14_ p[9] 2.62e-21
C2893 _52_/a_93_21# VPWR -0.00838f
C2894 _49_/a_75_199# b[1] 0.00805f
C2895 _11_ _39_/a_47_47# 3.9e-19
C2896 _16_ _55_/a_217_297# 0.0017f
C2897 _24_ _12_ 1.67e-19
C2898 VGND _52_/a_256_47# -0.00161f
C2899 _33_/a_296_53# net10 8.22e-20
C2900 _32_/a_303_47# VPWR 6.03e-19
C2901 VPWR b[2] 0.262f
C2902 _15_ b[3] 1.89e-19
C2903 p[0] output17/a_27_47# 0.00805f
C2904 net15 _03_ 4.26e-20
C2905 net13 _29_/a_29_53# 0.00104f
C2906 output18/a_27_47# _06_ 0.0114f
C2907 _26_/a_111_297# _22_ 0.00137f
C2908 net16 _24_ 6.93e-19
C2909 output17/a_27_47# _05_ 1.12e-19
C2910 _07_ _08_ 0.348f
C2911 _53_/a_29_53# VPWR 0.00821f
C2912 p[12] _41_/a_145_75# 0.00339f
C2913 net1 p[6] 3.12e-20
C2914 net3 _11_ 0.165f
C2915 net5 net8 0.48f
C2916 _24_ _22_ 0.0846f
C2917 net11 _52_/a_93_21# 2.8e-19
C2918 net19 p[9] 0.0731f
C2919 _49_/a_544_297# net7 2.72e-19
C2920 _43_/a_193_413# _12_ 7.94e-22
C2921 net18 p[5] 1.98e-19
C2922 net11 b[2] 1.46e-19
C2923 net3 _37_/a_303_47# 0.00133f
C2924 _50_/a_615_93# _20_ 8.8e-19
C2925 net15 p[10] 0.00989f
C2926 p[11] _22_ 3.13e-20
C2927 _44_/a_256_47# _14_ 0.00124f
C2928 _10_ _03_ 0.00244f
C2929 _45_/a_109_297# VPWR -0.011f
C2930 p[3] b[1] 0.00382f
C2931 _53_/a_29_53# net11 8.31e-19
C2932 _37_/a_27_47# net2 0.0692f
C2933 _39_/a_47_47# _02_ 0.0127f
C2934 output19/a_27_47# net2 0.00168f
C2935 _26_/a_29_53# _29_/a_29_53# 0.00121f
C2936 net13 _30_/a_215_297# 0.0246f
C2937 _43_/a_193_413# _22_ 0.00133f
C2938 _10_ _50_/a_223_47# 0.0295f
C2939 input9/a_75_212# input13/a_27_47# 0.00732f
C2940 net15 VGND 0.222f
C2941 net5 _42_/a_109_93# 0.00109f
C2942 input3/a_27_47# _22_ 5.13e-20
C2943 net12 net8 0.00458f
C2944 _14_ net19 0.00714f
C2945 _34_/a_377_297# _03_ 3.13e-20
C2946 _27_/a_27_297# net17 0.00181f
C2947 net3 _02_ 9.52e-20
C2948 net7 _43_/a_27_47# 6.31e-19
C2949 net6 _43_/a_469_47# 4.85e-21
C2950 VPWR _09_ 0.297f
C2951 _16_ _43_/a_27_47# 2.47e-19
C2952 _11_ _17_ 0.197f
C2953 _43_/a_193_413# _04_ 5.67e-21
C2954 _45_/a_109_297# net11 7.46e-20
C2955 net18 _03_ 2.07e-21
C2956 net5 _18_ 0.0426f
C2957 output17/a_27_47# net10 1.31e-20
C2958 input3/a_27_47# _04_ 3.55e-19
C2959 net5 _45_/a_193_297# 0.00935f
C2960 _50_/a_343_93# _17_ 0.0015f
C2961 net3 _42_/a_209_311# 0.029f
C2962 _12_ net4 0.105f
C2963 _04_ 0 0.341f
C2964 net9 0 0.285f
C2965 _03_ 0 0.36f
C2966 net10 0 0.422f
C2967 _30_/a_109_53# 0 0.159f
C2968 _30_/a_215_297# 0 0.142f
C2969 _05_ 0 0.152f
C2970 net8 0 0.394f
C2971 _31_/a_285_297# 0 0.00137f
C2972 _31_/a_35_297# 0 0.255f
C2973 _06_ 0 0.79f
C2974 _32_/a_27_47# 0 0.175f
C2975 _11_ 0 0.267f
C2976 _50_/a_343_93# 0 0.172f
C2977 _50_/a_223_47# 0 0.141f
C2978 _50_/a_27_47# 0 0.259f
C2979 _07_ 0 0.288f
C2980 _33_/a_209_311# 0 0.143f
C2981 _33_/a_109_93# 0 0.158f
C2982 _08_ 0 0.131f
C2983 _34_/a_285_47# 0 0.0174f
C2984 _34_/a_47_47# 0 0.199f
C2985 _23_ 0 0.106f
C2986 _09_ 0 0.142f
C2987 _35_/a_489_413# 0 0.0254f
C2988 _35_/a_226_47# 0 0.162f
C2989 _35_/a_76_199# 0 0.141f
C2990 p[9] 0 0.241f
C2991 input15/a_27_47# 0 0.208f
C2992 _24_ 0 0.135f
C2993 _12_ 0 0.387f
C2994 _52_/a_250_297# 0 0.0278f
C2995 _52_/a_93_21# 0 0.151f
C2996 _10_ 0 0.643f
C2997 _36_/a_27_47# 0 0.175f
C2998 _53_/a_29_53# 0 0.18f
C2999 p[8] 0 0.33f
C3000 input14/a_27_47# 0 0.208f
C3001 _37_/a_27_47# 0 0.175f
C3002 p[7] 0 0.227f
C3003 input13/a_27_47# 0 0.208f
C3004 net18 0 0.207f
C3005 _25_ 0 0.191f
C3006 _54_/a_75_212# 0 0.21f
C3007 _38_/a_27_47# 0 0.175f
C3008 net19 0 0.187f
C3009 _22_ 0 0.215f
C3010 _14_ 0 0.228f
C3011 _15_ 0 0.336f
C3012 _55_/a_217_297# 0 0.00117f
C3013 _55_/a_80_21# 0 0.21f
C3014 p[6] 0 0.207f
C3015 input12/a_27_47# 0 0.208f
C3016 p[3] 0 0.236f
C3017 input9/a_75_212# 0 0.21f
C3018 _39_/a_285_47# 0 0.0174f
C3019 _39_/a_47_47# 0 0.199f
C3020 p[5] 0 0.267f
C3021 input11/a_27_47# 0 0.208f
C3022 p[2] 0 0.218f
C3023 input8/a_27_47# 0 0.208f
C3024 p[4] 0 0.327f
C3025 input10/a_27_47# 0 0.208f
C3026 net7 0 0.463f
C3027 p[1] 0 0.22f
C3028 input7/a_27_47# 0 0.208f
C3029 p[14] 0 0.24f
C3030 input6/a_27_47# 0 0.208f
C3031 net5 0 0.824f
C3032 p[13] 0 0.394f
C3033 input5/a_841_47# 0 0.0929f
C3034 input5/a_664_47# 0 0.13f
C3035 input5/a_558_47# 0 0.164f
C3036 input5/a_381_47# 0 0.11f
C3037 input5/a_62_47# 0 0.169f
C3038 p[12] 0 0.36f
C3039 input4/a_75_212# 0 0.21f
C3040 p[11] 0 0.248f
C3041 input3/a_27_47# 0 0.208f
C3042 net2 0 0.825f
C3043 p[10] 0 0.278f
C3044 input2/a_27_47# 0 0.208f
C3045 net1 0 0.342f
C3046 p[0] 0 0.312f
C3047 input1/a_75_212# 0 0.21f
C3048 b[3] 0 0.247f
C3049 output19/a_27_47# 0 0.543f
C3050 b[2] 0 0.515f
C3051 output18/a_27_47# 0 0.543f
C3052 b[1] 0 0.39f
C3053 net17 0 0.172f
C3054 output17/a_27_47# 0 0.543f
C3055 _41_/a_59_75# 0 0.177f
C3056 b[0] 0 0.528f
C3057 output16/a_27_47# 0 0.543f
C3058 _16_ 0 0.125f
C3059 _42_/a_209_311# 0 0.143f
C3060 _42_/a_109_93# 0 0.158f
C3061 _17_ 0 0.251f
C3062 _43_/a_193_413# 0 0.136f
C3063 _43_/a_27_47# 0 0.224f
C3064 net6 0 0.531f
C3065 net4 0 0.324f
C3066 _26_/a_29_53# 0 0.18f
C3067 _01_ 0 0.15f
C3068 net14 0 0.516f
C3069 net3 0 0.464f
C3070 net15 0 0.452f
C3071 _27_/a_27_297# 0 0.163f
C3072 _18_ 0 0.143f
C3073 _44_/a_250_297# 0 0.0278f
C3074 _44_/a_93_21# 0 0.151f
C3075 net16 0 0.231f
C3076 _13_ 0 0.133f
C3077 _45_/a_193_297# 0 0.0011f
C3078 _45_/a_109_297# 0 7.11e-19
C3079 _45_/a_27_47# 0 0.216f
C3080 _00_ 0 0.377f
C3081 net11 0 0.775f
C3082 net12 0 0.531f
C3083 net13 0 0.382f
C3084 _29_/a_29_53# 0 0.18f
C3085 _19_ 0 0.118f
C3086 _47_/a_299_297# 0 0.0348f
C3087 _47_/a_81_21# 0 0.147f
C3088 VPWR 0 40.3f
C3089 VGND 0 13.7f
C3090 _48_/a_27_47# 0 0.177f
C3091 _21_ 0 0.29f
C3092 _20_ 0 0.238f
C3093 _02_ 0 0.45f
C3094 _49_/a_201_297# 0 0.00345f
C3095 _49_/a_75_199# 0 0.205f
.ends

