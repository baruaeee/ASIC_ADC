magic
tech sky130A
timestamp 1706270542
<< pwell >>
rect -243 -126 243 126
<< nmos >>
rect -145 -21 145 21
<< ndiff >>
rect -174 15 -145 21
rect -174 -15 -168 15
rect -151 -15 -145 15
rect -174 -21 -145 -15
rect 145 15 174 21
rect 145 -15 151 15
rect 168 -15 174 15
rect 145 -21 174 -15
<< ndiffc >>
rect -168 -15 -151 15
rect 151 -15 168 15
<< psubdiff >>
rect -225 60 -208 91
rect -225 -91 -208 -60
<< psubdiffcont >>
rect -225 -60 -208 60
<< poly >>
rect -145 57 145 65
rect -145 40 -137 57
rect 137 40 145 57
rect -145 21 145 40
rect -145 -40 145 -21
rect -145 -57 -137 -40
rect 137 -57 145 -40
rect -145 -65 145 -57
<< polycont >>
rect -137 40 137 57
rect -137 -57 137 -40
<< locali >>
rect -225 60 -208 91
rect -145 40 -137 57
rect 137 40 145 57
rect -168 15 -151 23
rect -168 -23 -151 -15
rect 151 15 168 23
rect 151 -23 168 -15
rect -145 -57 -137 -40
rect 137 -57 145 -40
rect -225 -91 -208 -60
<< viali >>
rect -137 40 137 57
rect -168 -15 -151 15
rect 151 -15 168 15
rect -137 -57 137 -40
<< metal1 >>
rect -143 57 143 60
rect -143 40 -137 57
rect 137 40 143 57
rect -143 37 143 40
rect -171 15 -148 21
rect -171 -15 -168 15
rect -151 -15 -148 15
rect -171 -21 -148 -15
rect 148 15 171 21
rect 148 -15 151 15
rect 168 -15 171 15
rect 148 -21 171 -15
rect -143 -40 143 -37
rect -143 -57 -137 -40
rect 137 -57 143 -40
rect -143 -60 143 -57
<< properties >>
string FIXED_BBOX -216 -99 216 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 2.9 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
