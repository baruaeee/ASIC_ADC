** sch_path: /home/exotic/Desktop/ASIC_ADC/xschem/Vth_sch/Pre_layout/th06.sch
**.subckt th06 Vin Vout
*.ipin Vin
*.opin Vout
VDD VDD GND 1.8
Vin Vin GND pulse(0 0.2 0ns 1ns 1ns 5ns 10ns)
V_logic_high V_LH GND 1.25
V_logic_low V_LL GND 0.5
x1 VDD Vin Vout GND th06
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.save all





.dc Vin 0 1.8 0.01
*.tran 1n 30n
.control
run
set color0=white
set color1=black
plot Vin Vout V_LH V_LL
set xbrushwidth=3
.save all
.endc
.end


**** end user architecture code
**.ends

* NGSPICE file created from th06.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_L7T3GD a_n33_n130# a_15_n42# a_n175_n216# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n42# a_n33_n130# 0.0209f
C1 a_n33_n130# a_15_n42# 0.0209f
C2 a_n73_n42# a_15_n42# 0.0699f
C3 a_15_n42# a_n175_n216# 0.0729f
C4 a_n73_n42# a_n175_n216# 0.0729f
C5 a_n33_n130# a_n175_n216# 0.338f
.ends

.subckt sky130_fd_pr__pfet_01v8_NZD9V2 w_n243_n261# a_47_n42# a_n47_n139# a_n105_n42#
+ VSUBS
X0 a_47_n42# a_n47_n139# a_n105_n42# w_n243_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.47
C0 a_n47_n139# w_n243_n261# 0.27f
C1 a_47_n42# a_n105_n42# 0.0406f
C2 a_47_n42# w_n243_n261# 0.0499f
C3 a_47_n42# a_n47_n139# 0.00866f
C4 w_n243_n261# a_n105_n42# 0.0499f
C5 a_n47_n139# a_n105_n42# 0.00866f
C6 a_47_n42# VSUBS 0.0297f
C7 a_n105_n42# VSUBS 0.0297f
C8 a_n47_n139# VSUBS 0.168f
C9 w_n243_n261# VSUBS 1.17f
.ends

.subckt sky130_fd_pr__pfet_01v8_3PDS9J a_n102_n42# a_44_n42# a_n44_n139# w_n240_n261#
+ VSUBS
X0 a_44_n42# a_n44_n139# a_n102_n42# w_n240_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.44
C0 a_n44_n139# w_n240_n261# 0.261f
C1 a_44_n42# a_n102_n42# 0.0423f
C2 a_44_n42# w_n240_n261# 0.0499f
C3 a_44_n42# a_n44_n139# 0.00823f
C4 w_n240_n261# a_n102_n42# 0.0499f
C5 a_n44_n139# a_n102_n42# 0.00823f
C6 a_44_n42# VSUBS 0.0296f
C7 a_n102_n42# VSUBS 0.0296f
C8 a_n44_n139# VSUBS 0.16f
C9 w_n240_n261# VSUBS 1.15f
.ends

.subckt sky130_fd_pr__nfet_01v8_97T34Z a_n73_n46# a_n175_n220# a_n33_n134# a_15_n46#
X0 a_15_n46# a_n33_n134# a_n73_n46# a_n175_n220# sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.5 as=0.133 ps=1.5 w=0.46 l=0.15
C0 a_n73_n46# a_n33_n134# 0.0212f
C1 a_n33_n134# a_15_n46# 0.0212f
C2 a_n73_n46# a_15_n46# 0.0763f
C3 a_15_n46# a_n175_n220# 0.0769f
C4 a_n73_n46# a_n175_n220# 0.0769f
C5 a_n33_n134# a_n175_n220# 0.338f
.ends

.subckt th06 Vp Vin V06 Vn
XXM0 Vin m1_528_n874# Vn Vn sky130_fd_pr__nfet_01v8_L7T3GD
XXM1 Vp m1_528_n874# Vin Vp Vn sky130_fd_pr__pfet_01v8_NZD9V2
XXM2 Vp V06 m1_528_n874# Vp Vn sky130_fd_pr__pfet_01v8_3PDS9J
XXM3 Vn Vn m1_528_n874# V06 sky130_fd_pr__nfet_01v8_97T34Z
C0 m1_528_n874# V06 0.135f
C1 m1_528_n874# Vp 0.467f
C2 Vin V06 2.39e-21
C3 Vin Vp 0.192f
C4 m1_528_n874# Vin 0.224f
C5 V06 Vp 0.109f
C6 Vin Vn 0.726f
C7 V06 Vn 0.353f
C8 m1_528_n874# Vn 0.971f
C9 Vp Vn 2.62f
.ends


.GLOBAL VDD
.GLOBAL GND
.GLOBAL V_LH
.GLOBAL V_LL
.end
