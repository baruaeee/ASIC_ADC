magic
tech sky130A
magscale 1 2
timestamp 1704739411
<< pwell >>
rect -201 -2298 201 2298
<< psubdiff >>
rect -165 2228 -69 2262
rect 69 2228 165 2262
rect -165 2166 -131 2228
rect 131 2166 165 2228
rect -165 -2228 -131 -2166
rect 131 -2228 165 -2166
rect -165 -2262 -69 -2228
rect 69 -2262 165 -2228
<< psubdiffcont >>
rect -69 2228 69 2262
rect -165 -2166 -131 2166
rect 131 -2166 165 2166
rect -69 -2262 69 -2228
<< xpolycontact >>
rect -35 1700 35 2132
rect -35 -2132 35 -1700
<< xpolyres >>
rect -35 -1700 35 1700
<< locali >>
rect -165 2228 -69 2262
rect 69 2228 165 2262
rect -165 2166 -131 2228
rect 131 2166 165 2228
rect -165 -2228 -131 -2166
rect 131 -2228 165 -2166
rect -165 -2262 -69 -2228
rect 69 -2262 165 -2228
<< viali >>
rect -19 1717 19 2114
rect -19 -2114 19 -1717
<< metal1 >>
rect -25 2114 25 2126
rect -25 1717 -19 2114
rect 19 1717 25 2114
rect -25 1705 25 1717
rect -25 -1717 25 -1705
rect -25 -2114 -19 -1717
rect 19 -2114 25 -1717
rect -25 -2126 25 -2114
<< properties >>
string FIXED_BBOX -148 -2245 148 2245
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 17.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 98.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
