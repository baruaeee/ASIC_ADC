magic
tech sky130A
magscale 1 2
timestamp 1705501067
<< metal1 >>
rect 29058 10082 33964 10084
rect 29058 10015 33966 10082
rect 32218 9840 32287 10015
rect 33766 9772 33966 10015
rect 26274 9590 26280 9648
rect 26349 9590 26355 9648
rect 33303 9494 33309 9557
rect 33378 9494 33461 9557
rect 31856 9110 31862 9179
rect 31931 9110 32036 9179
rect 34966 9126 35149 9127
rect 34966 9062 35084 9126
rect 35148 9062 35154 9126
rect 33168 8728 33206 8770
rect 33200 8707 33206 8728
rect 33270 8707 33276 8770
rect 31483 8552 31760 8610
rect 28983 8464 29041 8470
rect 28983 8400 29041 8406
rect 31624 8319 31693 8422
rect 31624 8250 31629 8319
rect 31687 8250 31693 8319
rect 33399 8257 33513 8277
rect 31629 8243 31687 8249
rect 32139 8216 32193 8257
rect 33307 8216 33513 8257
rect 32139 8162 33513 8216
rect 32141 7847 32195 8162
rect 27671 7793 33851 7847
rect 27671 7719 27725 7793
rect 27401 7665 27725 7719
rect 28475 7513 28529 7793
rect 28869 7445 28923 7793
rect 28869 7387 28939 7445
rect 28885 7190 28939 7387
rect 30039 7361 30093 7793
rect 31284 7355 31342 7793
rect 33797 7685 33851 7793
rect 35686 7438 35692 7498
rect 35761 7438 35767 7498
rect 35696 7352 35756 7438
rect 35634 7292 35756 7352
rect 31860 7248 31932 7254
rect 28872 7136 28878 7190
rect 28947 7136 28953 7190
rect 31856 7188 31862 7248
rect 31931 7188 31937 7248
rect 29077 6992 29139 6994
rect 29068 6934 29074 6992
rect 29143 6934 29149 6992
rect 31860 6984 31932 7188
rect 27630 6906 27691 6911
rect 27620 6854 27626 6906
rect 27695 6854 27701 6906
rect 27630 6736 27691 6854
rect 29077 6743 29139 6934
rect 30476 6871 30534 6877
rect 30476 6796 30534 6802
rect 28845 6082 28912 6209
rect 30144 6194 30204 6402
rect 31636 6314 31918 6348
rect 31636 6288 31858 6314
rect 31852 6254 31858 6288
rect 31918 6254 31924 6314
rect 31982 6224 32046 6260
rect 30134 6134 30140 6194
rect 30209 6134 30215 6194
rect 31982 6184 32056 6224
rect 30986 6098 31042 6164
rect 31974 6124 31980 6184
rect 32049 6124 32056 6184
rect 31982 6122 32056 6124
rect 28838 6030 28844 6082
rect 28913 6030 28919 6082
rect 28845 6023 28912 6030
rect 31838 5848 33208 5908
rect 33584 5848 34984 5908
rect 31838 5736 31898 5848
rect 30894 5676 31898 5736
rect 30522 5642 30582 5648
rect 30894 5642 30954 5676
rect 27874 5607 27934 5613
rect 28178 5602 30522 5642
rect 27934 5582 30522 5602
rect 30582 5582 30954 5642
rect 27934 5542 28238 5582
rect 27874 5532 27934 5538
rect 28178 4946 28238 5542
rect 29824 4966 29884 5582
rect 30522 5576 30582 5582
rect 30894 5268 30954 5582
rect 30894 5208 31572 5268
rect 31512 4820 31572 5208
rect 34924 5048 34984 5848
rect 29214 4562 29220 4622
rect 29289 4562 29295 4622
rect 30672 4577 30846 4658
rect 29224 4484 29284 4562
rect 30672 4538 30753 4577
rect 27402 4082 27481 4289
rect 28958 4284 29526 4484
rect 30664 4478 30670 4538
rect 30755 4478 30761 4538
rect 30672 4468 30753 4478
rect 30366 4401 30434 4458
rect 30366 4400 30534 4401
rect 30366 4322 30616 4400
rect 30426 4320 30616 4322
rect 30548 4264 30616 4320
rect 30542 4212 30548 4264
rect 30617 4212 30623 4264
rect 30548 4204 30616 4212
rect 31989 4131 32049 4137
rect 27393 3998 27399 4082
rect 27483 3998 27489 4082
rect 31987 4064 31989 4129
rect 32049 4064 32270 4129
rect 31989 4056 32049 4062
rect 28108 3838 29210 3922
rect 28108 3604 28192 3838
rect 29126 3740 29210 3838
rect 31738 3830 31790 3836
rect 29861 3740 29919 3803
rect 29126 3703 29919 3740
rect 30819 3703 30877 3795
rect 31631 3748 31738 3827
rect 31790 3748 31804 3827
rect 31738 3739 31790 3745
rect 29126 3656 30877 3703
rect 28855 3199 28939 3205
rect 28672 3115 28855 3199
rect 28939 3115 28942 3199
rect 28855 3109 28942 3115
rect 27539 2484 27600 2784
rect 28858 2728 28942 3109
rect 29474 2812 29558 3656
rect 29861 3645 30877 3656
rect 30857 3291 31035 3349
rect 30857 2877 30915 3291
rect 31260 3224 31317 3324
rect 34837 3272 34895 3471
rect 31260 3167 31825 3224
rect 34830 3220 34836 3272
rect 34896 3220 34902 3272
rect 34837 3217 34895 3220
rect 31768 2907 31825 3167
rect 32008 3074 32065 3076
rect 32002 3020 32008 3074
rect 32064 3020 32070 3074
rect 32008 2907 32065 3020
rect 31768 2850 32272 2907
rect 32008 2633 32065 2850
rect 31594 2627 31638 2628
rect 31594 2624 31683 2627
rect 31542 2621 31692 2624
rect 27521 2400 27527 2484
rect 27611 2400 27617 2484
rect 28278 1345 28330 1351
rect 28274 1280 28278 1340
rect 28486 1340 28546 2560
rect 31542 2552 31626 2621
rect 31683 2552 31692 2621
rect 32008 2576 33168 2633
rect 31542 2548 31692 2552
rect 31594 2546 31683 2548
rect 32135 2527 32192 2533
rect 32128 2458 32135 2527
rect 32192 2458 32198 2527
rect 32128 2329 32198 2458
rect 33111 2361 33168 2576
rect 33111 2327 34181 2361
rect 30193 2276 30279 2277
rect 30193 2220 30298 2276
rect 30063 2134 30298 2220
rect 33111 2200 33177 2327
rect 33143 2199 33177 2200
rect 30063 2132 30279 2134
rect 29758 2072 29998 2079
rect 29758 2018 29930 2072
rect 29999 2018 30005 2072
rect 30057 2056 30063 2132
rect 30139 2121 30279 2132
rect 30139 2056 30145 2121
rect 35524 2051 35578 2057
rect 29758 2011 29998 2018
rect 35383 1983 35524 2050
rect 35578 1983 35585 2050
rect 35524 1976 35578 1982
rect 32615 1783 33539 1913
rect 29018 1340 29078 1548
rect 30760 1434 30934 1494
rect 30760 1384 30868 1434
rect 30748 1381 30868 1384
rect 31664 1381 34904 1436
rect 30748 1376 34904 1381
rect 30748 1373 33755 1376
rect 30748 1340 31724 1373
rect 28330 1320 31724 1340
rect 28330 1280 30868 1320
rect 28278 1270 28330 1276
<< via1 >>
rect 26280 9590 26349 9648
rect 33309 9494 33378 9557
rect 31862 9110 31931 9179
rect 35084 9062 35148 9126
rect 33206 8707 33270 8770
rect 28983 8406 29041 8464
rect 31629 8249 31687 8319
rect 35692 7438 35761 7498
rect 28878 7136 28947 7190
rect 31862 7188 31931 7248
rect 29074 6934 29143 6992
rect 27626 6854 27695 6906
rect 30476 6802 30534 6871
rect 31858 6254 31918 6314
rect 30140 6134 30209 6194
rect 31980 6124 32049 6184
rect 28844 6030 28913 6082
rect 27874 5538 27934 5607
rect 30522 5582 30582 5642
rect 29220 4562 29289 4622
rect 30670 4478 30755 4538
rect 30548 4212 30617 4264
rect 27399 3998 27483 4082
rect 31989 4062 32049 4131
rect 31738 3745 31790 3830
rect 28855 3115 28939 3199
rect 34836 3220 34896 3272
rect 32008 3020 32064 3074
rect 27527 2400 27611 2484
rect 28278 1276 28330 1345
rect 31626 2552 31683 2621
rect 32135 2458 32192 2527
rect 29930 2018 29999 2072
rect 30063 2056 30139 2132
rect 35524 1982 35578 2051
<< metal2 >>
rect 26280 10243 29383 10312
rect 26280 9648 26349 10243
rect 29314 10219 29383 10243
rect 29314 10150 33966 10219
rect 26280 9584 26349 9590
rect 31862 9179 31931 10150
rect 33309 9557 33378 10150
rect 33309 9488 33378 9494
rect 35084 9166 35148 9170
rect 35079 9126 35088 9166
rect 35144 9126 35153 9166
rect 35079 9110 35084 9126
rect 35148 9110 35153 9126
rect 28977 8406 28983 8464
rect 29041 8463 29400 8464
rect 29041 8407 29343 8463
rect 29399 8407 29408 8463
rect 29041 8406 29400 8407
rect 31677 8319 31736 8323
rect 31623 8249 31629 8319
rect 31687 8314 31741 8319
rect 31736 8255 31741 8314
rect 31687 8249 31741 8255
rect 31677 8246 31736 8249
rect 31862 7725 31931 9110
rect 35084 9056 35148 9062
rect 33206 8770 33270 8776
rect 33201 8707 33206 8722
rect 33270 8707 33275 8722
rect 33201 8666 33210 8707
rect 33266 8666 33275 8707
rect 33206 8662 33270 8666
rect 27846 7656 31931 7725
rect 27846 7569 27915 7656
rect 27626 7500 27915 7569
rect 27626 6906 27695 7500
rect 28878 7190 28947 7196
rect 28874 7136 28878 7142
rect 28947 7136 28951 7142
rect 28874 7083 28883 7136
rect 28942 7083 28951 7136
rect 28878 7078 28947 7083
rect 29074 6992 29143 7656
rect 29074 6928 29143 6934
rect 27626 6848 27695 6854
rect 30378 6871 30447 7656
rect 31862 7248 31931 7656
rect 35692 7544 35761 7549
rect 35688 7498 35697 7544
rect 35756 7498 35765 7544
rect 35688 7485 35692 7498
rect 35761 7485 35765 7498
rect 35692 7432 35761 7438
rect 31862 7182 31931 7188
rect 30378 6802 30476 6871
rect 30534 6802 30540 6871
rect 31858 6314 31918 6320
rect 31851 6254 31858 6268
rect 31918 6254 31925 6268
rect 31851 6212 31860 6254
rect 31916 6212 31925 6254
rect 31858 6210 31918 6212
rect 30140 6194 30209 6200
rect 30140 6122 30209 6134
rect 31980 6184 32049 6190
rect 28844 6082 28913 6088
rect 30136 6063 30145 6122
rect 30204 6063 30213 6122
rect 30140 6058 30209 6063
rect 28844 6020 28913 6030
rect 28840 5961 28849 6020
rect 28908 5961 28917 6020
rect 28844 5956 28913 5961
rect 30582 5642 30638 5649
rect 27811 5607 27870 5611
rect 27806 5602 27874 5607
rect 27806 5542 27811 5602
rect 27870 5542 27874 5602
rect 27806 5538 27874 5542
rect 27934 5538 27940 5607
rect 30516 5582 30522 5642
rect 30582 5640 30640 5642
rect 30638 5584 30640 5640
rect 30582 5582 30640 5584
rect 30582 5575 30638 5582
rect 27811 5533 27870 5538
rect 31980 5334 32049 6124
rect 29220 5265 32049 5334
rect 29220 4622 29289 5265
rect 27399 4082 27483 4088
rect 27399 3992 27411 3998
rect 27402 3955 27411 3992
rect 27470 3992 27483 3998
rect 27470 3955 27479 3992
rect 27406 3950 27475 3955
rect 29220 3571 29289 4562
rect 30670 4538 30755 4544
rect 30670 4462 30755 4478
rect 30666 4387 30675 4462
rect 30750 4387 30759 4462
rect 30670 4382 30755 4387
rect 30548 4264 30617 4270
rect 30548 4186 30617 4212
rect 30544 4127 30553 4186
rect 30612 4127 30621 4186
rect 31980 4131 32049 5265
rect 30548 4122 30617 4127
rect 31980 4062 31989 4131
rect 32049 4062 32055 4131
rect 31980 3830 32049 4062
rect 31732 3745 31738 3830
rect 31790 3758 32049 3830
rect 31790 3745 32048 3758
rect 28862 3502 29289 3571
rect 28862 3199 28931 3502
rect 28849 3115 28855 3199
rect 28939 3115 28945 3199
rect 31882 2621 31951 3745
rect 34836 3272 34896 3278
rect 34829 3220 34836 3222
rect 34896 3220 34903 3222
rect 34829 3166 34838 3220
rect 34894 3166 34903 3220
rect 34836 3164 34896 3166
rect 31999 3062 32008 3118
rect 32064 3062 32073 3118
rect 32008 3014 32064 3020
rect 31620 2552 31626 2621
rect 31683 2552 31951 2621
rect 31882 2527 31951 2552
rect 27527 2484 27611 2490
rect 31882 2458 32135 2527
rect 32192 2458 32198 2527
rect 27527 2394 27539 2400
rect 27530 2365 27539 2394
rect 27598 2394 27611 2400
rect 27598 2365 27607 2394
rect 27534 2360 27603 2365
rect 30063 2132 30139 2138
rect 29930 2072 29999 2078
rect 30062 2056 30063 2076
rect 29926 1959 29935 2018
rect 29994 1959 30003 2018
rect 30062 2017 30071 2056
rect 30130 2017 30139 2056
rect 35581 2051 35640 2055
rect 30066 2012 30135 2017
rect 35518 1982 35524 2051
rect 35578 2046 35645 2051
rect 35578 1987 35581 2046
rect 35640 1987 35645 2046
rect 35578 1982 35645 1987
rect 35581 1978 35640 1982
rect 29930 1954 29999 1959
rect 28198 1345 28257 1349
rect 28193 1340 28278 1345
rect 28193 1281 28198 1340
rect 28257 1281 28278 1340
rect 28193 1276 28278 1281
rect 28330 1276 28336 1345
rect 28198 1272 28257 1276
<< via2 >>
rect 35088 9126 35144 9166
rect 35088 9110 35144 9126
rect 29343 8407 29399 8463
rect 31677 8255 31687 8314
rect 31687 8255 31736 8314
rect 33210 8707 33266 8722
rect 33210 8666 33266 8707
rect 28883 7136 28942 7142
rect 28883 7083 28942 7136
rect 35697 7498 35756 7544
rect 35697 7485 35756 7498
rect 31860 6254 31916 6268
rect 31860 6212 31916 6254
rect 30145 6063 30204 6122
rect 28849 5961 28908 6020
rect 27811 5542 27870 5602
rect 30582 5584 30638 5640
rect 27411 3998 27470 4014
rect 27411 3955 27470 3998
rect 30675 4387 30750 4462
rect 30553 4127 30612 4186
rect 34838 3220 34894 3222
rect 34838 3166 34894 3220
rect 32008 3074 32064 3118
rect 32008 3062 32064 3074
rect 27539 2400 27598 2424
rect 27539 2365 27598 2400
rect 30071 2056 30130 2076
rect 29935 1959 29994 2018
rect 30071 2017 30130 2056
rect 35581 1987 35640 2046
rect 28198 1281 28257 1340
<< metal3 >>
rect 35086 10082 35302 10142
rect 35086 9171 35146 10082
rect 35083 9166 35149 9171
rect 35083 9110 35088 9166
rect 35144 9110 35149 9166
rect 35083 9105 35149 9110
rect 33205 8722 33271 8727
rect 33205 8666 33210 8722
rect 33266 8666 33271 8722
rect 33205 8661 33271 8666
rect 29340 8470 29400 8476
rect 29332 8466 29338 8470
rect 29330 8464 29338 8466
rect 29266 8406 29338 8464
rect 29402 8464 29408 8470
rect 29402 8406 29410 8464
rect 29266 8404 29410 8406
rect 29270 8402 29404 8404
rect 31672 8314 31741 8319
rect 31672 8255 31677 8314
rect 31736 8255 31864 8314
rect 31672 8254 31864 8255
rect 31672 8250 31741 8254
rect 31804 7988 31864 8254
rect 33208 8124 33268 8661
rect 35370 8124 35430 9748
rect 33208 8064 35430 8124
rect 35536 7988 35596 9396
rect 31804 7928 35596 7988
rect 35696 7549 35756 9322
rect 35692 7544 35761 7549
rect 35692 7485 35697 7544
rect 35756 7485 35761 7544
rect 35692 7480 35761 7485
rect 28878 7143 28947 7147
rect 28877 7142 28948 7143
rect 28877 7083 28883 7142
rect 28942 7083 28948 7142
rect 28877 7058 28948 7083
rect 28874 6994 28880 7058
rect 28944 6994 28950 7058
rect 35918 6968 35978 8898
rect 35622 6908 35978 6968
rect 31855 6268 31921 6273
rect 31855 6212 31860 6268
rect 31916 6212 31921 6268
rect 31855 6207 31921 6212
rect 30140 6122 30209 6127
rect 30140 6063 30145 6122
rect 30204 6063 30209 6122
rect 30140 6058 30209 6063
rect 31858 6084 31918 6207
rect 28844 6020 28913 6025
rect 28844 5961 28849 6020
rect 28908 5961 28913 6020
rect 28844 5956 28913 5961
rect 27732 5607 27796 5610
rect 27729 5604 27875 5607
rect 27729 5540 27732 5604
rect 27796 5602 27875 5604
rect 27796 5542 27811 5602
rect 27870 5542 27875 5602
rect 27796 5540 27875 5542
rect 27729 5537 27875 5540
rect 27732 5534 27796 5537
rect 28848 5466 28908 5956
rect 30144 5498 30204 6058
rect 31858 6024 32106 6084
rect 31858 6020 31918 6024
rect 32046 5718 32106 6024
rect 35622 5718 35682 6908
rect 32046 5658 35682 5718
rect 35810 6702 36322 6762
rect 30422 5644 30486 5650
rect 30577 5642 30643 5645
rect 30486 5640 30643 5642
rect 30486 5584 30582 5640
rect 30638 5584 30643 5640
rect 30486 5582 30643 5584
rect 30422 5574 30486 5580
rect 30577 5579 30643 5582
rect 35810 5580 35870 6702
rect 31050 5520 35870 5580
rect 35982 6458 36310 6518
rect 31050 5498 31110 5520
rect 28848 5406 29982 5466
rect 30144 5438 31110 5498
rect 35982 5420 36042 6458
rect 29922 5348 29982 5406
rect 31264 5360 36042 5420
rect 31264 5348 31324 5360
rect 29922 5288 31324 5348
rect 30670 4462 30755 4467
rect 30670 4387 30675 4462
rect 30750 4387 30755 4462
rect 30670 4382 30755 4387
rect 30548 4186 30617 4191
rect 30548 4127 30553 4186
rect 30612 4127 30617 4186
rect 30548 4122 30617 4127
rect 27406 4014 27475 4019
rect 27406 3955 27411 4014
rect 27470 3955 27475 4014
rect 27406 3950 27475 3955
rect 27410 3800 27470 3950
rect 30552 3910 30612 4122
rect 30682 3210 30742 4382
rect 34836 3227 34896 3228
rect 34833 3222 34899 3227
rect 30682 3150 31116 3210
rect 31056 3104 31116 3150
rect 31998 3148 32004 3212
rect 32068 3148 32074 3212
rect 34833 3166 34838 3222
rect 34894 3166 34899 3222
rect 34833 3161 34899 3166
rect 32000 3118 32069 3148
rect 31056 3044 31696 3104
rect 32000 3099 32008 3118
rect 32003 3062 32008 3099
rect 32064 3062 32069 3118
rect 32003 3057 32069 3062
rect 31636 2776 31696 3044
rect 31636 2716 31798 2776
rect 27538 2429 27598 2433
rect 27534 2424 27603 2429
rect 27534 2365 27539 2424
rect 27598 2365 27603 2424
rect 27534 2360 27603 2365
rect 31738 2380 31798 2716
rect 34836 2576 34896 3161
rect 34836 2516 36154 2576
rect 27538 2278 27598 2360
rect 31738 2320 32028 2380
rect 30066 2076 30135 2081
rect 29930 2018 29999 2023
rect 29930 1959 29935 2018
rect 29994 1959 29999 2018
rect 30066 2017 30071 2076
rect 30130 2017 30135 2076
rect 30066 2012 30135 2017
rect 29930 1954 29999 1959
rect 29934 1790 29994 1954
rect 30070 1788 30130 2012
rect 28104 1345 28168 1348
rect 28102 1342 28262 1345
rect 28102 1278 28104 1342
rect 28168 1340 28262 1342
rect 28168 1281 28198 1340
rect 28257 1281 28262 1340
rect 28168 1278 28262 1281
rect 28102 1276 28262 1278
rect 31968 1334 32028 2320
rect 35576 2046 35645 2051
rect 35748 2046 36192 2047
rect 35576 1987 35581 2046
rect 35640 1987 36192 2046
rect 35576 1986 36192 1987
rect 35576 1982 35645 1986
rect 28104 1272 28168 1276
rect 31968 1274 36228 1334
<< via3 >>
rect 29338 8463 29402 8470
rect 29338 8407 29343 8463
rect 29343 8407 29399 8463
rect 29399 8407 29402 8463
rect 29338 8406 29402 8407
rect 28880 6994 28944 7058
rect 27732 5540 27796 5604
rect 30422 5580 30486 5644
rect 32004 3148 32068 3212
rect 28104 1278 28168 1342
<< metal4 >>
rect 29337 8470 29403 8471
rect 29337 8406 29338 8470
rect 29402 8406 29403 8470
rect 29337 8405 29403 8406
rect 29340 7608 29400 8405
rect 29340 7548 30330 7608
rect 28879 7058 28945 7059
rect 28879 6994 28880 7058
rect 28944 6994 28945 7058
rect 28879 6993 28945 6994
rect 28882 6530 28942 6993
rect 28882 6470 29122 6530
rect 27731 5604 27797 5605
rect 27731 5602 27732 5604
rect 27300 5542 27732 5602
rect 27300 1340 27360 5542
rect 27731 5540 27732 5542
rect 27796 5540 27797 5604
rect 27731 5539 27797 5540
rect 29062 5564 29122 6470
rect 30270 5642 30330 7548
rect 30421 5644 30487 5645
rect 30421 5642 30422 5644
rect 30270 5582 30422 5642
rect 30421 5580 30422 5582
rect 30486 5580 30487 5644
rect 30421 5579 30487 5580
rect 29062 5504 29400 5564
rect 29340 5190 29400 5504
rect 29340 5130 31876 5190
rect 31816 3934 31876 5130
rect 31816 3874 32066 3934
rect 32006 3213 32066 3874
rect 32003 3212 32069 3213
rect 32003 3148 32004 3212
rect 32068 3148 32069 3212
rect 32003 3147 32069 3148
rect 28103 1342 28169 1343
rect 28103 1340 28104 1342
rect 27300 1280 28104 1340
rect 28103 1278 28104 1280
rect 28168 1278 28169 1342
rect 28103 1277 28169 1278
use th09  th09_0
timestamp 1705440721
transform 1 0 31258 0 1 9576
box 670 -1498 1918 398
use th02  x16
timestamp 1705440580
transform 1 0 31040 0 1 4594
box 1100 -1960 4395 680
use th03  x17
timestamp 1705440596
transform -1 0 32014 0 -1 2072
box 414 -920 1840 706
use th04  x18
timestamp 1705440610
transform -1 0 32004 0 1 4580
box 279 -1300 1216 476
use th05  x19
timestamp 1705440623
transform -1 0 29462 0 1 4794
box 394 -966 2064 258
use th06  x20
timestamp 1705440654
transform -1 0 29068 0 -1 2576
box 308 -1110 1542 62
use th07  x21
timestamp 1705440679
transform 1 0 29030 0 1 5058
box 296 -1290 1462 -44
use th08  x22
timestamp 1705440694
transform 1 0 28494 0 -1 1540
box 330 -1392 1396 54
use th10  x24
timestamp 1705440736
transform 1 0 28612 0 -1 6332
box 394 -1164 1590 790
use th11  x25
timestamp 1705440755
transform 1 0 27384 0 -1 6988
box 160 -636 1584 1464
use th12  x26
timestamp 1705481551
transform 1 0 30095 0 -1 6400
box 375 -1092 1662 716
use th13  x27
timestamp 1705440792
transform 1 0 33074 0 1 9416
box 240 -1200 2062 556
use th14  x28
timestamp 1705440829
transform 1 0 31552 0 -1 6548
box 300 -1200 4172 772
use th15  x29
timestamp 1705440844
transform 1 0 25327 0 1 8330
box 915 -950 6436 1862
use preamp  x30
timestamp 1705440528
transform 1 0 31712 0 -1 2152
box 398 -255 1470 780
use th01  x31
timestamp 1705440556
transform 1 0 32796 0 -1 1194
box 618 -1168 2664 -180
<< end >>
