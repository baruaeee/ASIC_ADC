magic
tech sky130A
magscale 1 2
timestamp 1706473616
<< error_p >>
rect -29 131 29 137
rect -29 97 -17 131
rect -29 91 29 97
rect -29 -97 29 -91
rect -29 -131 -17 -97
rect -29 -137 29 -131
<< nwell >>
rect -219 -269 219 269
<< pmos >>
rect -23 -50 23 50
<< pdiff >>
rect -81 38 -23 50
rect -81 -38 -69 38
rect -35 -38 -23 38
rect -81 -50 -23 -38
rect 23 38 81 50
rect 23 -38 35 38
rect 69 -38 81 38
rect 23 -50 81 -38
<< pdiffc >>
rect -69 -38 -35 38
rect 35 -38 69 38
<< nsubdiff >>
rect -183 -27 -149 35
rect -183 -199 -149 -137
<< nsubdiffcont >>
rect -183 -137 -149 -27
<< poly >>
rect -33 131 33 147
rect -33 97 -17 131
rect 17 97 33 131
rect -33 81 33 97
rect -23 50 23 81
rect -23 -81 23 -50
rect -33 -97 33 -81
rect -33 -131 -17 -97
rect 17 -131 33 -97
rect -33 -147 33 -131
<< polycont >>
rect -17 97 17 131
rect -17 -131 17 -97
<< locali >>
rect -33 97 -17 131
rect 17 97 33 131
rect -69 38 -35 54
rect -183 -27 -149 35
rect -69 -54 -35 -38
rect 35 38 69 54
rect 35 -54 69 -38
rect -33 -131 -17 -97
rect 17 -131 33 -97
rect -183 -199 -149 -137
<< viali >>
rect -17 97 17 131
rect -69 -38 -35 38
rect 35 -38 69 38
rect -17 -131 17 -97
<< metal1 >>
rect -29 131 29 137
rect -29 97 -17 131
rect 17 97 29 131
rect -29 91 29 97
rect -75 38 -29 50
rect -75 -38 -69 38
rect -35 -38 -29 38
rect -75 -50 -29 -38
rect 29 38 75 50
rect 29 -38 35 38
rect 69 -38 75 38
rect 29 -50 75 -38
rect -29 -97 29 -91
rect -29 -131 -17 -97
rect 17 -131 29 -97
rect -29 -137 29 -131
<< properties >>
string FIXED_BBOX -166 -216 166 216
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 0.227 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
