magic
tech sky130A
magscale 1 2
timestamp 1702941823
<< checkpaint >>
rect 735 -925 3963 2099
<< error_s >>
rect 1626 1139 1679 1142
rect 1608 1106 1679 1139
rect 1626 1072 1697 1106
rect 1439 1037 1497 1043
rect 584 999 619 1033
rect 1293 1016 1327 1034
rect 585 980 619 999
rect 604 583 619 980
rect 638 946 673 980
rect 638 583 672 946
rect 638 549 653 583
rect 1257 530 1327 1016
rect 1439 1003 1451 1037
rect 1439 997 1497 1003
rect 1439 613 1497 619
rect 1439 579 1451 613
rect 1439 573 1497 579
rect 1257 494 1310 530
rect 1626 477 1696 1072
rect 1808 1004 1866 1010
rect 1808 970 1820 1004
rect 1808 964 1866 970
rect 1808 560 1866 566
rect 1808 526 1820 560
rect 1808 520 1866 526
rect 1626 441 1679 477
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_XYZSMQ  XM1
timestamp 0
transform 1 0 1837 0 1 765
box -211 -377 211 377
use sky130_fd_pr__nfet_01v8_2V6S9N  XM3
timestamp 0
transform 1 0 2349 0 1 587
box -354 -252 354 252
use sky130_fd_pr__pfet_01v8_AZD98U  XM7
timestamp 0
transform 1 0 301 0 1 808
box -354 -261 354 261
use sky130_fd_pr__pfet_01v8_AZD98U  XM9
timestamp 0
transform 1 0 956 0 1 755
box -354 -261 354 261
use sky130_fd_pr__nfet_01v8_T8HSQ7  XM10
timestamp 0
transform 1 0 1468 0 1 808
box -211 -367 211 367
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
