magic
tech sky130A
magscale 1 2
timestamp 1706197322
<< error_p >>
rect 422 215 456 246
<< pwell >>
rect -446 -252 446 252
<< nmos >>
rect -250 -42 250 42
<< ndiff >>
rect -308 30 -250 42
rect -308 -30 -296 30
rect -262 -30 -250 30
rect -308 -42 -250 -30
rect 250 30 308 42
rect 250 -30 262 30
rect 296 -30 308 30
rect 250 -42 308 -30
<< ndiffc >>
rect -296 -30 -262 30
rect 262 -30 296 30
<< psubdiff >>
rect -410 182 -259 216
rect 422 215 456 246
rect -410 120 -376 182
rect -410 -182 -376 -120
rect 376 -182 410 129
rect -410 -216 -314 -182
rect 314 -216 410 -182
<< psubdiffcont >>
rect -410 -120 -376 120
rect -314 -216 314 -182
<< poly >>
rect -250 114 250 130
rect -250 80 -234 114
rect 234 80 250 114
rect -250 42 250 80
rect -250 -80 250 -42
rect -250 -114 -234 -80
rect 234 -114 250 -80
rect -250 -130 250 -114
<< polycont >>
rect -234 80 234 114
rect -234 -114 234 -80
<< locali >>
rect -410 182 -265 216
rect -410 120 -376 182
rect 376 161 455 195
rect -250 80 -234 114
rect 234 80 250 114
rect -296 30 -262 46
rect -296 -46 -262 -30
rect 262 30 296 46
rect 262 -46 296 -30
rect -250 -114 -234 -80
rect 234 -114 250 -80
rect -410 -182 -376 -120
rect 376 -182 410 161
rect -410 -216 -314 -182
rect 314 -216 410 -182
<< viali >>
rect -234 80 234 114
rect -296 -30 -262 30
rect 262 -30 296 30
rect -234 -114 234 -80
<< metal1 >>
rect -246 114 246 120
rect -246 80 -234 114
rect 234 80 246 114
rect -246 74 246 80
rect -302 30 -256 42
rect -302 -30 -296 30
rect -262 -30 -256 30
rect -302 -42 -256 -30
rect 256 30 302 42
rect 256 -30 262 30
rect 296 -30 302 30
rect 256 -42 302 -30
rect -246 -80 246 -74
rect -246 -114 -234 -80
rect 234 -114 246 -80
rect -246 -120 246 -114
<< properties >>
string FIXED_BBOX -392 -198 392 198
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 2.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
