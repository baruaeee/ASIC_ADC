magic
tech sky130A
magscale 1 2
timestamp 1702941822
<< checkpaint >>
rect -84 -872 2858 2152
<< error_s >>
rect 356 1006 391 1024
rect 356 999 427 1006
rect 357 970 427 999
rect 374 936 445 970
rect 725 963 760 970
rect 725 936 796 963
rect 374 583 444 936
rect 726 927 796 936
rect 743 893 814 927
rect 556 868 614 874
rect 556 834 568 868
rect 556 828 614 834
rect 556 666 614 672
rect 556 632 568 666
rect 556 626 614 632
rect 374 547 427 583
rect 743 530 813 893
rect 743 494 796 530
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_NZD9V2  XM1
timestamp 0
transform 1 0 986 0 1 702
box -243 -261 243 261
use sky130_fd_pr__nfet_01v8_L7T3GD  XM3
timestamp 0
transform 1 0 1387 0 1 640
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_3PDS9J  XM7
timestamp 0
transform 1 0 187 0 1 808
box -240 -261 240 261
use sky130_fd_pr__nfet_01v8_97T34Z  XM10
timestamp 0
transform 1 0 585 0 1 750
box -211 -256 211 256
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
