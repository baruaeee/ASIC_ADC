** sch_path: /home/exotic/Desktop/ASIC_ADC/xschem/Vth_sch/Pre_layout/th14.sch
**.subckt th14 Vin Vout
*.ipin Vin
*.opin Vout
VDD VDD GND 1.8
Vin Vin GND pulse(0 0.2 0ns 1ns 1ns 5ns 10ns)
V_logic_high V_LH GND 1.25
V_logic_low V_LL GND 0.5
x1 VDD Vout Vin GND th14
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.save all





.dc Vin 0 1.8 0.01
*.tran 1n 30n
.control
run
set color0=white
set color1=black
plot Vin Vout V_LH V_LL
set xbrushwidth=3
.save all
.endc
.end


**** end user architecture code
**.ends

* NGSPICE file created from th14.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_XJ7SDL a_15_n450# w_n211_n669# a_n73_n450# a_n33_n547#
+ VSUBS
X0 a_15_n450# a_n33_n547# a_n73_n450# w_n211_n669# sky130_fd_pr__pfet_01v8 ad=1.3 pd=9.58 as=1.3 ps=9.58 w=4.5 l=0.15
C0 a_n73_n450# w_n211_n669# 0.295f
C1 a_15_n450# a_n33_n547# 0.0407f
C2 w_n211_n669# a_n33_n547# 0.242f
C3 a_n73_n450# a_n33_n547# 0.0407f
C4 a_15_n450# w_n211_n669# 0.295f
C5 a_n73_n450# a_15_n450# 0.718f
C6 a_15_n450# VSUBS 0.191f
C7 a_n73_n450# VSUBS 0.191f
C8 a_n33_n547# VSUBS 0.122f
C9 w_n211_n669# VSUBS 2.46f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFMUVB a_n608_n42# a_550_n42# a_n710_n216# a_n550_n130#
X0 a_550_n42# a_n550_n130# a_n608_n42# a_n710_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=5.5
C0 a_550_n42# a_n550_n130# 0.0242f
C1 a_n550_n130# a_n608_n42# 0.0242f
C2 a_550_n42# a_n608_n42# 0.00526f
C3 a_550_n42# a_n710_n216# 0.0873f
C4 a_n608_n42# a_n710_n216# 0.0873f
C5 a_n550_n130# a_n710_n216# 3.19f
.ends

.subckt sky130_fd_pr__pfet_01v8_UJPVTG w_n211_n769# a_n73_n550# a_n33_n647# a_15_n550#
+ VSUBS
X0 a_15_n550# a_n33_n647# a_n73_n550# w_n211_n769# sky130_fd_pr__pfet_01v8 ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.15
C0 a_n73_n550# w_n211_n769# 0.356f
C1 a_15_n550# a_n33_n647# 0.0449f
C2 w_n211_n769# a_n33_n647# 0.242f
C3 a_n73_n550# a_n33_n647# 0.0449f
C4 a_15_n550# w_n211_n769# 0.356f
C5 a_n73_n550# a_15_n550# 0.877f
C6 a_15_n550# VSUBS 0.232f
C7 a_n73_n550# VSUBS 0.232f
C8 a_n33_n647# VSUBS 0.122f
C9 w_n211_n769# VSUBS 2.81f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GTR a_n608_n42# a_550_n42# w_n746_n261# a_n550_n139#
+ VSUBS
X0 a_550_n42# a_n550_n139# a_n608_n42# w_n746_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=5.5
C0 a_n608_n42# w_n746_n261# 0.0498f
C1 a_550_n42# a_n550_n139# 0.0242f
C2 w_n746_n261# a_n550_n139# 1.82f
C3 a_n608_n42# a_n550_n139# 0.0242f
C4 a_550_n42# w_n746_n261# 0.0498f
C5 a_n608_n42# a_550_n42# 0.00526f
C6 a_550_n42# VSUBS 0.037f
C7 a_n608_n42# VSUBS 0.037f
C8 a_n550_n139# VSUBS 1.44f
C9 w_n746_n261# VSUBS 3.22f
.ends

.subckt sky130_fd_pr__nfet_01v8_9GNSAM a_n73_n550# a_n175_n724# a_15_n550# a_n33_n638#
X0 a_15_n550# a_n33_n638# a_n73_n550# a_n175_n724# sky130_fd_pr__nfet_01v8 ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.15
C0 a_15_n550# a_n33_n638# 0.0468f
C1 a_n33_n638# a_n73_n550# 0.0468f
C2 a_15_n550# a_n73_n550# 0.877f
C3 a_15_n550# a_n175_n724# 0.588f
C4 a_n73_n550# a_n175_n724# 0.588f
C5 a_n33_n638# a_n175_n724# 0.352f
.ends

.subckt th14 Vp Vout Vin Vn
XXM0 m1_1594_n962# Vp Vn Vn Vn sky130_fd_pr__pfet_01v8_XJ7SDL
XXM1 m1_710_n388# m1_1594_n962# Vn Vin sky130_fd_pr__nfet_01v8_ZFMUVB
XXM2 Vp m1_710_n388# Vin Vp Vn sky130_fd_pr__pfet_01v8_UJPVTG
XXM3 Vp m1_2498_n384# Vp m1_710_n388# Vn sky130_fd_pr__pfet_01v8_VZ9GTR
XXM4 m1_2498_n384# Vout Vp m1_710_n388# Vn sky130_fd_pr__pfet_01v8_VZ9GTR
XXM5 Vn Vn Vout m1_710_n388# sky130_fd_pr__nfet_01v8_9GNSAM
C0 Vn m1_2498_n384# 3.16e-24
C1 Vn Vp 0.876f
C2 Vin m1_2498_n384# 1.46e-19
C3 Vin Vp 0.214f
C4 Vin Vn 0.0583f
C5 m1_1594_n962# Vp 0.237f
C6 m1_1594_n962# Vn 0.111f
C7 m1_710_n388# Vout 0.191f
C8 m1_1594_n962# Vin 0.166f
C9 m1_710_n388# m1_2498_n384# 0.768f
C10 m1_710_n388# Vp 0.755f
C11 m1_710_n388# Vn 0.459f
C12 m1_710_n388# Vin 0.365f
C13 m1_2498_n384# Vout 0.0142f
C14 Vp Vout 0.125f
C15 Vn Vout 0.0354f
C16 m1_1594_n962# m1_710_n388# 0.00647f
C17 Vp m1_2498_n384# 0.276f
C18 Vin 0 3.4f
C19 Vn 0 0.831f
C20 Vout 0 0.854f
C21 m1_2498_n384# 0 0.297f
C22 m1_710_n388# 0 3.52f
C23 Vp 0 11.9f
C24 m1_1594_n962# 0 0.292f
.ends


.GLOBAL VDD
.GLOBAL GND
.GLOBAL V_LH
.GLOBAL V_LL
.end
