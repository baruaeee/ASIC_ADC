magic
tech sky130A
magscale 1 2
timestamp 1704752409
<< locali >>
rect -20 854 126 1024
rect 1402 848 1552 1020
rect 2358 852 2508 1024
rect 2842 844 2988 1020
rect 352 184 722 360
rect 1406 184 1552 356
rect 2364 188 2510 360
rect 3010 188 3158 362
<< metal1 >>
rect 2338 1520 2538 1686
rect -55 1450 543 1520
rect 2338 1486 3977 1520
rect 2475 1453 3977 1486
rect -55 476 15 1450
rect 2491 1295 2525 1453
rect 61 1261 2875 1295
rect 61 1027 95 1261
rect 156 1151 324 1152
rect 156 1117 417 1151
rect 156 1085 323 1117
rect 383 1027 417 1117
rect 61 993 127 1027
rect 62 851 127 993
rect 351 851 417 1027
rect 62 850 96 851
rect 383 791 417 851
rect 635 1027 669 1261
rect 1473 1217 2427 1219
rect 1263 1185 2427 1217
rect 1263 1183 1849 1185
rect 635 849 705 1027
rect 924 1024 996 1028
rect 1263 1024 1297 1183
rect 924 990 1297 1024
rect 1473 1035 1507 1183
rect 924 890 996 990
rect 1268 905 1274 914
rect 929 851 996 890
rect 962 850 996 851
rect 1133 871 1274 905
rect 1133 791 1167 871
rect 1268 862 1274 871
rect 1326 862 1332 914
rect 1473 847 1553 1035
rect 1810 1023 1844 1024
rect 1775 989 1844 1023
rect 1775 881 1809 989
rect 1810 881 1844 989
rect 2070 881 2135 1025
rect 2393 1021 2427 1185
rect 1775 848 1844 881
rect 1775 847 1843 848
rect 155 757 1167 791
rect 383 583 417 757
rect 1289 717 1751 787
rect 383 549 1017 583
rect -55 409 921 476
rect -55 361 15 409
rect 983 361 1017 549
rect -55 181 131 361
rect 352 184 722 360
rect 501 29 568 184
rect 945 183 1017 361
rect 1163 234 1229 235
rect 1163 182 1170 234
rect 1222 182 1229 234
rect 1163 160 1229 182
rect 1054 29 1254 160
rect 501 -38 1254 29
rect 1054 -40 1254 -38
rect 1289 -107 1359 717
rect 1809 473 1843 847
rect 1581 407 1843 473
rect 1809 361 1843 407
rect 1490 359 1524 360
rect 1490 221 1553 359
rect 1489 187 1553 221
rect 1489 184 1524 187
rect 1489 -15 1523 184
rect 1777 183 1843 361
rect 2069 847 2135 881
rect 2359 847 2427 1021
rect 2839 877 2875 1261
rect 3226 1168 3278 1174
rect 3151 1146 3226 1155
rect 3017 1116 3226 1146
rect 3278 1146 3281 1155
rect 3278 1116 3283 1146
rect 3017 1112 3283 1116
rect 3017 1081 3185 1112
rect 3226 1110 3278 1112
rect 2921 877 2989 1023
rect 2069 569 2103 847
rect 2839 843 2989 877
rect 3213 879 3278 1023
rect 2165 757 2333 789
rect 2548 757 2748 814
rect 2163 723 2748 757
rect 2164 722 2332 723
rect 2548 614 2748 723
rect 2069 535 2557 569
rect 2839 565 2873 843
rect 3213 831 3309 879
rect 3275 782 3309 831
rect 3257 730 3263 782
rect 3315 730 3321 782
rect 3275 619 3309 730
rect 3275 615 3332 619
rect 3370 615 3570 788
rect 3275 588 3570 615
rect 3275 581 3447 588
rect 2069 363 2103 535
rect 2523 497 2557 535
rect 2740 531 2873 565
rect 2616 510 2668 516
rect 2523 463 2616 497
rect 2069 183 2141 363
rect 2365 253 2443 361
rect 2365 205 2399 253
rect 2403 205 2443 253
rect 2523 283 2557 463
rect 2616 452 2668 458
rect 2740 411 2774 531
rect 3060 461 3066 513
rect 3118 477 3124 513
rect 3188 477 3356 478
rect 3118 461 3356 477
rect 3067 444 3356 461
rect 3067 443 3355 444
rect 3187 413 3355 443
rect 3413 363 3447 581
rect 2649 283 2717 361
rect 2523 249 2717 283
rect 2365 171 2443 205
rect 2649 185 2717 249
rect 2801 251 2866 362
rect 3090 361 3124 362
rect 2801 185 2889 251
rect 3090 189 3159 361
rect 3381 215 3447 363
rect 3090 186 3125 189
rect 3381 187 3567 215
rect 2803 173 2889 185
rect 1581 103 1751 133
rect 2167 103 2337 137
rect 1581 69 2337 103
rect 1582 68 1751 69
rect 2409 -15 2443 171
rect 2724 88 2790 146
rect 2855 106 2889 173
rect 2841 54 2847 106
rect 2899 54 2905 106
rect 1489 -49 2443 -15
rect 109 -177 1359 -107
rect 2409 -143 2443 -49
rect 2658 -134 2710 -128
rect 2409 -177 2658 -143
rect 109 -237 545 -177
rect 2649 -186 2658 -177
rect 3091 -142 3125 186
rect 3405 185 3567 187
rect 3413 181 3567 185
rect 2946 -143 3378 -142
rect 2710 -186 3378 -143
rect 2649 -213 3378 -186
rect 2649 -233 2719 -213
rect 112 -450 544 -237
rect 1549 -303 2719 -233
rect 2945 -283 3378 -213
rect 3037 -285 3107 -283
rect 112 -706 546 -450
rect 3533 -637 3567 181
rect 3531 -645 3975 -637
rect 3531 -707 3977 -645
<< via1 >>
rect 1274 862 1326 914
rect 1170 182 1222 234
rect 3226 1116 3278 1168
rect 3263 730 3315 782
rect 2616 458 2668 510
rect 3066 461 3118 513
rect 2847 54 2899 106
rect 2658 -186 2710 -134
<< metal2 >>
rect 3220 1157 3226 1168
rect 2545 1155 3226 1157
rect 2544 1127 3226 1155
rect 2544 1125 2765 1127
rect 2544 1067 2575 1125
rect 3220 1116 3226 1127
rect 3278 1116 3284 1168
rect 1274 914 1326 920
rect 2544 903 2574 1067
rect 1326 873 2574 903
rect 1274 856 1326 862
rect 3263 782 3315 788
rect 3263 724 3315 730
rect 3066 513 3118 519
rect 2610 458 2616 510
rect 2668 505 2674 510
rect 2668 468 3066 505
rect 2668 466 2690 468
rect 2668 458 2674 466
rect 3066 455 3118 461
rect 1182 279 1309 309
rect 1182 264 1212 279
rect 1180 240 1212 264
rect 1170 234 1222 240
rect 1170 176 1222 182
rect 1279 -145 1309 279
rect 2847 106 2899 112
rect 2847 48 2899 54
rect 2652 -145 2658 -134
rect 1279 -175 2658 -145
rect 2533 -854 2563 -175
rect 2652 -186 2658 -175
rect 2710 -186 2716 -134
rect 2856 -681 2890 48
rect 3272 -681 3306 724
rect 2856 -715 3307 -681
rect 2492 -949 2501 -854
rect 2596 -949 2605 -854
rect 2856 -1103 2890 -715
rect 3272 -883 3306 -715
rect 3272 -917 3603 -883
rect 3273 -918 3307 -917
rect 3387 -945 3461 -917
rect 3387 -951 3459 -945
rect 3387 -1020 3390 -951
rect 3459 -1020 3461 -991
rect 3569 -1020 3603 -917
rect 3387 -1025 3461 -1020
rect 3390 -1029 3459 -1025
rect 3552 -1029 3621 -1020
rect 2855 -1177 2890 -1103
rect 3552 -1107 3621 -1098
rect 2855 -1178 2961 -1177
rect 4242 -1178 4251 -1167
rect 2855 -1212 4251 -1178
rect 2855 -1215 2997 -1212
rect 4242 -1223 4251 -1212
rect 4310 -1223 4319 -1167
<< via2 >>
rect 2501 -949 2596 -854
rect 3390 -1020 3459 -951
rect 3552 -1098 3621 -1029
rect 4251 -1223 4310 -1167
<< metal3 >>
rect 2496 -854 2601 -849
rect 2496 -925 2501 -854
rect 2494 -949 2501 -925
rect 2596 -925 2601 -854
rect 2596 -949 2603 -925
rect 2494 -1030 2603 -949
rect 3380 -951 3475 -940
rect 3380 -1020 3390 -951
rect 3459 -1020 3475 -951
rect 3380 -1096 3475 -1020
rect 3547 -1026 3626 -1024
rect 3547 -1029 3704 -1026
rect 3547 -1098 3552 -1029
rect 3621 -1098 3841 -1029
rect 3547 -1103 3841 -1098
rect 3548 -1124 3841 -1103
rect 3380 -1175 3475 -1169
rect 4246 -1167 4315 -1162
rect 4246 -1223 4251 -1167
rect 4310 -1223 4315 -1167
rect 4246 -1393 4315 -1223
rect 4229 -1399 4333 -1393
rect 4229 -1509 4333 -1503
<< via3 >>
rect 3380 -1169 3475 -1096
rect 4229 -1503 4333 -1399
<< metal4 >>
rect 3124 -1096 3476 -1095
rect 3124 -1168 3380 -1096
rect 3379 -1169 3380 -1168
rect 3475 -1169 3476 -1096
rect 3379 -1170 3476 -1169
rect 4228 -1399 4334 -1398
rect 4228 -1430 4229 -1399
rect 4156 -1461 4229 -1430
rect 3944 -1503 4229 -1461
rect 4333 -1503 4334 -1399
rect 3944 -1534 4334 -1503
use sky130_fd_pr__nfet_01v8_69TQ3K  XM1 ~/Desktop/ASIC_ADC/magic/th01
timestamp 1704730646
transform 1 0 2252 0 1 274
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_3HMWVM  XM2 ~/Desktop/ASIC_ADC/magic/th01
timestamp 1704730646
transform 1 0 1664 0 1 935
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_69TQ3K  XM3
timestamp 1704730646
transform 1 0 1666 0 1 272
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_3HMWVM  XM4
timestamp 1704730646
transform 1 0 2248 0 1 935
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_3HMWVM  XM5
timestamp 1704730646
transform 1 0 818 0 1 939
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_PSFW3M  XM6 ~/Desktop/ASIC_ADC/magic/th01
timestamp 1704730646
transform 1 0 2758 0 1 274
box -226 -310 226 310
use sky130_fd_pr__pfet_01v8_3HMWVM  XM7
timestamp 1704730646
transform 1 0 3102 0 1 933
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_69TQ3K  XM8
timestamp 1704730646
transform 1 0 3270 0 1 274
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_3HMWVM  XM9
timestamp 1704730646
transform 1 0 240 0 1 939
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_69TQ3K  XM10
timestamp 1704730646
transform 1 0 834 0 1 272
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_69TQ3K  XM11
timestamp 1704730646
transform 1 0 242 0 1 272
box -296 -310 296 310
use sky130_fd_pr__res_xhigh_po_0p35_FM7VE8  XR1 ~/Desktop/ASIC_ADC/magic/th01
timestamp 1704730646
transform 0 -1 2046 1 0 -671
box -201 -2098 201 2098
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR2
timestamp 1704748838
transform 0 -1 1046 1 0 -249
box -201 -1098 201 1098
use sky130_fd_pr__res_xhigh_po_0p35_FM7VE8  XR3
timestamp 1704730646
transform 0 -1 2044 1 0 1485
box -201 -2098 201 2098
<< labels >>
flabel metal1 2338 1486 2538 1686 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 1054 -40 1254 160 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 2548 614 2748 814 0 FreeSans 256 0 0 0 vin
port 1 nsew
flabel metal1 3370 588 3570 788 0 FreeSans 256 0 0 0 Vout
port 2 nsew
<< end >>
