* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : inv03f                                       *
* Netlisted  : Sun Dec  1 20:08:24 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733080094010                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733080094010 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=2.95e-07 W=7.65e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733080094010

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733080094011                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733080094011 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=3.45e-07 W=6.3e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733080094011

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv03f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv03f A VDD VSS Y
** N=9 EP=4 FDC=2
X2 VSS Y A nfet_01v8_CDNS_733080094010 $T=365 640 0 0 $X=-40 $Y=490
X3 VDD Y A pfet_01v8_CDNS_733080094011 $T=335 2845 0 0 $X=-110 $Y=2665
.ends inv03f
