* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : inv03f                                       *
* Netlisted  : Mon Nov 18 14:04:23 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv03f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv03f
** N=4 EP=0 FDC=0
.ends inv03f
