magic
tech sky130A
magscale 1 2
timestamp 1706392731
<< metal1 >>
rect 3737 593 9365 627
rect 3737 -889 3771 593
rect 4191 571 4219 593
rect 9211 567 9353 593
rect 9285 555 9353 567
rect 9420 526 9620 626
rect 5899 456 5933 457
rect 5858 404 5864 456
rect 5916 404 5933 456
rect 5877 391 5933 404
rect 5877 357 6005 391
rect 5877 305 5911 357
rect 6772 324 6778 376
rect 6830 324 6836 376
rect 5583 151 5617 261
rect 6781 229 6828 324
rect 5583 117 5655 151
rect 5621 46 5655 117
rect 5612 -154 5712 46
rect 8382 -40 8434 -34
rect 8291 -83 8382 -49
rect 8382 -98 8434 -92
rect 6882 -113 7082 -98
rect 6882 -147 7279 -113
rect 6882 -198 7082 -147
rect 8576 -164 8676 36
rect 5578 -257 5785 -220
rect 8656 -402 8828 -340
rect 4474 -799 4574 -674
rect 5150 -771 5350 -750
rect 5748 -752 5785 -418
rect 8628 -440 8828 -402
rect 7375 -752 7409 -615
rect 8654 -752 8688 -440
rect 9740 -624 9940 -524
rect 4335 -833 4574 -799
rect 3737 -923 3817 -889
rect 4335 -901 4369 -833
rect 4474 -874 4574 -833
rect 4911 -776 5350 -771
rect 5400 -776 10185 -752
rect 4911 -805 10185 -776
rect 4911 -851 4945 -805
rect 5150 -823 10185 -805
rect 5150 -850 5350 -823
rect 5400 -848 10185 -823
rect 3783 -1181 3817 -923
rect 3769 -2666 3803 -1191
rect 4014 -2206 4214 -2106
rect 4959 -2219 4993 -1021
rect 3721 -2745 3755 -2711
rect 3789 -2745 3803 -2666
<< via1 >>
rect 5864 404 5916 456
rect 6778 324 6830 376
rect 8382 -92 8434 -40
<< metal2 >>
rect 3847 775 6055 809
rect 3847 -597 3881 775
rect 6021 726 6055 775
rect 3948 676 5912 720
rect 6021 692 10056 726
rect 3948 -488 3992 676
rect 5868 462 5912 676
rect 5864 456 5916 462
rect 5864 398 5916 404
rect 6787 382 6821 692
rect 6778 376 6830 382
rect 6778 318 6830 324
rect 8391 -40 8425 692
rect 10021 213 10055 692
rect 8376 -92 8382 -40
rect 8434 -92 8440 -40
rect 3948 -532 4140 -488
rect 3657 -631 3881 -597
rect 3657 -1707 3691 -631
rect 4125 -1707 4159 -1589
rect 3657 -1741 4159 -1707
rect 3657 -3445 3691 -1741
rect 4059 -3445 4093 -3347
rect 3657 -3479 4093 -3445
rect 3657 -3483 3691 -3479
use preamp  preamp_0
timestamp 1706271137
transform -1 0 7242 0 1 -714
box 394 136 1494 1340
use th09  th09_0
timestamp 1706236419
transform -1 0 8710 0 1 104
box 368 -754 1692 526
use th10  th10_0
timestamp 1706270854
transform 0 -1 4222 1 0 -1906
box 270 -794 1168 452
use th12  th12_0
timestamp 1706270854
transform 0 -1 3916 1 0 -3690
box 278 -1078 1572 236
use th13  th13_0
timestamp 1706270854
transform -1 0 10614 0 1 -20
box 438 -680 2042 646
use th15  th15_0
timestamp 1706388900
transform 1 0 3594 0 1 -46
box 468 -522 2070 674
<< labels >>
flabel metal1 9420 526 9620 626 0 FreeSans 256 0 0 0 Vp
port 1 nsew
flabel metal1 9740 -624 9940 -524 0 FreeSans 256 0 0 0 Vin
port 0 nsew
flabel metal1 8576 -164 8676 36 0 FreeSans 256 270 0 0 V13
port 14 nsew
flabel metal1 6882 -198 7082 -98 0 FreeSans 256 180 0 0 V09
port 10 nsew
flabel metal1 5612 -154 5712 46 0 FreeSans 256 90 0 0 V15
port 16 nsew
flabel metal1 5150 -850 5350 -750 0 FreeSans 256 180 0 0 Vn
port 17 nsew
flabel metal1 4474 -874 4574 -674 0 FreeSans 256 90 0 0 V10
port 11 nsew
flabel metal1 4014 -2206 4214 -2106 0 FreeSans 256 0 0 0 V12
port 13 nsew
<< end >>
