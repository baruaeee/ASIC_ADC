magic
tech sky130A
magscale 1 2
timestamp 1706323418
<< metal1 >>
rect 22568 7996 22620 8002
rect 22568 7938 22620 7944
rect 25332 7922 25384 7928
rect 25332 7864 25384 7870
rect 24194 7849 24246 7855
rect 24194 7791 24246 7797
rect 22454 7456 22490 7522
rect 22454 7420 22588 7456
rect 22516 7396 22588 7420
rect 22552 7160 22588 7396
rect 25762 7157 25796 7556
rect 22159 6418 22211 6424
rect 22159 6357 22211 6363
rect 22351 6009 22497 6043
rect 22351 5835 22385 6009
rect 22063 5801 22385 5835
rect 22154 5176 22480 5204
rect 22154 5040 22182 5176
rect 22346 4928 22561 4976
rect 22346 4256 22394 4928
rect 22188 4208 22394 4256
rect 22072 3892 22124 3898
rect 22072 3834 22124 3840
rect 22037 3133 22351 3167
rect 22317 2797 22351 3133
rect 22317 2763 22505 2797
<< via1 >>
rect 22568 7944 22620 7996
rect 25332 7870 25384 7922
rect 24194 7797 24246 7849
rect 22159 6363 22211 6418
rect 22072 3840 22124 3892
<< metal2 >>
rect 22562 7944 22568 7996
rect 22620 7944 22706 7996
rect 25326 7870 25332 7922
rect 25384 7913 25390 7922
rect 25384 7879 25447 7913
rect 25384 7870 25390 7879
rect 24188 7843 24194 7849
rect 24000 7802 24194 7843
rect 24188 7797 24194 7802
rect 24246 7797 24252 7849
rect 22210 6418 22266 6427
rect 22153 6363 22159 6418
rect 22210 6353 22266 6362
rect 22190 3892 22246 3901
rect 22066 3840 22072 3892
rect 22124 3880 22130 3892
rect 22124 3852 22190 3880
rect 22124 3840 22130 3852
rect 22190 3827 22246 3836
<< via2 >>
rect 22210 6363 22211 6418
rect 22211 6363 22266 6418
rect 22210 6362 22266 6363
rect 22190 3836 22246 3892
<< metal3 >>
rect 22354 6758 22468 6818
rect 22205 6420 22271 6423
rect 22354 6420 22414 6758
rect 22205 6418 22414 6420
rect 22205 6362 22210 6418
rect 22266 6362 22414 6418
rect 22205 6360 22414 6362
rect 22205 6357 22271 6360
rect 22185 3894 22251 3897
rect 22314 3894 22374 4158
rect 22185 3892 22374 3894
rect 22185 3836 22190 3892
rect 22246 3836 22374 3892
rect 22185 3834 22374 3836
rect 22185 3831 22251 3834
use therm  therm_0
timestamp 1706321462
transform 1 0 21385 0 1 600
box -1 1094 7123 7902
use Analog  x1
timestamp 1706323418
transform 1 0 0 0 1 7400
box 20556 -6558 28914 1285
<< end >>
