** sch_path: /home/exotic/Desktop/ASIC_ADC/xschem/Vth_sch/test_logic_1.sch
**.subckt test_logic_1 b[3],b[2],b[1],b[0]
*.opin b[3],b[2],b[1],b[0]
VDD VDD GND 1.8
V0 p0 GND pulse(0.45 1.3 10ns 1ns 1ns 150ns)
V1 p1 GND pulse(0.45 1.3 20ns 1ns 1ns 140ns)
V2 p2 GND pulse(0.45 1.3 30ns 1ns 1ns 130ns)
V3 p3 GND pulse(0.45 1.3 40ns 1ns 1ns 120ns)
V4 p4 GND pulse(0.45 1.3 50ns 1ns 1ns 110ns)
V5 p5 GND pulse(0.45 1.3 60ns 1ns 1ns 100ns)
V6 p6 GND pulse(0.45 1.3 70ns 1ns 1ns 90ns)
V7 p7 GND pulse(0.45 1.3 70ns 1ns 1ns 90ns)
V8 p8 GND pulse(0.45 1.3 80ns 1ns 1ns 80ns)
V9 p9 GND pulse(0.45 1.3 90ns 1ns 1ns 70ns)
V10 p10 GND pulse(0.45 1.3 100ns 1ns 1ns 60ns)
V11 p11 GND pulse(0.45 1.3 110ns 1ns 1ns 50ns)
V12 p12 GND pulse(0.45 1.3 120ns 1ns 1ns 40ns)
V13 p13 GND pulse(0.45 1.3 130ns 1ns 1ns 30ns)
V14 p14 GND pulse(0.45 1.3 140ns 1ns 1ns 10ns)
x1 GND VDD pb[0] b[1] b[2] b[3] p0 p10 p11 p12 p13 p14 p1 p2 p3 p4 p5 p6 p7 p8 p9 therm


**** begin user architecture code


*vvpwr vpwr 0 dc 1.8
*vvgnd vgnd 0 dc 0
*.dc Vin 0 1.8 0.01
.tran 1n 160n
.control
run
*set color0=white
*set color1=black
*plot Vin Vout V_LH V_LL
plot p0 p1 p2 p3 p4 p5 p6 p7 p8 p9 p10 p11 p12 p13 p14
set xbrushwidth=3
*.save all
.endc
.end


 .lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
*.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* NGSPICE file created from therm.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X a_208_47# a_75_199#
+ a_544_297# a_315_47# a_201_297#
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VGND a_315_47# 0.00427f
C1 a_201_297# a_75_199# 0.16f
C2 A2 VGND 0.0119f
C3 A3 a_208_47# 3.65e-19
C4 a_201_297# A1 0.011f
C5 X VGND 0.0609f
C6 a_75_199# A1 0.0696f
C7 VPWR VGND 0.0735f
C8 a_544_297# VGND 0.00256f
C9 a_201_297# B1 0.00594f
C10 VPB VGND 0.00772f
C11 a_208_47# a_75_199# 0.0159f
C12 a_201_297# C1 0.00243f
C13 a_75_199# B1 0.102f
C14 A3 A2 0.0747f
C15 a_75_199# C1 0.0628f
C16 A1 B1 0.0716f
C17 a_75_199# a_315_47# 0.0202f
C18 a_201_297# A2 0.0112f
C19 A3 X 0.00317f
C20 C1 A1 3.21e-19
C21 A3 VPWR 0.0181f
C22 VPB A3 0.0268f
C23 a_75_199# A2 0.0621f
C24 A1 a_315_47# 0.00313f
C25 a_201_297# X 0.0131f
C26 C1 B1 0.066f
C27 a_201_297# VPWR 0.211f
C28 a_544_297# a_201_297# 0.00702f
C29 VPB a_201_297# 0.00186f
C30 a_75_199# X 0.0959f
C31 A2 A1 0.0689f
C32 a_75_199# VPWR 0.109f
C33 a_544_297# a_75_199# 0.0176f
C34 VPB a_75_199# 0.0486f
C35 a_208_47# A2 0.00102f
C36 X A1 1.2e-19
C37 A3 VGND 0.0161f
C38 VPWR A1 0.0151f
C39 VPB A1 0.0306f
C40 a_208_47# X 1.91e-19
C41 a_208_47# VPWR 8.35e-19
C42 X B1 7.79e-20
C43 a_201_297# VGND 0.00403f
C44 A2 a_315_47# 0.00335f
C45 VPWR B1 0.0125f
C46 a_544_297# B1 1.13e-19
C47 VPB B1 0.0292f
C48 C1 X 5.14e-20
C49 a_75_199# VGND 0.362f
C50 C1 VPWR 0.0146f
C51 VPB C1 0.0394f
C52 VPWR a_315_47# 0.00154f
C53 VGND A1 0.0113f
C54 X A2 3.01e-19
C55 a_208_47# VGND 0.00302f
C56 A2 VPWR 0.0174f
C57 VPB A2 0.0376f
C58 A3 a_201_297# 0.00642f
C59 VGND B1 0.0171f
C60 A3 a_75_199# 0.163f
C61 X VPWR 0.0676f
C62 C1 VGND 0.0181f
C63 a_544_297# X 2.35e-19
C64 VPB X 0.0107f
C65 a_544_297# VPWR 0.0105f
C66 VPB VPWR 0.0749f
C67 VGND VNB 0.437f
C68 VPWR VNB 0.365f
C69 X VNB 0.0906f
C70 C1 VNB 0.148f
C71 B1 VNB 0.0947f
C72 A1 VNB 0.101f
C73 A2 VNB 0.11f
C74 A3 VNB 0.0908f
C75 VPB VNB 0.782f
C76 a_201_297# VNB 0.00345f
C77 a_75_199# VNB 0.205f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_181_47# a_109_47# a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPWR X 0.0766f
C1 A a_109_47# 6.45e-19
C2 a_27_47# VPWR 0.145f
C3 VPB VPWR 0.0795f
C4 B VPWR 0.128f
C5 VGND VPWR 0.0475f
C6 A a_27_47# 0.157f
C7 A VPB 0.0426f
C8 C a_181_47# 0.00151f
C9 A B 0.0869f
C10 VGND A 0.0154f
C11 C X 0.0149f
C12 a_27_47# a_109_47# 0.00517f
C13 C a_27_47# 0.186f
C14 a_27_47# a_181_47# 0.00401f
C15 A VPWR 0.0185f
C16 VGND a_109_47# 0.00123f
C17 C VPB 0.0347f
C18 C B 0.0746f
C19 VGND C 0.0703f
C20 a_27_47# X 0.087f
C21 VGND a_181_47# 0.00261f
C22 VPB X 0.0121f
C23 B X 0.00111f
C24 VGND X 0.0708f
C25 VPWR a_109_47# 3.29e-19
C26 VPB a_27_47# 0.0501f
C27 C VPWR 0.00464f
C28 a_27_47# B 0.0625f
C29 VGND a_27_47# 0.134f
C30 VPWR a_181_47# 3.97e-19
C31 VPB B 0.0836f
C32 VGND VPB 0.00604f
C33 VGND B 0.00714f
C34 VGND VNB 0.3f
C35 X VNB 0.0923f
C36 C VNB 0.12f
C37 A VNB 0.174f
C38 VPWR VNB 0.274f
C39 B VNB 0.102f
C40 VPB VNB 0.516f
C41 a_27_47# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
C0 VGND VPWR 0.353f
C1 VGND VPB 0.0797f
C2 VPWR VPB 0.0625f
C3 VPWR VNB 0.47f
C4 VGND VNB 0.427f
C5 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VGND VPWR 0.546f
C1 VGND VPB 0.116f
C2 VPWR VPB 0.0787f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_384_47# a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
C0 a_299_297# VPB 0.0111f
C1 VGND VPWR 0.0579f
C2 A2 VPWR 0.0201f
C3 a_81_21# a_299_297# 0.0821f
C4 VGND A2 0.0495f
C5 B1 a_299_297# 0.00863f
C6 A1 a_299_297# 0.0585f
C7 VPWR VPB 0.068f
C8 X VPWR 0.0847f
C9 VGND VPB 0.00713f
C10 a_384_47# a_81_21# 0.00138f
C11 A1 a_384_47# 0.00884f
C12 A2 VPB 0.0373f
C13 VGND X 0.0512f
C14 a_81_21# VPWR 0.146f
C15 B1 VPWR 0.0196f
C16 A1 VPWR 0.0209f
C17 VGND a_81_21# 0.173f
C18 B1 VGND 0.0181f
C19 A1 VGND 0.0786f
C20 a_384_47# a_299_297# 1.48e-19
C21 a_81_21# A2 7.47e-19
C22 A1 A2 0.0921f
C23 a_299_297# VPWR 0.202f
C24 X VPB 0.0108f
C25 VGND a_299_297# 0.00772f
C26 a_81_21# VPB 0.0593f
C27 B1 VPB 0.0387f
C28 a_299_297# A2 0.0468f
C29 A1 VPB 0.0264f
C30 X a_81_21# 0.112f
C31 B1 X 3.04e-20
C32 a_384_47# VPWR 4.08e-19
C33 VGND a_384_47# 0.00366f
C34 B1 a_81_21# 0.148f
C35 A1 a_81_21# 0.0568f
C36 B1 A1 0.0817f
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 VPWR VGND 0.0423f
C1 Y VGND 0.155f
C2 VPB VGND 0.00649f
C3 A VGND 0.0638f
C4 Y VPWR 0.209f
C5 VPB VPWR 0.0521f
C6 A VPWR 0.0631f
C7 VPB Y 0.0061f
C8 A Y 0.0894f
C9 VPB A 0.0742f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X a_29_53# a_183_297# a_111_297#
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 B VPWR 0.147f
C1 C VPWR 0.00457f
C2 X a_29_53# 0.0991f
C3 B C 0.0802f
C4 X VGND 0.036f
C5 X VPB 0.0109f
C6 VPWR a_29_53# 0.0833f
C7 VGND VPWR 0.0459f
C8 VPB VPWR 0.0649f
C9 B a_29_53# 0.121f
C10 X A 0.00127f
C11 B VGND 0.0152f
C12 B VPB 0.0962f
C13 A VPWR 0.00936f
C14 a_111_297# VPWR 5.94e-19
C15 C a_29_53# 0.0857f
C16 a_183_297# VPWR 8.13e-19
C17 C VGND 0.0161f
C18 C VPB 0.0396f
C19 B A 0.0787f
C20 C A 0.0343f
C21 VGND a_29_53# 0.217f
C22 VPB a_29_53# 0.0491f
C23 VPB VGND 0.00724f
C24 A a_29_53# 0.242f
C25 a_111_297# a_29_53# 0.005f
C26 a_183_297# a_29_53# 0.00868f
C27 A VGND 0.0187f
C28 a_111_297# VGND 3.96e-19
C29 a_183_297# VGND 5.75e-19
C30 VPB A 0.0377f
C31 X VPWR 0.0885f
C32 B X 6.52e-19
C33 a_111_297# A 0.00223f
C34 a_183_297# A 0.00239f
C35 VGND VNB 0.306f
C36 X VNB 0.0882f
C37 A VNB 0.117f
C38 C VNB 0.16f
C39 B VNB 0.117f
C40 VPWR VNB 0.253f
C41 VPB VNB 0.516f
C42 a_29_53# VNB 0.18f
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 Y VGND 0.154f
C1 Y B 0.0877f
C2 VPB VGND 0.00456f
C3 VPB B 0.0367f
C4 Y VPWR 0.0995f
C5 Y a_109_297# 0.0113f
C6 B VGND 0.0451f
C7 Y A 0.0471f
C8 VPB VPWR 0.0449f
C9 VPWR VGND 0.0314f
C10 a_109_297# VGND 0.00128f
C11 B VPWR 0.0148f
C12 VPB A 0.0415f
C13 A VGND 0.0486f
C14 B A 0.0584f
C15 a_109_297# VPWR 0.00638f
C16 A VPWR 0.0528f
C17 VPB Y 0.0139f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
C0 VPB VPWR 0.0858f
C1 VPB VGND 0.161f
C2 VGND VPWR 0.903f
C3 VPWR VNB 0.867f
C4 VGND VNB 0.761f
C5 VPB VNB 0.605f
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X a_193_297# a_465_47#
+ a_205_47# a_109_297# a_27_47#
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
C0 A1 B1 0.0609f
C1 A1 A2 0.0692f
C2 a_109_297# C1 0.00739f
C3 a_109_297# VPWR 0.15f
C4 C1 B1 6.46e-19
C5 C1 A2 9.03e-21
C6 VPWR B1 0.00982f
C7 VPWR A2 0.0209f
C8 a_109_297# X 3.99e-19
C9 A1 C1 1.77e-20
C10 a_109_297# a_193_297# 0.0927f
C11 A1 VPWR 0.0161f
C12 a_109_297# B2 0.0133f
C13 X B1 9.58e-20
C14 X A2 0.00157f
C15 VPWR a_205_47# 1.62e-19
C16 a_193_297# B1 0.00869f
C17 A2 a_193_297# 0.00683f
C18 A1 X 2.77e-19
C19 B2 B1 0.0784f
C20 A1 a_465_47# 7.06e-19
C21 VPWR C1 0.0139f
C22 a_109_297# a_27_47# 0.0961f
C23 VGND a_109_297# 0.00284f
C24 VPB a_109_297# 0.00421f
C25 A1 a_193_297# 0.0109f
C26 X C1 5.03e-20
C27 a_27_47# B1 0.112f
C28 A2 a_27_47# 0.153f
C29 VGND B1 0.0133f
C30 VGND A2 0.0168f
C31 VPB B1 0.0321f
C32 VPB A2 0.027f
C33 VPWR X 0.0897f
C34 VPWR a_465_47# 5.05e-19
C35 C1 B2 0.0726f
C36 A1 a_27_47# 0.0984f
C37 VGND A1 0.0126f
C38 VPB A1 0.0343f
C39 VPWR a_193_297# 0.169f
C40 VPWR B2 0.00842f
C41 a_27_47# a_205_47# 0.00762f
C42 VGND a_205_47# 0.00156f
C43 X a_465_47# 1.56e-19
C44 C1 a_27_47# 0.0792f
C45 VGND C1 0.0196f
C46 X a_193_297# 0.00367f
C47 VPB C1 0.0367f
C48 X B2 6.77e-20
C49 VPWR a_27_47# 0.099f
C50 VGND VPWR 0.0722f
C51 VPB VPWR 0.0799f
C52 B2 a_193_297# 0.00126f
C53 X a_27_47# 0.0921f
C54 VGND X 0.061f
C55 a_27_47# a_465_47# 0.013f
C56 VGND a_465_47# 0.00257f
C57 VPB X 0.0113f
C58 a_27_47# a_193_297# 0.144f
C59 VGND a_193_297# 0.00438f
C60 VPB a_193_297# 0.00774f
C61 B2 a_27_47# 0.0959f
C62 VGND B2 0.0174f
C63 VPB B2 0.0256f
C64 a_109_297# B1 0.00736f
C65 A1 a_109_297# 1.05e-19
C66 VGND a_27_47# 0.395f
C67 VPB a_27_47# 0.0512f
C68 VGND VPB 0.00844f
C69 VGND VNB 0.437f
C70 X VNB 0.0919f
C71 VPWR VNB 0.364f
C72 A2 VNB 0.0896f
C73 A1 VNB 0.106f
C74 B1 VNB 0.108f
C75 B2 VNB 0.0887f
C76 C1 VNB 0.139f
C77 VPB VNB 0.782f
C78 a_193_297# VNB 0.0011f
C79 a_109_297# VNB 7.11e-19
C80 a_27_47# VNB 0.216f
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X a_256_47# a_584_47#
+ a_93_21# a_250_297# a_346_47#
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
C0 A1 B2 3.14e-19
C1 B2 a_250_297# 0.0344f
C2 A3 a_250_297# 0.00602f
C3 a_584_47# a_250_297# 2.43e-19
C4 A1 X 6.03e-20
C5 a_256_47# A3 4.42e-19
C6 A1 B1 0.0965f
C7 A1 a_93_21# 0.0641f
C8 A3 B2 9.12e-20
C9 a_250_297# X 5.42e-19
C10 B1 a_250_297# 0.0125f
C11 a_346_47# B1 5.39e-20
C12 a_93_21# a_250_297# 0.188f
C13 a_346_47# a_93_21# 0.0119f
C14 A1 A2 0.0971f
C15 VPWR A1 0.016f
C16 VPB A1 0.0296f
C17 VGND A1 0.0133f
C18 a_256_47# B1 2.07e-20
C19 a_256_47# a_93_21# 0.0114f
C20 A2 a_250_297# 0.0129f
C21 B1 B2 0.0823f
C22 a_346_47# A2 0.00252f
C23 VPWR a_250_297# 0.313f
C24 A3 X 2.45e-19
C25 VPWR a_346_47# 0.00109f
C26 VPB a_250_297# 0.00616f
C27 VGND a_250_297# 0.0072f
C28 VGND a_346_47# 0.00514f
C29 a_93_21# B2 0.0147f
C30 A3 B1 7.88e-22
C31 A3 a_93_21# 0.124f
C32 a_256_47# A2 0.00256f
C33 VPWR a_256_47# 9.47e-19
C34 VGND a_256_47# 0.00394f
C35 a_584_47# B1 0.00143f
C36 a_584_47# a_93_21# 0.00278f
C37 A2 B2 1.46e-19
C38 VPWR B2 0.0108f
C39 VPB B2 0.0355f
C40 VGND B2 0.0469f
C41 A3 A2 0.0788f
C42 VPWR A3 0.0158f
C43 VPB A3 0.0291f
C44 VGND A3 0.00974f
C45 B1 X 3.83e-20
C46 a_93_21# X 0.0841f
C47 VPWR a_584_47# 9.47e-19
C48 VGND a_584_47# 0.00683f
C49 a_93_21# B1 0.0774f
C50 A2 X 1.19e-19
C51 VPWR X 0.0849f
C52 VPB X 0.0108f
C53 VGND X 0.06f
C54 A2 B1 1.44e-20
C55 VPWR B1 0.01f
C56 VPB B1 0.0276f
C57 VGND B1 0.0344f
C58 a_93_21# A2 0.0747f
C59 VPWR a_93_21# 0.0907f
C60 VPB a_93_21# 0.0485f
C61 VGND a_93_21# 0.251f
C62 A1 a_250_297# 0.0129f
C63 A1 a_346_47# 0.00465f
C64 VPWR A2 0.0133f
C65 VPB A2 0.0287f
C66 VPWR VPB 0.0756f
C67 VGND A2 0.0114f
C68 VPWR VGND 0.076f
C69 VPB VGND 0.00788f
C70 VGND VNB 0.465f
C71 VPWR VNB 0.365f
C72 X VNB 0.0937f
C73 B2 VNB 0.14f
C74 B1 VNB 0.101f
C75 A1 VNB 0.0951f
C76 A2 VNB 0.0921f
C77 A3 VNB 0.0929f
C78 VPB VNB 0.782f
C79 a_250_297# VNB 0.0278f
C80 a_93_21# VNB 0.151f
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X a_277_297# a_205_297# a_27_297#
+ a_109_297#
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 A C 0.028f
C1 A X 0.00133f
C2 a_277_297# C 5.54e-19
C3 X a_277_297# 6.43e-20
C4 a_109_297# VGND 7.58e-19
C5 B C 0.0917f
C6 B X 6.42e-19
C7 A a_277_297# 2.28e-19
C8 VGND C 0.0191f
C9 VGND X 0.0354f
C10 A B 0.0639f
C11 A VGND 0.016f
C12 B a_277_297# 2.29e-19
C13 VGND a_277_297# 4.65e-19
C14 a_205_297# C 0.00261f
C15 D C 0.0954f
C16 VGND B 0.0159f
C17 a_109_297# a_27_297# 0.00695f
C18 VPWR a_109_297# 9.23e-19
C19 A D 2.13e-19
C20 a_27_297# C 0.158f
C21 X a_27_297# 0.0991f
C22 VPB C 0.0338f
C23 VPB X 0.0109f
C24 VPWR C 0.00723f
C25 VPWR X 0.0878f
C26 B D 0.00287f
C27 A a_27_297# 0.163f
C28 VPB A 0.033f
C29 VPWR A 0.00769f
C30 VGND a_205_297# 3.36e-19
C31 VGND D 0.0517f
C32 a_27_297# a_277_297# 0.00876f
C33 VPWR a_277_297# 7.48e-19
C34 B a_27_297# 0.159f
C35 VPB B 0.106f
C36 VPWR B 0.193f
C37 VGND a_27_297# 0.235f
C38 VPB VGND 0.00796f
C39 VPWR VGND 0.0546f
C40 a_27_297# a_205_297# 0.00412f
C41 VPWR a_205_297# 5.16e-19
C42 D a_27_297# 0.054f
C43 VPB D 0.0405f
C44 VPWR D 0.00503f
C45 a_109_297# C 0.00356f
C46 VPB a_27_297# 0.0517f
C47 VPWR a_27_297# 0.084f
C48 VPB VPWR 0.075f
C49 VGND VNB 0.367f
C50 X VNB 0.0883f
C51 A VNB 0.109f
C52 C VNB 0.105f
C53 D VNB 0.175f
C54 B VNB 0.115f
C55 VPWR VNB 0.29f
C56 VPB VNB 0.605f
C57 a_27_297# VNB 0.163f
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
C0 VPB VPWR 0.137f
C1 VGND VPWR 1.57f
C2 VPB VGND 0.35f
C3 VPWR VNB 1.67f
C4 VGND VNB 1.47f
C5 VPB VNB 1.14f
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X a_369_47# a_469_47#
+ a_297_47# a_193_413# a_27_47#
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
C0 C VPWR 0.0182f
C1 C a_193_413# 0.0389f
C2 VPWR a_369_47# 6.65e-19
C3 C VPB 0.0742f
C4 a_193_413# a_369_47# 0.00181f
C5 a_469_47# VPWR 7.77e-19
C6 C VGND 0.0395f
C7 C X 0.00479f
C8 a_469_47# a_193_413# 0.00109f
C9 C D 0.183f
C10 a_193_413# VPWR 0.281f
C11 VGND a_369_47# 0.00505f
C12 VPB VPWR 0.0818f
C13 a_469_47# VGND 0.00551f
C14 a_469_47# X 0.001f
C15 VPB a_193_413# 0.0644f
C16 C B 0.164f
C17 a_469_47# D 0.00183f
C18 VGND VPWR 0.0727f
C19 VPWR X 0.0586f
C20 B a_369_47# 0.00129f
C21 D VPWR 0.0186f
C22 a_193_413# VGND 0.0915f
C23 a_193_413# X 0.108f
C24 a_297_47# VPWR 2.82e-19
C25 VPB VGND 0.0123f
C26 a_193_413# D 0.155f
C27 VPB X 0.0108f
C28 a_193_413# a_297_47# 0.00137f
C29 VPB D 0.0763f
C30 B VPWR 0.0186f
C31 A_N VPWR 0.02f
C32 a_27_47# VPWR 0.106f
C33 VGND X 0.0588f
C34 a_193_413# B 0.144f
C35 A_N a_193_413# 0.00151f
C36 D VGND 0.0372f
C37 a_27_47# a_193_413# 0.125f
C38 D X 0.0168f
C39 a_297_47# VGND 0.00183f
C40 VPB B 0.089f
C41 A_N VPB 0.0832f
C42 a_27_47# VPB 0.092f
C43 B VGND 0.037f
C44 A_N VGND 0.0205f
C45 a_27_47# VGND 0.103f
C46 a_297_47# B 0.00353f
C47 C a_369_47# 0.00448f
C48 a_469_47# C 0.00202f
C49 a_27_47# B 0.0794f
C50 A_N a_27_47# 0.237f
C51 VGND VNB 0.456f
C52 X VNB 0.0934f
C53 VPWR VNB 0.368f
C54 D VNB 0.123f
C55 C VNB 0.108f
C56 B VNB 0.12f
C57 A_N VNB 0.198f
C58 VPB VNB 0.782f
C59 a_193_413# VNB 0.136f
C60 a_27_47# VNB 0.224f
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X a_109_93# a_368_53# a_209_311#
+ a_296_53#
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
C0 a_296_53# VPWR 1.15e-19
C1 C VGND 0.0678f
C2 VPWR VGND 0.0657f
C3 A_N VGND 0.045f
C4 VGND VPB 0.00909f
C5 a_368_53# VGND 0.0031f
C6 X VGND 0.0647f
C7 VPWR C 0.005f
C8 a_296_53# a_209_311# 0.0049f
C9 a_109_93# a_296_53# 1.84e-19
C10 a_209_311# VGND 0.131f
C11 C A_N 7.6e-19
C12 a_109_93# VGND 0.0784f
C13 C VPB 0.0339f
C14 B VGND 0.00796f
C15 VPWR A_N 0.0513f
C16 C a_368_53# 0.00415f
C17 VPWR VPB 0.104f
C18 C X 0.0176f
C19 VPWR a_368_53# 4.26e-19
C20 VPWR X 0.0732f
C21 A_N VPB 0.111f
C22 C a_209_311# 0.19f
C23 a_109_93# C 3.91e-20
C24 B C 0.0671f
C25 X A_N 1.44e-19
C26 X VPB 0.0119f
C27 VPWR a_209_311# 0.155f
C28 a_109_93# VPWR 0.0984f
C29 B VPWR 0.131f
C30 a_209_311# A_N 0.00515f
C31 a_209_311# VPB 0.0515f
C32 a_109_93# A_N 0.117f
C33 a_109_93# VPB 0.0652f
C34 B A_N 2.03e-19
C35 B VPB 0.0914f
C36 a_209_311# a_368_53# 0.0026f
C37 X a_209_311# 0.0877f
C38 B X 0.00119f
C39 a_296_53# VGND 6.07e-19
C40 a_109_93# a_209_311# 0.168f
C41 B a_209_311# 0.0609f
C42 a_109_93# B 0.0802f
C43 VGND VNB 0.44f
C44 X VNB 0.0925f
C45 C VNB 0.114f
C46 B VNB 0.101f
C47 VPWR VNB 0.342f
C48 A_N VNB 0.197f
C49 VPB VNB 0.693f
C50 a_209_311# VNB 0.143f
C51 a_109_93# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
C0 X VPWR 0.317f
C1 X VGND 0.216f
C2 VPB VPWR 0.0632f
C3 VPB VGND 0.00583f
C4 a_27_47# VPWR 0.219f
C5 a_27_47# VGND 0.148f
C6 X VPB 0.0122f
C7 X a_27_47# 0.328f
C8 A VPWR 0.022f
C9 VGND A 0.0431f
C10 a_27_47# VPB 0.139f
C11 X A 0.014f
C12 VPB A 0.0321f
C13 a_27_47# A 0.195f
C14 VGND VPWR 0.057f
C15 VGND VNB 0.358f
C16 X VNB 0.067f
C17 VPWR VNB 0.308f
C18 A VNB 0.148f
C19 VPB VNB 0.605f
C20 a_27_47# VNB 0.543f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
C0 A VPWR 0.0362f
C1 A B 0.0971f
C2 a_59_75# VPWR 0.15f
C3 a_59_75# B 0.143f
C4 A a_59_75# 0.0809f
C5 X VPWR 0.111f
C6 B X 0.00276f
C7 VPB VPWR 0.0729f
C8 B VPB 0.0629f
C9 A X 1.68e-19
C10 A VPB 0.0806f
C11 VGND VPWR 0.0461f
C12 VGND B 0.0115f
C13 a_145_75# VPWR 6.31e-19
C14 a_59_75# X 0.109f
C15 VGND A 0.0147f
C16 a_59_75# VPB 0.0563f
C17 VPB X 0.0127f
C18 VGND a_59_75# 0.116f
C19 a_145_75# a_59_75# 0.00658f
C20 VGND X 0.0993f
C21 a_145_75# X 5.76e-19
C22 VGND VPB 0.008f
C23 B VPWR 0.0117f
C24 VGND a_145_75# 0.00468f
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y a_297_297# a_191_297#
+ a_109_297#
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPWR B 0.0887f
C1 A B 0.11f
C2 VPWR D 0.0128f
C3 B C 0.173f
C4 B VPB 0.0304f
C5 B VGND 0.0191f
C6 A VPWR 0.0483f
C7 D C 0.0523f
C8 VPB D 0.0376f
C9 VPWR a_109_297# 0.00576f
C10 B a_297_297# 0.0132f
C11 VPWR C 0.0509f
C12 a_191_297# B 0.00223f
C13 Y B 0.0403f
C14 VGND D 0.0456f
C15 VPWR VPB 0.0524f
C16 A C 0.00268f
C17 VPWR VGND 0.0492f
C18 A VPB 0.041f
C19 A VGND 0.0526f
C20 Y D 0.108f
C21 a_109_297# C 0.0062f
C22 VPWR a_297_297# 0.00317f
C23 a_191_297# VPWR 0.0049f
C24 Y VPWR 0.0561f
C25 VPB C 0.0299f
C26 VGND a_109_297# 0.00181f
C27 VGND C 0.0184f
C28 A a_297_297# 3.16e-19
C29 Y A 0.0175f
C30 VGND VPB 0.0048f
C31 a_191_297# C 0.0195f
C32 Y a_109_297# 0.0122f
C33 Y C 0.125f
C34 Y VPB 0.0127f
C35 VGND a_297_297# 8.1e-19
C36 a_191_297# VGND 9.29e-19
C37 Y VGND 0.151f
C38 Y a_297_297# 1.24e-19
C39 a_191_297# Y 0.00142f
C40 VGND VNB 0.322f
C41 VPWR VNB 0.276f
C42 Y VNB 0.0645f
C43 A VNB 0.174f
C44 B VNB 0.0968f
C45 C VNB 0.0911f
C46 D VNB 0.159f
C47 VPB VNB 0.516f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X a_75_212#
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 VGND VPWR 0.0289f
C1 VGND a_75_212# 0.105f
C2 A VPWR 0.0217f
C3 A a_75_212# 0.178f
C4 VGND A 0.0184f
C5 X VPWR 0.0896f
C6 a_75_212# X 0.107f
C7 VGND X 0.0545f
C8 VPB VPWR 0.0355f
C9 VPB a_75_212# 0.0571f
C10 A X 8.48e-19
C11 VPB VGND 0.00507f
C12 VPB A 0.0525f
C13 VPB X 0.0128f
C14 a_75_212# VPWR 0.134f
C15 VGND VNB 0.207f
C16 VPWR VNB 0.176f
C17 X VNB 0.0942f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_75_212# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 VGND X 0.0546f
C1 VGND a_27_47# 0.105f
C2 A X 8.48e-19
C3 A a_27_47# 0.181f
C4 VGND A 0.0184f
C5 VPWR X 0.0897f
C6 a_27_47# VPWR 0.135f
C7 VGND VPWR 0.029f
C8 VPB X 0.0128f
C9 VPB a_27_47# 0.0592f
C10 A VPWR 0.0215f
C11 VPB VGND 0.00505f
C12 VPB A 0.0524f
C13 VPB VPWR 0.0355f
C14 a_27_47# X 0.107f
C15 VGND VNB 0.207f
C16 X VNB 0.0941f
C17 VPWR VNB 0.175f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_27_47# VNB 0.208f
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X a_664_47# a_841_47#
+ a_381_47# a_62_47# a_558_47#
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPB a_62_47# 0.0515f
C1 VPB a_664_47# 0.043f
C2 VPB a_381_47# 0.0447f
C3 a_62_47# X 0.156f
C4 a_62_47# A 0.244f
C5 VPB X 0.126f
C6 VPB A 0.105f
C7 VPB a_841_47# 0.0108f
C8 a_664_47# X 6.67e-19
C9 a_62_47# VGND 0.144f
C10 VPWR a_62_47# 0.149f
C11 a_381_47# X 0.318f
C12 a_381_47# A 5.42e-19
C13 a_664_47# a_841_47# 0.134f
C14 VPB VGND 0.008f
C15 VPWR VPB 0.103f
C16 a_558_47# VPB 0.115f
C17 X A 0.0142f
C18 a_664_47# VGND 0.125f
C19 VPWR a_664_47# 0.131f
C20 a_558_47# a_664_47# 0.314f
C21 a_381_47# VGND 0.125f
C22 VPWR a_381_47# 0.134f
C23 a_558_47# a_381_47# 0.16f
C24 VGND X 0.106f
C25 VGND A 0.0176f
C26 VPWR X 0.108f
C27 VPWR A 0.0174f
C28 a_558_47# X 0.0144f
C29 a_841_47# VGND 0.0585f
C30 VPWR a_841_47# 0.0614f
C31 a_558_47# a_841_47# 0.00368f
C32 VPWR VGND 0.0902f
C33 a_558_47# VGND 0.0816f
C34 VPWR a_558_47# 0.084f
C35 VGND VNB 0.537f
C36 VPWR VNB 0.439f
C37 X VNB 0.163f
C38 A VNB 0.198f
C39 VPB VNB 0.959f
C40 a_841_47# VNB 0.0929f
C41 a_664_47# VNB 0.13f
C42 a_558_47# VNB 0.164f
C43 a_381_47# VNB 0.11f
C44 a_62_47# VNB 0.169f
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y a_129_47# a_47_47# a_285_47#
+ a_377_297#
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 A VPWR 0.0349f
C1 VPWR B 0.0408f
C2 A B 0.236f
C3 Y VPWR 0.107f
C4 A Y 0.00181f
C5 VPWR a_377_297# 0.00559f
C6 VPWR a_47_47# 0.273f
C7 Y B 0.00334f
C8 VPWR VPB 0.0718f
C9 A a_47_47# 0.0307f
C10 A VPB 0.0822f
C11 a_377_297# B 0.00254f
C12 B a_47_47# 0.356f
C13 VPB B 0.0643f
C14 VPWR a_285_47# 0.00255f
C15 a_129_47# VPWR 9.47e-19
C16 VGND VPWR 0.0665f
C17 Y a_377_297# 0.00188f
C18 Y a_47_47# 0.143f
C19 A a_285_47# 0.0353f
C20 VGND A 0.0635f
C21 Y VPB 0.00878f
C22 a_285_47# B 0.067f
C23 a_129_47# B 0.00236f
C24 VGND B 0.0389f
C25 a_377_297# a_47_47# 0.00899f
C26 VPB a_47_47# 0.0444f
C27 Y a_285_47# 0.0439f
C28 VGND Y 0.0381f
C29 a_285_47# a_47_47# 0.0175f
C30 a_129_47# a_47_47# 0.00369f
C31 VGND a_377_297# 0.00125f
C32 VGND a_47_47# 0.104f
C33 a_285_47# VPB 5.53e-19
C34 VGND VPB 0.00568f
C35 VGND a_285_47# 0.211f
C36 a_129_47# VGND 0.00547f
C37 VGND VNB 0.4f
C38 Y VNB 0.0783f
C39 VPWR VNB 0.352f
C40 A VNB 0.217f
C41 B VNB 0.212f
C42 VPB VNB 0.693f
C43 a_285_47# VNB 0.0174f
C44 a_47_47# VNB 0.199f
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X a_472_297# a_80_21#
+ a_300_47# a_217_297#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
C0 VGND A1 0.0147f
C1 a_80_21# A2 0.128f
C2 a_80_21# a_217_297# 0.127f
C3 A1 A2 0.0881f
C4 a_217_297# A1 0.0124f
C5 VGND a_472_297# 0.00188f
C6 a_80_21# A1 0.111f
C7 a_472_297# a_217_297# 0.00517f
C8 VGND C1 0.0176f
C9 VGND B1 0.0175f
C10 a_80_21# a_472_297# 0.0164f
C11 VGND VPB 0.00775f
C12 a_217_297# C1 0.00262f
C13 a_217_297# B1 0.00651f
C14 VPB A2 0.0384f
C15 a_217_297# VPB 0.00494f
C16 a_80_21# C1 0.079f
C17 a_80_21# B1 0.0964f
C18 VGND VPWR 0.0665f
C19 X VGND 0.0654f
C20 a_300_47# VGND 0.00536f
C21 A1 B1 0.0834f
C22 a_80_21# VPB 0.0661f
C23 VPWR A2 0.0161f
C24 a_217_297# VPWR 0.197f
C25 X A2 6.82e-19
C26 X a_217_297# 0.00271f
C27 VPB A1 0.0266f
C28 a_472_297# B1 1.87e-19
C29 a_80_21# VPWR 0.119f
C30 X a_80_21# 0.118f
C31 a_300_47# a_80_21# 0.00997f
C32 VPWR A1 0.0149f
C33 X A1 3.62e-19
C34 a_300_47# A1 5.95e-19
C35 C1 B1 0.0846f
C36 VPB C1 0.0379f
C37 VPB B1 0.0267f
C38 a_472_297# VPWR 0.00703f
C39 X a_472_297# 2.6e-19
C40 VPWR C1 0.0137f
C41 VPWR B1 0.0129f
C42 X C1 7.15e-20
C43 X B1 1.18e-19
C44 VPB VPWR 0.0754f
C45 X VPB 0.0118f
C46 VGND A2 0.0191f
C47 VGND a_217_297# 0.00342f
C48 a_80_21# VGND 0.293f
C49 X VPWR 0.0884f
C50 a_217_297# A2 0.0135f
C51 a_300_47# VPWR 8.53e-19
C52 X a_300_47# 5.31e-19
C53 VGND VNB 0.385f
C54 VPWR VNB 0.325f
C55 X VNB 0.0899f
C56 C1 VNB 0.144f
C57 B1 VNB 0.0899f
C58 A1 VNB 0.0905f
C59 A2 VNB 0.108f
C60 VPB VNB 0.693f
C61 a_217_297# VNB 0.00117f
C62 a_80_21# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPB a_27_47# 0.082f
C1 C B 0.161f
C2 C D 0.18f
C3 VPB VGND 0.00852f
C4 a_27_47# B 0.13f
C5 D a_27_47# 0.107f
C6 VPB VPWR 0.077f
C7 VGND B 0.0453f
C8 VGND D 0.0898f
C9 C a_27_47# 0.0516f
C10 VPWR B 0.0231f
C11 VPWR D 0.0207f
C12 C VGND 0.0408f
C13 VPB A 0.0907f
C14 C VPWR 0.021f
C15 VGND a_27_47# 0.132f
C16 a_197_47# B 0.00623f
C17 B a_109_47# 0.00153f
C18 VPWR a_27_47# 0.326f
C19 A B 0.0839f
C20 C a_197_47# 0.00123f
C21 C a_109_47# 1.72e-20
C22 VPWR VGND 0.0662f
C23 X VPB 0.0111f
C24 a_197_47# a_27_47# 0.00167f
C25 a_27_47# a_109_47# 0.00578f
C26 A a_27_47# 0.153f
C27 VGND a_197_47# 0.00387f
C28 VGND a_109_47# 0.00223f
C29 a_303_47# D 0.00119f
C30 X D 0.00746f
C31 VPWR a_197_47# 5.24e-19
C32 VGND A 0.0151f
C33 VPWR a_109_47# 4.66e-19
C34 a_303_47# C 0.00527f
C35 VPWR A 0.044f
C36 a_303_47# a_27_47# 0.00119f
C37 X a_27_47# 0.0754f
C38 a_303_47# VGND 0.00381f
C39 X VGND 0.0903f
C40 a_303_47# VPWR 4.83e-19
C41 X VPWR 0.0945f
C42 VPB B 0.0643f
C43 VPB D 0.0782f
C44 C VPB 0.0609f
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X a_489_413# a_226_47#
+ a_556_47# a_226_297# a_76_199#
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VGND B1 0.0471f
C1 a_226_47# a_76_199# 0.188f
C2 a_226_47# a_489_413# 0.00579f
C3 B1 a_76_199# 0.00185f
C4 a_489_413# B1 0.0382f
C5 VGND a_226_297# 5.63e-19
C6 a_226_297# a_76_199# 0.00354f
C7 VGND VPWR 0.0743f
C8 VGND X 0.0627f
C9 VGND B2 0.0335f
C10 a_226_47# a_226_297# 0.00128f
C11 VGND VPB 0.0128f
C12 VPWR a_76_199# 0.2f
C13 a_489_413# VPWR 0.143f
C14 a_76_199# X 0.0995f
C15 B2 a_76_199# 0.0626f
C16 a_489_413# B2 0.0541f
C17 VPB a_76_199# 0.0817f
C18 a_489_413# VPB 0.015f
C19 a_226_47# VPWR 0.0187f
C20 a_226_47# X 0.0108f
C21 VGND A2_N 0.0174f
C22 A1_N VGND 0.0261f
C23 a_556_47# VGND 0.00639f
C24 a_226_47# B2 0.0975f
C25 VPWR B1 0.0188f
C26 a_226_47# VPB 0.111f
C27 B2 B1 0.182f
C28 A2_N a_76_199# 0.0125f
C29 A1_N a_76_199# 0.119f
C30 a_556_47# a_76_199# 0.0017f
C31 VPB B1 0.0803f
C32 a_226_297# VPWR 8.54e-19
C33 a_226_47# A2_N 0.141f
C34 A1_N a_226_47# 0.0209f
C35 VPWR X 0.0589f
C36 B2 VPWR 0.0161f
C37 VPB VPWR 0.0951f
C38 VPB X 0.0113f
C39 A1_N a_226_297# 0.00184f
C40 VPB B2 0.0645f
C41 A2_N VPWR 0.00449f
C42 A2_N X 2.55e-19
C43 A1_N VPWR 0.00672f
C44 A1_N X 0.00211f
C45 a_556_47# VPWR 7.24e-19
C46 a_556_47# B2 0.00291f
C47 VPB A2_N 0.0327f
C48 A1_N VPB 0.0339f
C49 VGND a_76_199# 0.108f
C50 VGND a_489_413# 0.0058f
C51 a_226_47# VGND 0.149f
C52 A1_N A2_N 0.11f
C53 a_489_413# a_76_199# 0.0473f
C54 VGND VNB 0.462f
C55 A2_N VNB 0.103f
C56 A1_N VNB 0.111f
C57 VPWR VNB 0.369f
C58 X VNB 0.0975f
C59 B1 VNB 0.206f
C60 B2 VNB 0.106f
C61 VPB VNB 0.782f
C62 a_489_413# VNB 0.0254f
C63 a_226_47# VNB 0.162f
C64 a_76_199# VNB 0.141f
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X a_515_93# a_223_47#
+ a_615_93# a_343_93# a_429_93# a_27_47#
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
C0 VGND A_N 0.0146f
C1 VGND C 0.025f
C2 B_N A_N 0.117f
C3 B_N C 9.56e-20
C4 VGND B_N 0.0427f
C5 a_223_47# A_N 0.00833f
C6 C a_223_47# 0.151f
C7 VGND a_223_47# 0.199f
C8 B_N a_223_47# 0.0431f
C9 D C 0.163f
C10 VGND X 0.0609f
C11 B_N X 4.64e-20
C12 VGND D 0.0414f
C13 B_N D 6.67e-20
C14 C a_343_93# 0.0397f
C15 D a_223_47# 4.03e-19
C16 a_27_47# A_N 0.0906f
C17 VGND a_429_93# 0.00122f
C18 VGND a_343_93# 0.0548f
C19 VPB A_N 0.0848f
C20 C VPB 0.0686f
C21 B_N a_343_93# 0.00112f
C22 D X 0.0193f
C23 VGND a_27_47# 0.0715f
C24 B_N a_27_47# 0.138f
C25 VGND VPB 0.0167f
C26 a_429_93# a_223_47# 0.00492f
C27 a_223_47# a_343_93# 0.269f
C28 B_N VPB 0.0646f
C29 a_27_47# a_223_47# 0.267f
C30 C a_615_93# 0.00407f
C31 X a_343_93# 0.126f
C32 a_515_93# C 0.00389f
C33 VPWR A_N 0.0318f
C34 VPB a_223_47# 0.0799f
C35 VPWR C 0.012f
C36 D a_343_93# 0.114f
C37 VGND a_615_93# 0.0044f
C38 a_515_93# VGND 0.00408f
C39 X VPB 0.0103f
C40 VGND VPWR 0.0906f
C41 VPWR B_N 0.0168f
C42 D VPB 0.081f
C43 a_515_93# a_223_47# 0.00482f
C44 VPWR a_223_47# 0.114f
C45 a_429_93# a_343_93# 0.00484f
C46 VPWR X 0.0582f
C47 a_27_47# a_343_93# 0.0406f
C48 VPB a_343_93# 0.0857f
C49 D a_615_93# 0.00564f
C50 VPWR D 0.0143f
C51 VPB a_27_47# 0.154f
C52 a_615_93# a_343_93# 0.00103f
C53 a_515_93# a_343_93# 0.00115f
C54 VPWR a_429_93# 5.19e-19
C55 VPWR a_343_93# 0.255f
C56 VPWR a_27_47# 0.0897f
C57 VPWR VPB 0.106f
C58 VPWR a_615_93# 8.49e-19
C59 a_515_93# VPWR 7.86e-19
C60 VGND VNB 0.553f
C61 X VNB 0.0908f
C62 VPWR VNB 0.453f
C63 D VNB 0.124f
C64 C VNB 0.107f
C65 B_N VNB 0.134f
C66 A_N VNB 0.144f
C67 VPB VNB 0.959f
C68 a_343_93# VNB 0.172f
C69 a_223_47# VNB 0.141f
C70 a_27_47# VNB 0.259f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 B a_35_297# 0.203f
C1 B a_285_297# 0.0553f
C2 a_117_297# a_35_297# 0.00641f
C3 B a_117_297# 0.00777f
C4 X a_35_297# 0.166f
C5 a_285_297# X 0.0712f
C6 VPB a_35_297# 0.0699f
C7 VPB a_285_297# 0.0133f
C8 B X 0.0149f
C9 a_117_297# X 2.25e-19
C10 a_285_47# a_35_297# 0.00723f
C11 B VPB 0.0697f
C12 B a_285_47# 3.98e-19
C13 VPB X 0.0154f
C14 a_35_297# VGND 0.177f
C15 a_285_297# VGND 0.00394f
C16 a_285_47# X 0.00206f
C17 VPWR a_35_297# 0.096f
C18 a_285_297# VPWR 0.246f
C19 B VGND 0.0304f
C20 A a_35_297# 0.0633f
C21 a_285_297# A 0.00749f
C22 a_117_297# VGND 0.00177f
C23 B VPWR 0.0703f
C24 a_117_297# VPWR 0.00852f
C25 B A 0.221f
C26 X VGND 0.173f
C27 VPWR X 0.0537f
C28 VPB VGND 0.00696f
C29 A X 0.00166f
C30 VPB VPWR 0.0689f
C31 a_285_47# VGND 0.00552f
C32 VPB A 0.051f
C33 a_285_47# VPWR 8.6e-19
C34 VPWR VGND 0.0643f
C35 A VGND 0.0325f
C36 A VPWR 0.0348f
C37 a_285_297# a_35_297# 0.025f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X a_465_297# a_297_297#
+ a_215_297# a_392_297# a_109_53#
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 VPB a_109_53# 0.0547f
C1 VPB VGND 0.0115f
C2 a_109_53# B 0.0246f
C3 C a_109_53# 0.0984f
C4 VPB A 0.0325f
C5 VGND B 0.0161f
C6 VGND C 0.0202f
C7 D_N a_109_53# 0.0889f
C8 A B 0.0666f
C9 A C 0.0281f
C10 D_N VGND 0.0531f
C11 VPB a_215_297# 0.0508f
C12 VPB VPWR 0.122f
C13 VGND a_109_53# 0.118f
C14 C a_392_297# 0.00267f
C15 C a_297_297# 0.00375f
C16 A a_109_53# 1.19e-19
C17 a_215_297# B 0.159f
C18 C a_215_297# 0.161f
C19 VPWR B 0.255f
C20 C VPWR 0.00753f
C21 A VGND 0.0158f
C22 X VPB 0.011f
C23 D_N a_215_297# 3.19e-19
C24 a_109_53# a_297_297# 7.06e-21
C25 D_N VPWR 0.0412f
C26 a_215_297# a_109_53# 0.0807f
C27 VGND a_392_297# 3.44e-19
C28 VGND a_297_297# 6.5e-19
C29 a_465_297# C 6.89e-19
C30 X B 6.65e-19
C31 VPWR a_109_53# 0.0418f
C32 VGND a_215_297# 0.237f
C33 VGND VPWR 0.075f
C34 A a_215_297# 0.157f
C35 A VPWR 0.0073f
C36 a_465_297# VGND 5.02e-19
C37 X VGND 0.0359f
C38 a_215_297# a_392_297# 0.00419f
C39 a_215_297# a_297_297# 0.00659f
C40 VPWR a_392_297# 5.29e-19
C41 VPWR a_297_297# 8.59e-19
C42 a_465_297# A 5.42e-19
C43 X A 0.00127f
C44 VPWR a_215_297# 0.0871f
C45 a_465_297# a_215_297# 0.00827f
C46 X a_215_297# 0.0991f
C47 a_465_297# VPWR 7.08e-19
C48 X VPWR 0.0885f
C49 VPB B 0.116f
C50 VPB C 0.0337f
C51 D_N VPB 0.0461f
C52 C B 0.0893f
C53 VGND VNB 0.469f
C54 X VNB 0.0884f
C55 A VNB 0.108f
C56 C VNB 0.101f
C57 D_N VNB 0.185f
C58 B VNB 0.101f
C59 VPWR VNB 0.399f
C60 VPB VNB 0.782f
C61 a_109_53# VNB 0.159f
C62 a_215_297# VNB 0.142f
.ends

.subckt therm VGND VPWR b[0] b[1] b[2] b[3] p[0] p[10] p[11] p[12] p[13] p[14] p[1]
+ p[2] p[3] p[4] p[5] p[6] p[7] p[8] p[9]
X_49_ net7 _02_ _19_ _20_ _21_ VGND VGND VPWR VPWR net17 _49_/a_208_47# _49_/a_75_199#
+ _49_/a_544_297# _49_/a_315_47# _49_/a_201_297# sky130_fd_sc_hd__a311o_1
X_48_ net11 _02_ _07_ VGND VGND VPWR VPWR _21_ _48_/a_181_47# _48_/a_109_47# _48_/a_27_47#
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ net5 _12_ _17_ VGND VGND VPWR VPWR _20_ _47_/a_384_47# _47_/a_81_21# _47_/a_299_297#
+ sky130_fd_sc_hd__a21o_1
X_46_ _04_ VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__inv_2
X_29_ net11 net13 net12 VGND VGND VPWR VPWR _03_ _29_/a_29_53# _29_/a_183_297# _29_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_28_ _00_ _01_ VGND VGND VPWR VPWR _02_ _28_/a_109_297# sky130_fd_sc_hd__nor2_1
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_45_ _02_ _09_ _12_ _13_ _18_ VGND VGND VPWR VPWR net16 _45_/a_193_297# _45_/a_465_47#
+ _45_/a_205_47# _45_/a_109_297# _45_/a_27_47# sky130_fd_sc_hd__a221o_1
X_44_ net14 _14_ _15_ _17_ net2 VGND VGND VPWR VPWR _18_ _44_/a_256_47# _44_/a_584_47#
+ _44_/a_93_21# _44_/a_250_297# _44_/a_346_47# sky130_fd_sc_hd__a32o_1
X_27_ net14 net15 net3 net2 VGND VGND VPWR VPWR _01_ _27_/a_277_297# _27_/a_205_297#
+ _27_/a_27_297# _27_/a_109_297# sky130_fd_sc_hd__or4_1
XFILLER_0_7_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_26_ net5 net4 net6 VGND VGND VPWR VPWR _00_ _26_/a_29_53# _26_/a_183_297# _26_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_43_ _00_ _06_ _10_ _16_ VGND VGND VPWR VPWR _17_ _43_/a_369_47# _43_/a_469_47# _43_/a_297_47#
+ _43_/a_193_413# _43_/a_27_47# sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_42_ net3 net15 net14 VGND VGND VPWR VPWR _16_ _42_/a_109_93# _42_/a_368_53# _42_/a_209_311#
+ _42_/a_296_53# sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_3_Left_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND VPWR VPWR b[0] output16/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_41_ _06_ _10_ VGND VGND VPWR VPWR _15_ _41_/a_145_75# _41_/a_59_75# sky130_fd_sc_hd__and2_1
Xoutput17 net17 VGND VGND VPWR VPWR b[1] output17/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_40_ net15 net3 net2 _00_ VGND VGND VPWR VPWR _14_ _40_/a_297_297# _40_/a_191_297#
+ _40_/a_109_297# sky130_fd_sc_hd__nor4_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput18 net18 VGND VGND VPWR VPWR b[2] output18/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_0_Left_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR b[3] output19/a_27_47# sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 p[0] VGND VGND VPWR VPWR net1 input1/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput2 p[10] VGND VGND VPWR VPWR net2 input2/a_27_47# sky130_fd_sc_hd__buf_1
Xinput3 p[11] VGND VGND VPWR VPWR net3 input3/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 p[12] VGND VGND VPWR VPWR net4 input4/a_75_212# sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 p[13] VGND VGND VPWR VPWR net5 input5/a_664_47# input5/a_841_47# input5/a_381_47#
+ input5/a_62_47# input5/a_558_47# sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_1_Left_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 p[14] VGND VGND VPWR VPWR net6 input6/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 p[1] VGND VGND VPWR VPWR net7 input7/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput10 p[4] VGND VGND VPWR VPWR net10 input10/a_27_47# sky130_fd_sc_hd__buf_1
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 p[2] VGND VGND VPWR VPWR net8 input8/a_27_47# sky130_fd_sc_hd__buf_1
Xinput11 p[5] VGND VGND VPWR VPWR net11 input11/a_27_47# sky130_fd_sc_hd__buf_1
X_39_ net5 net6 VGND VGND VPWR VPWR _13_ _39_/a_129_47# _39_/a_47_47# _39_/a_285_47#
+ _39_/a_377_297# sky130_fd_sc_hd__xnor2_1
Xinput9 p[3] VGND VGND VPWR VPWR net9 input9/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput12 p[6] VGND VGND VPWR VPWR net12 input12/a_27_47# sky130_fd_sc_hd__buf_1
X_55_ _14_ _15_ _20_ _22_ VGND VGND VPWR VPWR net19 _55_/a_472_297# _55_/a_80_21#
+ _55_/a_300_47# _55_/a_217_297# sky130_fd_sc_hd__a211o_1
X_38_ net4 _06_ _10_ _11_ VGND VGND VPWR VPWR _12_ _38_/a_109_47# _38_/a_197_47# _38_/a_303_47#
+ _38_/a_27_47# sky130_fd_sc_hd__and4_1
X_54_ _25_ VGND VGND VPWR VPWR net18 _54_/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput13 p[7] VGND VGND VPWR VPWR net13 input13/a_27_47# sky130_fd_sc_hd__buf_1
X_37_ net14 net15 net3 net2 VGND VGND VPWR VPWR _11_ _37_/a_109_47# _37_/a_197_47#
+ _37_/a_303_47# _37_/a_27_47# sky130_fd_sc_hd__and4_1
Xinput14 p[8] VGND VGND VPWR VPWR net14 input14/a_27_47# sky130_fd_sc_hd__buf_1
X_53_ _21_ _22_ _24_ VGND VGND VPWR VPWR _25_ _53_/a_29_53# _53_/a_183_297# _53_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_36_ net11 net10 net13 net12 VGND VGND VPWR VPWR _10_ _36_/a_109_47# _36_/a_197_47#
+ _36_/a_303_47# _36_/a_27_47# sky130_fd_sc_hd__and4_1
X_52_ _02_ _06_ _23_ _12_ net5 VGND VGND VPWR VPWR _24_ _52_/a_256_47# _52_/a_584_47#
+ _52_/a_93_21# _52_/a_250_297# _52_/a_346_47# sky130_fd_sc_hd__a32o_1
Xinput15 p[9] VGND VGND VPWR VPWR net15 input15/a_27_47# sky130_fd_sc_hd__buf_1
X_35_ _04_ _05_ _07_ _08_ VGND VGND VPWR VPWR _09_ _35_/a_489_413# _35_/a_226_47#
+ _35_/a_556_47# _35_/a_226_297# _35_/a_76_199# sky130_fd_sc_hd__a2bb2o_1
X_51_ _03_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__inv_2
X_34_ net11 net12 VGND VGND VPWR VPWR _08_ _34_/a_129_47# _34_/a_47_47# _34_/a_285_47#
+ _34_/a_377_297# sky130_fd_sc_hd__xnor2_1
X_33_ net13 _06_ net10 VGND VGND VPWR VPWR _07_ _33_/a_109_93# _33_/a_368_53# _33_/a_209_311#
+ _33_/a_296_53# sky130_fd_sc_hd__and3b_1
X_50_ net5 net6 _15_ _11_ VGND VGND VPWR VPWR _22_ _50_/a_515_93# _50_/a_223_47# _50_/a_615_93#
+ _50_/a_343_93# _50_/a_429_93# _50_/a_27_47# sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ net7 net1 net9 net8 VGND VGND VPWR VPWR _06_ _32_/a_109_47# _32_/a_197_47# _32_/a_303_47#
+ _32_/a_27_47# sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_5_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31_ net7 net8 VGND VGND VPWR VPWR _05_ _31_/a_117_297# _31_/a_285_297# _31_/a_285_47#
+ _31_/a_35_297# sky130_fd_sc_hd__xor2_1
X_30_ net9 net10 _03_ net1 VGND VGND VPWR VPWR _04_ _30_/a_465_297# _30_/a_297_297#
+ _30_/a_215_297# _30_/a_392_297# _30_/a_109_53# sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
C0 net8 _22_ 3.3e-20
C1 net13 _13_ 4e-21
C2 net6 b[3] 7.68e-19
C3 input5/a_664_47# p[1] 1.21e-20
C4 _00_ _50_/a_223_47# 0.00738f
C5 _10_ _53_/a_29_53# 0.00779f
C6 net6 _40_/a_191_297# 1.16e-20
C7 net3 _17_ 0.0698f
C8 _04_ input3/a_27_47# 3.55e-19
C9 _01_ p[13] 2.02e-20
C10 _20_ VPWR 0.342f
C11 VPWR _30_/a_297_297# -4.57e-19
C12 _42_/a_109_93# output17/a_27_47# 8.6e-21
C13 _15_ _55_/a_300_47# 1.42e-20
C14 _43_/a_369_47# _43_/a_193_413# -1.25e-19
C15 VPWR _09_ 0.297f
C16 p[9] VPWR 0.374f
C17 _30_/a_109_53# net9 0.0193f
C18 _02_ _01_ 0.106f
C19 _03_ _08_ 0.0144f
C20 input13/a_27_47# input9/a_75_212# 0.00732f
C21 _02_ _34_/a_47_47# 1.09e-19
C22 _19_ net7 0.0458f
C23 _15_ _50_/a_615_93# 0.00183f
C24 _35_/a_76_199# _33_/a_209_311# 9.95e-21
C25 _06_ _52_/a_584_47# 0.00218f
C26 net5 _52_/a_584_47# 0.0022f
C27 input2/a_27_47# net7 0.00213f
C28 _20_ _39_/a_129_47# 1.71e-20
C29 VPWR _19_ 0.0335f
C30 _02_ _30_/a_109_53# 5.03e-22
C31 _21_ input9/a_75_212# 1.17e-21
C32 _01_ net3 1.16e-19
C33 _35_/a_226_47# p[7] 2.82e-19
C34 net11 _04_ 0.078f
C35 net12 _36_/a_197_47# 4.67e-20
C36 _15_ _43_/a_193_413# 4.86e-19
C37 _01_ _17_ 1.46e-20
C38 _01_ _49_/a_201_297# 0.0105f
C39 input3/a_27_47# output17/a_27_47# 3.15e-19
C40 input14/a_27_47# _44_/a_250_297# 8.25e-21
C41 VPWR input2/a_27_47# 0.00872f
C42 net3 _27_/a_109_297# 5.45e-19
C43 net14 p[14] 6.11e-20
C44 _35_/a_226_47# _04_ 0.00551f
C45 b[3] _22_ 1.28e-19
C46 net14 _11_ 5e-19
C47 _15_ net2 9.8e-19
C48 _06_ _50_/a_515_93# 0.00244f
C49 net12 input10/a_27_47# 0.00115f
C50 _09_ _35_/a_226_297# 4.98e-19
C51 _55_/a_80_21# _43_/a_27_47# 1.56e-19
C52 _21_ _13_ 1.69e-19
C53 _20_ _28_/a_109_297# 0.00221f
C54 _45_/a_109_297# net16 5.1e-20
C55 _45_/a_27_47# _00_ 4.84e-20
C56 _47_/a_81_21# net2 4.95e-19
C57 input5/a_664_47# net8 0.0116f
C58 _06_ _43_/a_27_47# 0.0329f
C59 _44_/a_93_21# p[14] 2.82e-20
C60 _03_ net9 0.15f
C61 _44_/a_93_21# _11_ 4.78e-20
C62 net6 p[14] 0.00237f
C63 VPWR _34_/a_129_47# -9.47e-19
C64 _35_/a_489_413# _07_ 0.00429f
C65 _10_ _50_/a_515_93# 0.00129f
C66 input14/a_27_47# net19 1.44e-19
C67 net6 _11_ 0.0257f
C68 net11 b[2] 1.46e-19
C69 _44_/a_346_47# net2 1.64e-19
C70 net10 _36_/a_27_47# 0.0366f
C71 p[12] _15_ 0.0162f
C72 _14_ net17 2.4e-20
C73 _20_ net12 0.00437f
C74 b[2] _23_ 2.87e-20
C75 net12 _30_/a_297_297# 7.14e-21
C76 net12 _09_ 0.0374f
C77 _10_ _43_/a_27_47# 0.0279f
C78 _14_ _00_ 0.133f
C79 _35_/a_76_199# _11_ 6.99e-22
C80 _00_ _26_/a_29_53# 0.0466f
C81 VPWR _52_/a_346_47# -0.00109f
C82 _08_ net10 0.189f
C83 _13_ _52_/a_250_297# 5.43e-19
C84 _03_ _02_ 0.00474f
C85 _12_ _33_/a_209_311# 2.88e-20
C86 _55_/a_80_21# net8 1.84e-21
C87 _21_ _50_/a_223_47# 2.91e-21
C88 _13_ _53_/a_29_53# 9.05e-19
C89 net14 _50_/a_615_93# 1.69e-20
C90 _42_/a_209_311# _18_ 3.21e-19
C91 p[10] _05_ 6e-20
C92 _06_ net8 0.00282f
C93 _15_ _55_/a_217_297# 0.0474f
C94 _20_ _27_/a_27_297# 3.14e-20
C95 net5 net8 0.48f
C96 input4/a_75_212# input15/a_27_47# 1.1e-21
C97 net14 _43_/a_193_413# 1.11e-19
C98 input5/a_381_47# net17 1.37e-20
C99 _03_ net3 4.27e-20
C100 _31_/a_285_47# _05_ 5.61e-19
C101 net17 net7 0.2f
C102 _32_/a_27_47# _05_ 2.2e-20
C103 _03_ _49_/a_201_297# 0.00842f
C104 _10_ net8 5.86e-19
C105 net13 _26_/a_29_53# 2.23e-20
C106 net6 _50_/a_615_93# 1.43e-19
C107 _11_ _22_ 0.15f
C108 net14 net2 0.151f
C109 input8/a_27_47# _04_ 2.36e-22
C110 _00_ net7 8.12e-21
C111 _04_ _07_ 9.74e-20
C112 _43_/a_469_47# _17_ 0.00177f
C113 p[5] p[4] 0.385f
C114 _31_/a_117_297# net17 0.00149f
C115 _04_ _05_ 0.0352f
C116 p[9] net15 0.00306f
C117 _20_ net15 0.0021f
C118 _44_/a_93_21# _43_/a_193_413# 0.0161f
C119 VPWR net17 0.0371f
C120 _27_/a_27_297# _19_ 0.082f
C121 _29_/a_183_297# net9 3.51e-19
C122 net2 net1 1.64e-19
C123 net6 _43_/a_193_413# 2.41e-20
C124 net14 p[8] 0.00868f
C125 net10 net9 0.111f
C126 VPWR _00_ 0.416f
C127 input5/a_62_47# net8 2.05e-19
C128 _30_/a_215_297# _29_/a_29_53# 1.72e-19
C129 _21_ _24_ 0.0388f
C130 input2/a_27_47# _27_/a_27_297# 1.16e-19
C131 _26_/a_111_297# _00_ 3.7e-19
C132 _44_/a_93_21# net2 0.0273f
C133 input12/a_27_47# net1 7.44e-20
C134 net6 net2 0.00139f
C135 p[4] net10 0.00268f
C136 _55_/a_80_21# b[3] 3.55e-19
C137 _11_ _50_/a_27_47# 0.0592f
C138 _03_ _01_ 2.85e-19
C139 _20_ _50_/a_343_93# 0.00826f
C140 _12_ _11_ 0.195f
C141 b[3] _06_ 9.96e-21
C142 input1/a_75_212# output17/a_27_47# 0.0101f
C143 net15 _19_ 0.00628f
C144 _31_/a_35_297# net8 0.0408f
C145 _55_/a_300_47# _22_ 2.08e-19
C146 _45_/a_27_47# _21_ 1.18e-20
C147 net6 p[8] 5.98e-19
C148 _03_ _34_/a_47_47# 4.5e-20
C149 net13 net7 1.72e-19
C150 _06_ _40_/a_191_297# 5.84e-19
C151 _39_/a_285_47# net16 1.29e-19
C152 input5/a_558_47# _42_/a_209_311# 7.85e-20
C153 _00_ _39_/a_129_47# 1.63e-20
C154 _02_ net10 3.52e-19
C155 _02_ net16 8.94e-19
C156 _03_ _27_/a_109_297# 1.97e-20
C157 _05_ output17/a_27_47# 1.12e-19
C158 input2/a_27_47# net15 1.61e-19
C159 _06_ _33_/a_209_311# 0.0187f
C160 output19/a_27_47# net14 0.00142f
C161 p[10] _42_/a_209_311# 2.37e-20
C162 _20_ _36_/a_27_47# 0.00148f
C163 _11_ _45_/a_193_297# 0.0292f
C164 _10_ b[3] 3.27e-20
C165 net13 VPWR 0.599f
C166 _52_/a_250_297# _24_ 3.03e-19
C167 _48_/a_109_47# _06_ 9.47e-19
C168 net6 p[12] 0.0941f
C169 net13 p[3] 9.49e-19
C170 _03_ _30_/a_109_53# 0.0189f
C171 net14 _55_/a_217_297# 2.1e-19
C172 _13_ _43_/a_27_47# 1.66e-20
C173 _53_/a_29_53# _24_ 0.0835f
C174 net3 _29_/a_183_297# 7.38e-21
C175 _27_/a_205_297# _04_ 6.42e-19
C176 _43_/a_193_413# _22_ 0.00133f
C177 _09_ _08_ 0.103f
C178 output19/a_27_47# _44_/a_93_21# 7.25e-20
C179 net11 _54_/a_75_212# 0.00956f
C180 input5/a_62_47# b[3] 0.00324f
C181 output19/a_27_47# net6 0.00112f
C182 p[0] input7/a_27_47# 5.13e-20
C183 p[0] p[13] 1.88e-19
C184 VPWR _36_/a_303_47# -4.83e-19
C185 _04_ _42_/a_209_311# 9.84e-22
C186 net2 _22_ 1.93e-20
C187 _21_ output18/a_27_47# 0.00103f
C188 _05_ _33_/a_368_53# 9.2e-19
C189 net12 net17 2.11e-21
C190 _06_ _52_/a_256_47# 0.00157f
C191 p[9] input6/a_27_47# 0.0762f
C192 p[9] input15/a_27_47# 0.0196f
C193 input13/a_27_47# p[3] 0.00101f
C194 input13/a_27_47# VPWR 0.0696f
C195 input14/a_27_47# p[11] 0.00118f
C196 _47_/a_299_297# _11_ 0.00738f
C197 _52_/a_93_21# net6 2.33e-19
C198 input13/a_27_47# p[6] 1.07e-19
C199 b[1] net1 1.78e-20
C200 _34_/a_285_47# _48_/a_27_47# 6.66e-20
C201 _12_ _43_/a_193_413# 7.94e-22
C202 _21_ net7 3e-19
C203 net13 _35_/a_226_297# 6.88e-19
C204 _10_ _52_/a_256_47# 1.65e-19
C205 p[12] _22_ 2.13e-21
C206 net8 net19 1.15e-19
C207 _15_ _42_/a_109_93# 0.00367f
C208 p[9] _37_/a_27_47# 0.0117f
C209 input10/a_27_47# p[4] 0.0215f
C210 _18_ _32_/a_27_47# 1.18e-20
C211 _06_ p[14] 1.04e-19
C212 _52_/a_93_21# _35_/a_76_199# 6.83e-21
C213 VPWR _33_/a_109_93# -0.00817f
C214 net4 _11_ 0.0858f
C215 _12_ net2 1.02e-20
C216 net6 _40_/a_297_297# 7.47e-22
C217 _11_ _06_ 0.493f
C218 _04_ _18_ 1.94e-21
C219 _27_/a_277_297# net8 7.99e-20
C220 _27_/a_27_297# net17 0.00181f
C221 _34_/a_47_47# net10 0.0507f
C222 _21_ VPWR 0.871f
C223 net5 _11_ 0.207f
C224 _21_ p[3] 3.95e-21
C225 _03_ _34_/a_377_297# 3.13e-20
C226 _21_ p[6] 0.00203f
C227 _20_ net9 0.328f
C228 output18/a_27_47# _53_/a_29_53# 9.46e-19
C229 _30_/a_297_297# net9 7.83e-19
C230 _09_ net9 2.62e-19
C231 input14/a_27_47# VPWR 0.0735f
C232 net11 _30_/a_215_297# 1.04e-19
C233 _10_ p[14] 1.53e-19
C234 net13 net12 0.363f
C235 _44_/a_250_297# b[3] 0.0112f
C236 _10_ _11_ 0.176f
C237 _30_/a_109_53# net10 5.6e-20
C238 _34_/a_129_47# _08_ 3.29e-19
C239 _16_ _15_ 0.0607f
C240 _12_ p[12] 2.08e-20
C241 p[12] _50_/a_27_47# 1.34e-19
C242 net15 net17 5.19e-19
C243 _09_ _45_/a_465_47# 2.77e-19
C244 input3/a_27_47# _15_ 7.53e-19
C245 _02_ _20_ 0.1f
C246 net15 _00_ 0.00147f
C247 _26_/a_29_53# _52_/a_584_47# 7.45e-20
C248 _02_ _09_ 0.297f
C249 _06_ _55_/a_300_47# 2.5e-20
C250 _52_/a_93_21# _22_ 0.0347f
C251 net14 _37_/a_109_47# 1.71e-19
C252 net14 _29_/a_29_53# 1.61e-20
C253 net12 _36_/a_303_47# 1.37e-19
C254 VPWR _52_/a_250_297# 0.019f
C255 input5/a_664_47# net2 8.11e-20
C256 p[10] input5/a_558_47# 1.09e-19
C257 _34_/a_285_47# _07_ 0.00975f
C258 _34_/a_285_47# _05_ 7.85e-21
C259 VPWR _53_/a_29_53# 0.00821f
C260 _54_/a_75_212# _38_/a_27_47# 2.67e-19
C261 b[3] net19 0.0439f
C262 _29_/a_29_53# net1 9.76e-19
C263 _06_ _50_/a_615_93# 0.00264f
C264 input7/a_27_47# _19_ 3.12e-21
C265 _20_ net3 4.07e-19
C266 input13/a_27_47# net12 0.0163f
C267 _09_ _35_/a_556_47# 3.74e-19
C268 _55_/a_80_21# _43_/a_193_413# 2.54e-19
C269 p[9] net3 1.63e-19
C270 _02_ _19_ 0.213f
C271 _45_/a_109_297# _00_ 4.86e-20
C272 _00_ _50_/a_343_93# 0.102f
C273 input2/a_27_47# input7/a_27_47# 1.62e-19
C274 _20_ _49_/a_201_297# 5.24e-21
C275 net6 _29_/a_29_53# 1.4e-20
C276 p[9] _17_ 1.03e-20
C277 _47_/a_299_297# net2 1.18e-19
C278 _20_ _17_ 0.102f
C279 _49_/a_201_297# _09_ 1.74e-20
C280 _06_ _43_/a_193_413# 0.0138f
C281 net11 _25_ 0.0262f
C282 input5/a_558_47# _04_ 1.25e-20
C283 net13 net15 8.84e-19
C284 _14_ _43_/a_27_47# 0.00938f
C285 _10_ _50_/a_615_93# 8.82e-19
C286 _52_/a_93_21# _12_ 0.0157f
C287 _25_ _23_ 0.00465f
C288 net5 _43_/a_193_413# 1.39e-20
C289 net14 _42_/a_109_93# 0.00351f
C290 _03_ _29_/a_183_297# 7.36e-19
C291 net12 _33_/a_109_93# 0.0435f
C292 p[10] _04_ 0.00306f
C293 _49_/a_75_199# _29_/a_29_53# 1.28e-19
C294 _35_/a_76_199# _29_/a_29_53# 9.88e-19
C295 _03_ net10 0.32f
C296 _21_ net12 0.23f
C297 _06_ net2 0.0108f
C298 _34_/a_377_297# net10 1.62e-19
C299 _10_ _43_/a_193_413# 0.0174f
C300 net5 net2 0.0616f
C301 _39_/a_47_47# _11_ 3.9e-19
C302 net3 _19_ 0.0129f
C303 VPWR _52_/a_584_47# -9.47e-19
C304 _52_/a_93_21# _45_/a_193_297# 6.01e-19
C305 p[1] net7 0.00514f
C306 input12/a_27_47# _06_ 5.3e-22
C307 _04_ p[7] 0.00142f
C308 _19_ _17_ 8.82e-21
C309 _44_/a_93_21# _42_/a_109_93# 1.25e-19
C310 input5/a_841_47# net1 1.33e-19
C311 _10_ net2 2.65e-19
C312 _20_ _01_ 0.161f
C313 _01_ _09_ 4.69e-21
C314 _04_ _32_/a_27_47# 1.43e-19
C315 VPWR p[1] 0.08f
C316 net14 _16_ 0.00266f
C317 _30_/a_215_297# _05_ 0.0453f
C318 net14 input3/a_27_47# 3.47e-19
C319 _15_ _55_/a_472_297# 0.00626f
C320 p[12] _06_ 0.0535f
C321 net4 p[12] 0.00758f
C322 _14_ net8 4.23e-19
C323 net5 p[12] 4.79e-20
C324 _43_/a_27_47# net7 6.31e-19
C325 net13 _36_/a_27_47# 0.0488f
C326 _02_ _52_/a_346_47# 0.00526f
C327 _29_/a_29_53# _22_ 2.24e-21
C328 VPWR _50_/a_515_93# -5.03e-19
C329 _13_ _11_ 0.164f
C330 p[10] output17/a_27_47# 0.118f
C331 input5/a_62_47# net2 0.0197f
C332 _52_/a_93_21# net18 8.21e-21
C333 _20_ _30_/a_109_53# 8.12e-19
C334 p[14] net19 0.101f
C335 _10_ p[12] 0.0993f
C336 _44_/a_93_21# _16_ 0.00354f
C337 _11_ net19 2.19e-19
C338 _55_/a_80_21# _55_/a_217_297# 1.42e-32
C339 output19/a_27_47# _06_ 1.53e-19
C340 _01_ _19_ 0.031f
C341 net13 _08_ 1.82e-19
C342 net6 _16_ 1.62e-20
C343 input5/a_62_47# p[8] 1.15e-19
C344 VPWR _43_/a_27_47# 0.0186f
C345 p[5] net10 0.00544f
C346 _37_/a_27_47# _00_ 6.15e-20
C347 _31_/a_35_297# net2 0.0635f
C348 _06_ _55_/a_217_297# 3.46e-19
C349 net4 _55_/a_217_297# 1.13e-19
C350 _27_/a_109_297# _19_ 7.54e-21
C351 net5 _55_/a_217_297# 8.84e-20
C352 net17 net9 1.26e-20
C353 net14 net11 9.95e-19
C354 _10_ output19/a_27_47# 3.23e-20
C355 _00_ net9 0.00501f
C356 _04_ output17/a_27_47# 0.027f
C357 input5/a_381_47# net8 7.48e-19
C358 _29_/a_29_53# _50_/a_27_47# 1.44e-20
C359 _42_/a_109_93# _22_ 1.21e-19
C360 _52_/a_93_21# net4 7.93e-20
C361 _52_/a_93_21# _06_ 0.0574f
C362 _10_ _55_/a_217_297# 1.43e-19
C363 _52_/a_93_21# net5 0.0124f
C364 net8 net7 0.295f
C365 net11 net1 1.13e-19
C366 _25_ _38_/a_27_47# 5.76e-19
C367 _11_ _50_/a_223_47# 0.0329f
C368 input7/a_27_47# net17 4.99e-20
C369 _31_/a_117_297# net8 5.91e-19
C370 input2/a_27_47# _30_/a_109_53# 1.54e-20
C371 _14_ b[3] 1.92e-19
C372 _02_ net17 0.0608f
C373 _35_/a_226_47# net1 1.3e-20
C374 _52_/a_93_21# _10_ 0.00534f
C375 _06_ _40_/a_297_297# 1.64e-19
C376 _14_ _40_/a_191_297# 2.4e-19
C377 _00_ _39_/a_285_47# 1.47e-21
C378 net11 net6 1.08e-19
C379 VPWR net8 0.703f
C380 net6 _23_ 2.13e-19
C381 _02_ _00_ 0.0269f
C382 net16 output16/a_27_47# 0.0101f
C383 net8 p[3] 0.0015f
C384 _44_/a_250_297# net2 0.0169f
C385 _21_ _36_/a_27_47# 0.0276f
C386 _48_/a_181_47# _06_ 6.4e-19
C387 _16_ _22_ 3.8e-19
C388 _13_ _43_/a_193_413# 5.58e-21
C389 _03_ _20_ 0.0794f
C390 net13 net9 0.035f
C391 _03_ _30_/a_297_297# 0.00117f
C392 _35_/a_76_199# net11 4e-19
C393 _49_/a_75_199# net11 4.49e-19
C394 _03_ _09_ 0.326f
C395 input3/a_27_47# _22_ 5.13e-20
C396 net3 net17 3.72e-19
C397 _43_/a_193_413# net19 3.31e-19
C398 _39_/a_47_47# p[12] 3.32e-19
C399 net13 p[4] 2.34e-20
C400 _21_ _08_ 0.00139f
C401 _35_/a_226_47# _49_/a_75_199# 8.73e-20
C402 _00_ net3 2.12e-19
C403 _37_/a_197_47# _15_ 3.02e-19
C404 p[11] b[3] 0.243f
C405 _00_ _17_ 0.0851f
C406 _11_ _24_ 7.29e-20
C407 net13 _02_ 0.00154f
C408 net2 net19 0.599f
C409 _27_/a_27_297# p[1] 2.27e-19
C410 _03_ _19_ 0.0019f
C411 p[5] input10/a_27_47# 0.0172f
C412 _31_/a_285_297# net1 5.85e-19
C413 p[8] net19 0.0268f
C414 _03_ input2/a_27_47# 2.71e-19
C415 _27_/a_205_297# _15_ 5.5e-20
C416 _45_/a_27_47# _11_ 0.0703f
C417 _31_/a_35_297# b[1] 3.21e-19
C418 net11 _22_ 6.82e-21
C419 output19/a_27_47# _44_/a_250_297# 6.42e-20
C420 input13/a_27_47# net9 2.42e-19
C421 _23_ _22_ 0.0186f
C422 VPWR b[3] 0.367f
C423 net15 p[1] 6.22e-20
C424 _29_/a_29_53# _06_ 0.00111f
C425 VPWR _40_/a_191_297# -6.82e-19
C426 net13 net3 3.25e-21
C427 _35_/a_226_47# _22_ 1.39e-20
C428 net5 _29_/a_29_53# 8.1e-20
C429 p[12] net19 6.8e-20
C430 input13/a_27_47# p[4] 7.37e-20
C431 _01_ net17 0.0988f
C432 _15_ _42_/a_209_311# 0.0521f
C433 _52_/a_93_21# _39_/a_47_47# 1.44e-20
C434 input10/a_27_47# net10 0.00321f
C435 _14_ p[14] 1.66e-20
C436 net13 _49_/a_201_297# 3.31e-19
C437 _33_/a_109_93# net9 0.00211f
C438 VPWR _33_/a_209_311# -0.0131f
C439 _01_ _00_ 0.00124f
C440 _14_ _11_ 0.0415f
C441 input1/a_75_212# net1 0.00208f
C442 _43_/a_369_47# _18_ 1.49e-19
C443 _21_ net9 0.0282f
C444 _10_ _29_/a_29_53# 5.17e-19
C445 net12 net8 0.00458f
C446 _07_ net1 6.08e-22
C447 input8/a_27_47# net1 0.0347f
C448 _26_/a_29_53# _11_ 1.09e-19
C449 _05_ net1 0.151f
C450 net11 _50_/a_27_47# 6.05e-21
C451 output19/a_27_47# net19 0.0279f
C452 p[2] _31_/a_285_297# 0.00156f
C453 _09_ _29_/a_183_297# 4.51e-20
C454 net11 _12_ 0.00799f
C455 _30_/a_109_53# net17 4.18e-20
C456 _20_ net10 3.23e-19
C457 b[0] b[2] 0.183f
C458 _12_ _23_ 0.00743f
C459 _09_ net10 0.037f
C460 _30_/a_297_297# net10 1.68e-19
C461 net16 _09_ 0.00707f
C462 _00_ _30_/a_109_53# 3.67e-20
C463 _06_ _42_/a_109_93# 5.53e-20
C464 _02_ _33_/a_109_93# 1.54e-21
C465 _35_/a_226_47# _12_ 8.38e-20
C466 _52_/a_93_21# _13_ 1.31e-19
C467 net5 _42_/a_109_93# 0.00109f
C468 input14/a_27_47# p[13] 1.37e-19
C469 _15_ _18_ 0.042f
C470 _02_ _21_ 0.397f
C471 _27_/a_27_297# net8 0.0108f
C472 p[11] p[14] 3.13e-20
C473 input8/a_27_47# _49_/a_75_199# 1.99e-20
C474 input5/a_841_47# _06_ 1.66e-19
C475 net13 _01_ 0.00228f
C476 _35_/a_76_199# _07_ 0.00226f
C477 _49_/a_75_199# _07_ 4.05e-21
C478 net14 _37_/a_197_47# 7e-19
C479 _45_/a_193_297# _23_ 4.13e-19
C480 _35_/a_76_199# _05_ 0.00238f
C481 p[11] _11_ 4.18e-20
C482 _14_ _55_/a_300_47# 8.09e-19
C483 net5 input5/a_841_47# 0.0221f
C484 VPWR _52_/a_256_47# -9.47e-19
C485 net13 _34_/a_47_47# 1.68e-19
C486 _28_/a_109_297# b[3] 7.49e-20
C487 _35_/a_226_47# _45_/a_193_297# 8.15e-21
C488 _47_/a_81_21# _18_ 7.96e-20
C489 p[2] _05_ 3.69e-19
C490 input8/a_27_47# p[2] 0.0159f
C491 _55_/a_80_21# _16_ 0.0143f
C492 net14 _27_/a_205_297# 3.63e-19
C493 net15 net8 0.2f
C494 _21_ _35_/a_556_47# 2.69e-19
C495 net4 _16_ 2.73e-20
C496 _16_ _06_ 0.00162f
C497 net11 input11/a_27_47# 0.00318f
C498 input2/a_27_47# net10 1.17e-20
C499 net13 _30_/a_109_53# 1.05e-19
C500 net5 _16_ 1.99e-20
C501 VPWR p[14] 0.0416f
C502 input14/a_27_47# net3 9.36e-19
C503 _02_ _52_/a_250_297# 0.0128f
C504 VPWR _11_ 0.352f
C505 _14_ _43_/a_193_413# 0.0297f
C506 net11 net18 0.00221f
C507 net14 _42_/a_209_311# 0.0238f
C508 _10_ _16_ 0.00486f
C509 _02_ _53_/a_29_53# 0.0388f
C510 _38_/a_27_47# _22_ 2.86e-19
C511 _07_ _22_ 1.19e-20
C512 _03_ net17 5.1e-19
C513 net12 _33_/a_209_311# 0.0769f
C514 _05_ _22_ 3.33e-21
C515 _03_ _00_ 2.31e-20
C516 _14_ net2 0.0104f
C517 _30_/a_215_297# _04_ 0.00225f
C518 input9/a_75_212# _29_/a_29_53# 9.7e-21
C519 _34_/a_129_47# net10 0.003f
C520 _39_/a_377_297# _11_ 2.57e-20
C521 net8 _50_/a_343_93# 7.25e-19
C522 _44_/a_93_21# _42_/a_209_311# 2.21e-19
C523 net11 _06_ 0.546f
C524 net6 _42_/a_209_311# 1.32e-20
C525 input5/a_558_47# _15_ 0.00166f
C526 _06_ _23_ 0.218f
C527 VPWR _55_/a_300_47# -4.61e-19
C528 input5/a_62_47# input3/a_27_47# 0.00179f
C529 _21_ _01_ 7.94e-19
C530 net5 net11 0.0129f
C531 net5 _23_ 0.0052f
C532 _36_/a_27_47# net8 1.52e-19
C533 _21_ _34_/a_47_47# 8.93e-19
C534 _50_/a_27_47# _38_/a_27_47# 2.37e-20
C535 _12_ _38_/a_27_47# 0.0527f
C536 _12_ _07_ 2.94e-23
C537 net14 _18_ 0.0147f
C538 _12_ _05_ 2.52e-19
C539 _35_/a_226_47# _06_ 0.00487f
C540 _43_/a_193_413# net7 3.49e-19
C541 _10_ net11 0.0109f
C542 _02_ _52_/a_584_47# 0.00389f
C543 net15 b[3] 0.00408f
C544 net13 _36_/a_109_47# 0.00126f
C545 _37_/a_109_47# net19 1.16e-20
C546 VPWR _50_/a_615_93# -5.34e-19
C547 _10_ _23_ 0.00192f
C548 _52_/a_93_21# _24_ 0.0211f
C549 p[11] net2 0.0204f
C550 _28_/a_109_297# _11_ 6.29e-19
C551 _03_ net13 0.271f
C552 net15 _40_/a_191_297# 8.41e-19
C553 input5/a_381_47# net2 0.0138f
C554 _44_/a_250_297# _42_/a_109_93# 6.38e-19
C555 input7/a_27_47# p[1] 0.0164f
C556 _21_ _30_/a_109_53# 3.31e-20
C557 _20_ _09_ 7.11e-19
C558 _10_ _35_/a_226_47# 1.25e-19
C559 _45_/a_193_297# _05_ 4.84e-22
C560 net2 net7 0.00234f
C561 output19/a_27_47# _14_ 1.43e-19
C562 _49_/a_544_297# _04_ 0.00204f
C563 _44_/a_93_21# _18_ 0.00485f
C564 _15_ _32_/a_27_47# 1.19e-19
C565 _45_/a_27_47# _52_/a_93_21# 1.18e-19
C566 VPWR _43_/a_193_413# 0.0063f
C567 p[11] p[8] 0.0023f
C568 _48_/a_27_47# _06_ 0.0251f
C569 net6 _18_ 0.166f
C570 _04_ _15_ 3.61e-20
C571 _14_ _55_/a_217_297# 0.0116f
C572 net12 _11_ 3.82e-21
C573 _41_/a_145_75# p[12] 0.00339f
C574 _47_/a_81_21# _32_/a_27_47# 5.06e-21
C575 VPWR net2 0.918f
C576 _34_/a_47_47# _53_/a_29_53# 5.88e-22
C577 _41_/a_59_75# _15_ 0.0139f
C578 _29_/a_29_53# _50_/a_223_47# 1.45e-20
C579 _20_ _19_ 0.00734f
C580 _44_/a_250_297# _16_ 3.25e-19
C581 _10_ _55_/a_472_297# 7.35e-21
C582 _35_/a_76_199# _18_ 6.82e-21
C583 _42_/a_209_311# _22_ 1.72e-19
C584 _10_ _48_/a_27_47# 4.55e-19
C585 _42_/a_109_93# net19 0.0448f
C586 _31_/a_285_297# _06_ 1.01e-20
C587 net17 net10 8.67e-21
C588 _09_ _19_ 4.8e-21
C589 VPWR p[8] 0.208f
C590 VPWR input12/a_27_47# 0.0646f
C591 _02_ _43_/a_27_47# 1.88e-21
C592 _44_/a_250_297# input3/a_27_47# 2.07e-19
C593 net18 _38_/a_27_47# 0.00997f
C594 input12/a_27_47# p[6] 0.0166f
C595 _37_/a_27_47# net8 6.66e-21
C596 _41_/a_59_75# _47_/a_81_21# 1.5e-19
C597 _37_/a_303_47# net2 4.41e-19
C598 _14_ _40_/a_297_297# 1.58e-19
C599 VPWR p[12] 0.0375f
C600 net13 p[5] 1.05e-19
C601 net8 net9 0.0605f
C602 _03_ _33_/a_109_93# 2.78e-19
C603 net14 input5/a_558_47# 0.0325f
C604 b[2] _25_ 0.0015f
C605 _03_ _21_ 0.0818f
C606 _16_ net19 0.206f
C607 _39_/a_47_47# _23_ 5.24e-21
C608 _55_/a_217_297# net7 1.04e-19
C609 _06_ _38_/a_27_47# 0.0172f
C610 net4 _38_/a_27_47# 0.0119f
C611 p[10] net14 3.02e-19
C612 _21_ _34_/a_377_297# 2.37e-19
C613 _06_ _07_ 0.185f
C614 _43_/a_27_47# _17_ 0.00131f
C615 input3/a_27_47# net19 0.00105f
C616 input5/a_558_47# net1 1.1e-19
C617 _18_ _22_ 0.0211f
C618 net15 p[14] 0.00132f
C619 input7/a_27_47# net8 2.03e-21
C620 input2/a_27_47# _19_ 5.26e-20
C621 p[13] net8 0.00345f
C622 _06_ _05_ 0.00724f
C623 _08_ _33_/a_209_311# 0.0122f
C624 net5 _38_/a_27_47# 1.76e-19
C625 output19/a_27_47# VPWR 0.0229f
C626 net15 _11_ 0.145f
C627 net11 input9/a_75_212# 1.1e-20
C628 input6/a_27_47# b[3] 4.02e-19
C629 net13 net10 0.375f
C630 b[3] input15/a_27_47# 1.77e-19
C631 p[10] net1 1.22e-19
C632 _44_/a_93_21# input5/a_558_47# 2.71e-19
C633 _02_ net8 0.334f
C634 VPWR _55_/a_217_297# -0.00133f
C635 _10_ _38_/a_27_47# 0.0133f
C636 _10_ _05_ 9.25e-21
C637 p[11] b[1] 1.84e-20
C638 _26_/a_183_297# _00_ 4.53e-19
C639 _10_ _07_ 2.19e-19
C640 p[7] net1 7.5e-20
C641 input13/a_27_47# p[5] 3.09e-19
C642 net14 _04_ 0.0863f
C643 net11 _13_ 2.34e-19
C644 _52_/a_93_21# VPWR -0.00838f
C645 _13_ _23_ 2.08e-20
C646 b[1] net7 0.005f
C647 _11_ _50_/a_343_93# 0.0384f
C648 _31_/a_117_297# b[1] 2.34e-19
C649 _32_/a_27_47# net1 0.0211f
C650 _50_/a_27_47# _18_ 0.0665f
C651 _45_/a_109_297# _11_ 0.00168f
C652 _12_ _18_ 0.0115f
C653 net3 net8 9.23e-19
C654 input5/a_664_47# _42_/a_209_311# 0.0124f
C655 _35_/a_226_47# _13_ 5.62e-21
C656 _01_ _43_/a_27_47# 9.77e-20
C657 _04_ net1 0.018f
C658 net15 _55_/a_300_47# 1.09e-19
C659 p[10] _49_/a_75_199# 2.29e-20
C660 _17_ net8 4.52e-20
C661 net12 input12/a_27_47# 0.0295f
C662 _49_/a_201_297# net8 7.3e-19
C663 VPWR b[1] 0.396f
C664 VPWR _40_/a_297_297# -5.42e-19
C665 _40_/a_109_297# net6 2.53e-20
C666 _44_/a_93_21# _04_ 4.47e-21
C667 input13/a_27_47# net10 8.86e-20
C668 _26_/a_29_53# _29_/a_29_53# 0.00121f
C669 _04_ net6 2.61e-20
C670 _33_/a_209_311# net9 4.33e-20
C671 input8/a_27_47# _31_/a_35_297# 0.00955f
C672 VPWR _48_/a_181_47# -3.35e-19
C673 b[3] p[13] 0.165f
C674 _27_/a_27_297# net2 0.0131f
C675 _06_ _33_/a_296_53# 1.11e-20
C676 _31_/a_35_297# _05_ 0.00649f
C677 _41_/a_59_75# net6 0.0373f
C678 _02_ b[3] 1.07e-19
C679 net13 _36_/a_197_47# 1.06e-19
C680 _49_/a_75_199# _04_ 0.0782f
C681 net10 _33_/a_109_93# 0.0336f
C682 _35_/a_76_199# _04_ 0.0269f
C683 _20_ net17 4e-20
C684 _21_ net10 0.0254f
C685 _55_/a_80_21# _42_/a_209_311# 0.0175f
C686 _21_ net16 1.89e-19
C687 net15 _43_/a_193_413# 0.00169f
C688 input5/a_664_47# _18_ 1.09e-20
C689 _20_ _00_ 0.271f
C690 _49_/a_208_47# net7 0.00312f
C691 _06_ _42_/a_209_311# 1.66e-19
C692 _00_ _09_ 9.35e-21
C693 p[2] _04_ 1.83e-20
C694 output17/a_27_47# net1 8.12e-19
C695 _14_ _42_/a_109_93# 0.00141f
C696 _01_ net8 0.0802f
C697 input6/a_27_47# p[14] 0.0155f
C698 _37_/a_109_47# p[11] 2.84e-20
C699 net5 _42_/a_209_311# 3.27e-21
C700 b[3] _44_/a_584_47# 0.00109f
C701 input15/a_27_47# p[14] 6.15e-19
C702 net15 net2 0.324f
C703 input15/a_27_47# _11_ 4.4e-19
C704 _29_/a_29_53# net7 6.01e-19
C705 net3 b[3] 0.0026f
C706 VPWR _49_/a_208_47# -5.93e-19
C707 net3 _40_/a_191_297# 1.89e-19
C708 net15 p[8] 3.39e-19
C709 input9/a_75_212# _05_ 1.24e-21
C710 input8/a_27_47# input9/a_75_212# 3.09e-20
C711 b[3] _17_ 0.00637f
C712 net17 _19_ 0.0211f
C713 _32_/a_27_47# _22_ 1.76e-19
C714 _37_/a_27_47# p[14] 1.37e-19
C715 _30_/a_109_53# net8 1.76e-20
C716 _40_/a_191_297# _17_ 4.35e-19
C717 net10 _52_/a_250_297# 2.86e-21
C718 VPWR _29_/a_29_53# 0.0299f
C719 _55_/a_80_21# _18_ 1.44e-20
C720 _04_ _22_ 1.76e-20
C721 VPWR _37_/a_109_47# -4.38e-19
C722 _37_/a_27_47# _11_ 0.0018f
C723 input2/a_27_47# net17 0.0398f
C724 _29_/a_29_53# p[3] 2.07e-19
C725 _14_ _16_ 0.0584f
C726 net2 _50_/a_343_93# 1.25e-20
C727 net13 _20_ 5.95e-19
C728 _54_/a_75_212# _25_ 0.0247f
C729 net15 p[12] 2.99e-19
C730 net13 _30_/a_297_297# 3.27e-20
C731 net13 _09_ 0.0379f
C732 _53_/a_29_53# net10 7.88e-22
C733 net16 _53_/a_29_53# 2.04e-20
C734 _06_ _18_ 0.54f
C735 net4 _18_ 0.023f
C736 _13_ _38_/a_27_47# 4.58e-19
C737 _24_ _23_ 0.012f
C738 _41_/a_59_75# _22_ 6.24e-22
C739 _11_ net9 5.39e-19
C740 _13_ _07_ 3.22e-23
C741 p[11] _42_/a_109_93# 4.55e-21
C742 input5/a_381_47# _42_/a_109_93# 0.00763f
C743 _13_ _05_ 2.57e-20
C744 _02_ _52_/a_256_47# 0.00344f
C745 net5 _18_ 0.0426f
C746 _45_/a_27_47# net11 3.64e-20
C747 _45_/a_27_47# _23_ 1.74e-19
C748 output19/a_27_47# net15 6.88e-19
C749 _10_ _18_ 0.133f
C750 _01_ b[3] 9.26e-20
C751 input5/a_841_47# net7 0.00193f
C752 net15 _55_/a_217_297# 7.79e-19
C753 _04_ _12_ 1.42e-19
C754 _04_ _50_/a_27_47# 2.07e-21
C755 net13 _19_ 4.45e-20
C756 _45_/a_27_47# _35_/a_226_47# 5.71e-21
C757 VPWR _42_/a_109_93# -0.00118f
C758 _02_ _11_ 0.0621f
C759 b[2] _22_ 0.0043f
C760 _16_ p[11] 2.17e-20
C761 _41_/a_59_75# _50_/a_27_47# 9.59e-22
C762 _41_/a_59_75# _12_ 0.00101f
C763 VPWR input5/a_841_47# 0.0775f
C764 p[11] input3/a_27_47# 0.0157f
C765 input15/a_27_47# _43_/a_193_413# 1.62e-20
C766 input13/a_27_47# _09_ 1.27e-21
C767 _34_/a_47_47# _33_/a_209_311# 0.017f
C768 _16_ net7 7.5e-20
C769 net11 _26_/a_29_53# 1.08e-20
C770 _03_ net8 0.0287f
C771 _35_/a_489_413# _06_ 9.22e-19
C772 _12_ _38_/a_109_47# 0.00179f
C773 net11 _29_/a_111_297# 8.27e-19
C774 input6/a_27_47# net2 0.0047f
C775 input15/a_27_47# net2 0.00296f
C776 net3 p[14] 0.00446f
C777 b[0] net6 2.52e-19
C778 net15 _40_/a_297_297# 4.08e-19
C779 net3 _11_ 0.165f
C780 _20_ _21_ 0.191f
C781 _09_ _33_/a_109_93# 7.36e-20
C782 _37_/a_27_47# _43_/a_193_413# 0.0102f
C783 VPWR _16_ 0.126f
C784 _17_ p[14] 5.46e-21
C785 net11 output18/a_27_47# 6.84e-20
C786 input6/a_27_47# p[8] 0.00139f
C787 _11_ _17_ 0.197f
C788 input5/a_664_47# _04_ 6.73e-21
C789 VPWR input3/a_27_47# 0.0687f
C790 _12_ b[2] 3.89e-20
C791 _10_ _35_/a_489_413# 3.41e-19
C792 _21_ _09_ 0.263f
C793 input15/a_27_47# p[8] 7.57e-19
C794 input5/a_558_47# _06_ 3.55e-19
C795 _02_ _55_/a_300_47# 0.00371f
C796 input14/a_27_47# p[9] 8.53e-21
C797 net12 _29_/a_29_53# 0.0132f
C798 net5 input5/a_558_47# 0.0597f
C799 _37_/a_27_47# net2 0.0692f
C800 net5 _32_/a_109_47# 5.69e-21
C801 _14_ _55_/a_472_297# 0.00192f
C802 input6/a_27_47# p[12] 2.78e-19
C803 p[12] input15/a_27_47# 5.48e-19
C804 p[10] net5 5.12e-21
C805 _37_/a_27_47# p[8] 9.82e-21
C806 net2 net9 3.64e-20
C807 net11 net7 1.77e-19
C808 _39_/a_47_47# _18_ 1.23e-19
C809 _42_/a_209_311# net19 0.0766f
C810 _07_ _24_ 5.67e-19
C811 _35_/a_226_47# net7 2.93e-20
C812 _06_ p[7] 0.00864f
C813 _02_ _43_/a_193_413# 9.4e-21
C814 _09_ _52_/a_250_297# 1.97e-20
C815 output19/a_27_47# input6/a_27_47# 0.107f
C816 _40_/a_109_297# _06_ 0.00175f
C817 p[0] p[1] 0.187f
C818 _06_ _32_/a_27_47# 0.00663f
C819 VPWR net11 0.996f
C820 _41_/a_59_75# _47_/a_299_297# 0.00146f
C821 input7/a_27_47# net2 3.24e-19
C822 net11 p[6] 0.0099f
C823 p[13] net2 0.0247f
C824 VPWR _23_ -0.00374f
C825 net5 _32_/a_27_47# 0.0961f
C826 _04_ _06_ 0.0136f
C827 _09_ _53_/a_29_53# 0.00642f
C828 input12/a_27_47# p[4] 8.26e-19
C829 _45_/a_27_47# _05_ 9.34e-23
C830 VPWR _35_/a_226_47# 0.00159f
C831 net5 _04_ 0.00476f
C832 _45_/a_27_47# _07_ 1.02e-20
C833 p[13] p[8] 0.00172f
C834 _47_/a_384_47# _15_ 0.00112f
C835 _03_ _33_/a_209_311# 8.38e-19
C836 _28_/a_109_297# _16_ 1.26e-19
C837 _10_ _32_/a_27_47# 0.00217f
C838 b[2] net18 0.0131f
C839 _41_/a_59_75# _06_ 0.0429f
C840 _13_ _18_ 0.019f
C841 _47_/a_81_21# _15_ 0.00332f
C842 _41_/a_59_75# net4 1.76e-19
C843 _41_/a_59_75# net5 2.41e-19
C844 _10_ _04_ 9.24e-20
C845 net10 net8 2.05e-21
C846 _02_ input12/a_27_47# 1.88e-19
C847 net3 _43_/a_193_413# 5.65e-20
C848 _44_/a_584_47# net2 0.0053f
C849 net4 _38_/a_109_47# 7.32e-19
C850 _18_ net19 4.89e-20
C851 _43_/a_193_413# _17_ 0.0503f
C852 _32_/a_197_47# net1 0.00142f
C853 p[10] _31_/a_35_297# 2.29e-19
C854 net13 net17 5.21e-20
C855 _27_/a_27_297# _42_/a_109_93# 1.35e-20
C856 _10_ _41_/a_59_75# 0.0172f
C857 _01_ _55_/a_300_47# 0.00113f
C858 net3 net2 0.519f
C859 b[0] _12_ 2.61e-20
C860 VPWR _48_/a_27_47# 0.0158f
C861 p[6] _48_/a_27_47# 2.22e-19
C862 VPWR _55_/a_472_297# 0.00488f
C863 _17_ net2 0.181f
C864 _31_/a_285_297# net7 0.00227f
C865 _30_/a_215_297# net1 0.00375f
C866 _32_/a_303_47# net1 1.45e-19
C867 b[2] _06_ 0.0116f
C868 _10_ _38_/a_109_47# 5.44e-19
C869 input5/a_62_47# _04_ 0.00345f
C870 net3 p[8] 2.53e-19
C871 net5 b[2] 7.33e-20
C872 net5 output17/a_27_47# 5.01e-20
C873 output18/a_27_47# _38_/a_27_47# 8.6e-19
C874 net14 _43_/a_369_47# 6.79e-21
C875 _31_/a_35_297# _32_/a_27_47# 9.17e-20
C876 _30_/a_215_297# net6 3.3e-21
C877 net15 _42_/a_109_93# 4.62e-19
C878 VPWR _31_/a_285_297# 0.0174f
C879 _50_/a_223_47# _18_ 0.0367f
C880 _31_/a_35_297# _04_ 1.89e-20
C881 _27_/a_27_297# _16_ 3.74e-22
C882 _01_ _43_/a_193_413# 8.16e-19
C883 _29_/a_29_53# _36_/a_27_47# 6.92e-20
C884 _42_/a_296_53# _15_ 1.28e-19
C885 net15 input5/a_841_47# 0.00585f
C886 _02_ _55_/a_217_297# 6.01e-19
C887 input1/a_75_212# net7 3.77e-19
C888 net11 net12 0.358f
C889 net12 _23_ 2.28e-21
C890 _05_ net7 0.0129f
C891 input8/a_27_47# net7 1.47e-19
C892 _01_ net2 2.72e-19
C893 net6 _43_/a_369_47# 3.62e-21
C894 _52_/a_93_21# _02_ 0.0957f
C895 net14 _15_ 0.225f
C896 output19/a_27_47# net3 0.00348f
C897 _35_/a_226_47# net12 8.29e-19
C898 _20_ _43_/a_27_47# 0.0124f
C899 VPWR input1/a_75_212# 0.0786f
C900 input5/a_62_47# output17/a_27_47# 1.02e-19
C901 _27_/a_109_297# net2 7.24e-20
C902 _06_ _33_/a_368_53# 1.7e-19
C903 net15 _16_ 0.214f
C904 _19_ p[1] 2.82e-20
C905 input9/a_75_212# p[7] 0.00102f
C906 p[13] b[1] 0.00115f
C907 _49_/a_544_297# net1 0.00175f
C908 net15 input3/a_27_47# 6.19e-20
C909 VPWR _38_/a_27_47# -0.0142f
C910 output19/a_27_47# _17_ 0.00122f
C911 input8/a_27_47# VPWR 0.0863f
C912 VPWR _05_ 0.127f
C913 VPWR _07_ 0.0728f
C914 net10 _33_/a_209_311# 0.0419f
C915 net3 _55_/a_217_297# 5.78e-20
C916 _05_ p[3] 5.83e-21
C917 input8/a_27_47# p[3] 0.0023f
C918 input5/a_558_47# net19 2.24e-20
C919 p[6] _07_ 1.26e-19
C920 net13 _36_/a_303_47# 5.5e-20
C921 input12/a_27_47# _34_/a_47_47# 2.17e-19
C922 input2/a_27_47# p[1] 0.0119f
C923 _21_ _00_ 9.26e-20
C924 _04_ input9/a_75_212# 7.69e-22
C925 _44_/a_250_297# _04_ 5.57e-21
C926 net11 _27_/a_27_297# 1.58e-20
C927 p[10] net19 1.26e-21
C928 _14_ _42_/a_209_311# 0.00142f
C929 _44_/a_93_21# _15_ 0.0168f
C930 _37_/a_197_47# p[11] 1.59e-19
C931 net14 _44_/a_346_47# 0.00464f
C932 _47_/a_81_21# net1 1.58e-21
C933 net6 _15_ 0.17f
C934 _30_/a_215_297# _22_ 2.46e-21
C935 _02_ _48_/a_181_47# 3.9e-19
C936 net12 _48_/a_27_47# 0.0126f
C937 net13 input13/a_27_47# 0.00139f
C938 net4 b[0] 0.0024f
C939 _13_ _04_ 1.17e-21
C940 _45_/a_27_47# _18_ 0.00347f
C941 net3 _40_/a_297_297# 2.54e-19
C942 net5 b[0] 2.76e-19
C943 net6 _47_/a_81_21# 2.14e-19
C944 _20_ net8 5.07e-19
C945 _30_/a_297_297# net8 2.42e-21
C946 net10 _52_/a_256_47# 8.13e-20
C947 _44_/a_93_21# _44_/a_346_47# -5.12e-20
C948 _04_ net19 2.07e-20
C949 net13 _33_/a_109_93# 0.0254f
C950 VPWR _37_/a_197_47# -3.27e-19
C951 _01_ _55_/a_217_297# 0.00112f
C952 _29_/a_29_53# net9 0.0205f
C953 net13 _21_ 0.13f
C954 _54_/a_75_212# net18 0.0143f
C955 _27_/a_277_297# _04_ 0.00113f
C956 net14 _42_/a_296_53# 2.18e-19
C957 _14_ _18_ 0.243f
C958 input5/a_381_47# _42_/a_209_311# 3.88e-19
C959 _41_/a_59_75# net19 3.1e-20
C960 _02_ _49_/a_208_47# 0.00193f
C961 VPWR _33_/a_296_53# -1.15e-19
C962 _26_/a_29_53# _18_ 5.26e-20
C963 VPWR _27_/a_205_297# 1.05e-19
C964 _19_ net8 0.0322f
C965 _45_/a_109_297# net11 7.46e-20
C966 _34_/a_285_47# _06_ 0.00598f
C967 _37_/a_27_47# _42_/a_109_93# 2.55e-20
C968 net16 _11_ 0.172f
C969 _02_ _29_/a_29_53# 6.76e-21
C970 _03_ net2 1.89e-19
C971 _15_ _22_ 0.0236f
C972 _25_ _22_ 5.39e-19
C973 _04_ _50_/a_223_47# 7.89e-22
C974 input2/a_27_47# net8 0.0207f
C975 net12 _07_ 0.18f
C976 _54_/a_75_212# _06_ 0.00727f
C977 net12 _05_ 0.0414f
C978 _45_/a_109_297# _35_/a_226_47# 1.59e-21
C979 VPWR _42_/a_209_311# -0.00753f
C980 _45_/a_27_47# _35_/a_489_413# 3.89e-21
C981 _37_/a_27_47# input5/a_841_47# 4.64e-20
C982 _16_ input15/a_27_47# 7.13e-19
C983 net14 net1 6.64e-20
C984 input13/a_27_47# _33_/a_109_93# 0.00348f
C985 net11 _36_/a_27_47# 0.0717f
C986 _47_/a_81_21# _22_ 7.25e-19
C987 _36_/a_27_47# _23_ 0.00118f
C988 _20_ b[3] 1.37e-19
C989 input5/a_841_47# net9 2.7e-19
C990 p[9] b[3] 0.0898f
C991 net14 _44_/a_93_21# 0.0646f
C992 net14 net6 2.82e-21
C993 _37_/a_109_47# net3 0.00212f
C994 net3 _29_/a_29_53# 1.68e-20
C995 _20_ _40_/a_191_297# 2.07e-20
C996 _18_ net7 2.58e-20
C997 net11 _08_ 8.83e-19
C998 _37_/a_109_47# _17_ 8.86e-21
C999 _37_/a_27_47# _16_ 2.07e-19
C1000 _08_ _23_ 1.81e-19
C1001 net17 p[1] 6.65e-20
C1002 _21_ _33_/a_109_93# 1.62e-20
C1003 _15_ _50_/a_27_47# 5.65e-19
C1004 _12_ _25_ 1.23e-20
C1005 _12_ _15_ 0.00833f
C1006 _09_ _33_/a_209_311# 3.79e-20
C1007 net14 _49_/a_75_199# 3.67e-19
C1008 _35_/a_226_47# _08_ 0.00117f
C1009 net12 _30_/a_392_297# 2.19e-20
C1010 input5/a_841_47# p[13] 1.73e-19
C1011 _12_ _47_/a_384_47# 9.51e-20
C1012 _02_ input5/a_841_47# 0.00591f
C1013 _39_/a_47_47# b[0] 2.04e-19
C1014 VPWR _18_ 0.0721f
C1015 _44_/a_93_21# net6 1.08e-20
C1016 _12_ _47_/a_81_21# 0.00158f
C1017 _49_/a_75_199# net1 0.00799f
C1018 net5 _32_/a_197_47# 5.61e-21
C1019 _01_ _49_/a_208_47# 2.13e-19
C1020 net3 _42_/a_109_93# 0.0435f
C1021 _30_/a_215_297# _06_ 2.03e-20
C1022 input3/a_27_47# p[13] 0.00499f
C1023 p[2] net1 0.0269f
C1024 net5 _30_/a_215_297# 8.27e-21
C1025 net12 _33_/a_296_53# 1.23e-20
C1026 _42_/a_109_93# _17_ 7.83e-20
C1027 _02_ _16_ 0.00564f
C1028 net5 _32_/a_303_47# 7.18e-21
C1029 _00_ _43_/a_27_47# 0.0431f
C1030 p[5] input12/a_27_47# 0.00359f
C1031 _01_ _29_/a_29_53# 8.33e-20
C1032 _52_/a_250_297# _33_/a_109_93# 5.17e-22
C1033 _35_/a_76_199# net6 4.6e-21
C1034 _48_/a_27_47# _08_ 2.58e-19
C1035 _03_ _52_/a_93_21# 0.00985f
C1036 input5/a_664_47# _15_ 9.15e-22
C1037 _04_ _49_/a_315_47# 7.71e-19
C1038 net10 net2 2.05e-20
C1039 b[0] _13_ 0.00299f
C1040 _10_ _30_/a_215_297# 5.66e-20
C1041 net14 _22_ 2.23e-19
C1042 net11 net9 0.136f
C1043 _21_ _53_/a_29_53# 0.00959f
C1044 _40_/a_109_297# _14_ -1.78e-33
C1045 _23_ net9 1.21e-19
C1046 _03_ b[1] 0.00143f
C1047 _43_/a_369_47# _06_ -2.02e-19
C1048 _25_ net18 0.0594f
C1049 input12/a_27_47# net10 0.00182f
C1050 _14_ _04_ 2.04e-21
C1051 b[2] _24_ 1.85e-19
C1052 net11 p[4] 0.0557f
C1053 _45_/a_109_297# _05_ 2.79e-22
C1054 _30_/a_109_53# _29_/a_29_53# 0.0103f
C1055 VPWR _35_/a_489_413# -0.00725f
C1056 net3 _16_ 1.77e-19
C1057 net1 _22_ 0.0129f
C1058 p[2] _49_/a_75_199# 1.06e-19
C1059 _35_/a_226_47# net9 1.22e-20
C1060 _26_/a_29_53# _04_ 2.3e-21
C1061 net3 input3/a_27_47# 0.03f
C1062 input5/a_558_47# net7 0.00358f
C1063 p[9] p[14] 0.4f
C1064 p[10] p[11] 0.00241f
C1065 _37_/a_197_47# net15 1.78e-19
C1066 _16_ _17_ 0.242f
C1067 _47_/a_299_297# _15_ 0.0103f
C1068 _20_ _11_ 0.268f
C1069 net17 net8 0.18f
C1070 _04_ _29_/a_111_297# 9.25e-19
C1071 _10_ _43_/a_369_47# 0.00199f
C1072 _09_ _11_ 0.0665f
C1073 p[9] _11_ 1.01e-19
C1074 input4/a_75_212# p[12] 0.02f
C1075 net6 _22_ 0.163f
C1076 p[10] net7 0.00481f
C1077 _36_/a_27_47# _05_ 3.67e-21
C1078 _55_/a_80_21# _15_ 0.107f
C1079 _02_ net11 0.0327f
C1080 _39_/a_285_47# _23_ 1.9e-20
C1081 _00_ net8 3.23e-19
C1082 _02_ _23_ 0.0641f
C1083 VPWR input5/a_558_47# 0.0083f
C1084 _27_/a_27_297# _42_/a_209_311# 4.7e-20
C1085 VPWR _32_/a_109_47# 0.00124f
C1086 _06_ _25_ 0.144f
C1087 _15_ _06_ 0.22f
C1088 net4 _15_ 0.00427f
C1089 _31_/a_35_297# _30_/a_215_297# 6.37e-19
C1090 _02_ _35_/a_226_47# 2.21e-19
C1091 net5 _25_ 6.42e-19
C1092 _35_/a_76_199# _22_ 6.58e-21
C1093 _49_/a_75_199# _22_ 9.85e-21
C1094 net12 _18_ 2.25e-21
C1095 net5 _15_ 0.0352f
C1096 _31_/a_285_47# net7 0.00132f
C1097 VPWR p[10] 0.177f
C1098 _08_ _05_ 0.00897f
C1099 _08_ _07_ 0.348f
C1100 net5 _47_/a_384_47# 0.00129f
C1101 _32_/a_27_47# net7 0.00559f
C1102 _47_/a_81_21# _06_ 0.0388f
C1103 net5 _47_/a_81_21# 4.59e-19
C1104 _10_ _25_ 0.0109f
C1105 _10_ _15_ 0.479f
C1106 _04_ net7 0.0602f
C1107 net15 _42_/a_209_311# 0.0157f
C1108 _01_ _16_ 3.24e-19
C1109 VPWR p[7] 0.0184f
C1110 _03_ _49_/a_208_47# 3.86e-19
C1111 net6 _50_/a_27_47# 0.0428f
C1112 _10_ _47_/a_384_47# 3.53e-19
C1113 _12_ net6 0.0891f
C1114 p[7] p[3] 0.169f
C1115 p[6] p[7] 0.217f
C1116 VPWR _31_/a_285_47# -2.91e-19
C1117 _49_/a_201_297# net11 1.42e-19
C1118 net13 net8 7.51e-20
C1119 VPWR _32_/a_27_47# 0.0395f
C1120 VPWR _40_/a_109_297# -4.23e-19
C1121 _02_ _48_/a_27_47# 0.00435f
C1122 _10_ _47_/a_81_21# 0.0061f
C1123 _52_/a_93_21# net10 7.84e-20
C1124 _02_ _55_/a_472_297# 1.25e-19
C1125 VPWR _04_ 0.456f
C1126 _49_/a_201_297# _35_/a_226_47# 1.66e-20
C1127 _03_ _29_/a_29_53# 0.0414f
C1128 net14 input5/a_664_47# 0.0179f
C1129 output18/a_27_47# b[2] 0.0141f
C1130 _04_ p[3] 8.93e-22
C1131 _35_/a_76_199# _12_ 6.84e-20
C1132 _20_ _50_/a_615_93# 8.8e-19
C1133 net6 _45_/a_193_297# 9.84e-20
C1134 _30_/a_215_297# input9/a_75_212# 6.24e-21
C1135 _10_ _44_/a_346_47# 9.13e-21
C1136 _00_ b[3] 1.04e-19
C1137 VPWR _41_/a_59_75# 0.0179f
C1138 input5/a_664_47# net1 2.41e-19
C1139 _02_ _31_/a_285_297# 5.86e-20
C1140 _35_/a_489_413# net12 3.97e-20
C1141 _20_ _43_/a_193_413# 0.00161f
C1142 input5/a_381_47# output17/a_27_47# 6.6e-20
C1143 p[9] _43_/a_193_413# 1.09e-19
C1144 input10/a_27_47# input12/a_27_47# 0.0154f
C1145 net17 _33_/a_209_311# 7.03e-21
C1146 VPWR _38_/a_109_47# -4.66e-19
C1147 net7 output17/a_27_47# 0.00185f
C1148 _07_ net9 1.39e-20
C1149 _44_/a_93_21# input5/a_664_47# 1.88e-20
C1150 net15 _18_ 0.0382f
C1151 input8/a_27_47# net9 3.71e-20
C1152 _05_ net9 0.124f
C1153 _01_ net11 3.82e-20
C1154 _20_ net2 8.83e-19
C1155 net11 _34_/a_47_47# 0.0309f
C1156 p[9] net2 0.00112f
C1157 _12_ _38_/a_197_47# 0.00173f
C1158 input7/a_27_47# input1/a_75_212# 3.2e-20
C1159 input1/a_75_212# p[13] 4.16e-19
C1160 net14 _55_/a_80_21# 4.7e-19
C1161 VPWR b[2] 0.262f
C1162 VPWR output17/a_27_47# 0.0263f
C1163 net14 _06_ 1.94e-19
C1164 _50_/a_27_47# _22_ 0.0276f
C1165 p[9] p[8] 0.0518f
C1166 _12_ _22_ 0.196f
C1167 input8/a_27_47# input7/a_27_47# 3.2e-20
C1168 net14 net4 2.21e-21
C1169 _19_ _43_/a_193_413# 4.85e-21
C1170 _55_/a_80_21# net1 1.8e-19
C1171 _02_ _38_/a_27_47# 0.00103f
C1172 net14 net5 0.0263f
C1173 input8/a_27_47# _02_ 5.08e-20
C1174 _02_ _07_ 0.0083f
C1175 _02_ _05_ 0.00163f
C1176 _04_ _35_/a_226_297# 4.51e-19
C1177 _18_ _50_/a_343_93# 0.0276f
C1178 net6 _47_/a_299_297# 3.63e-19
C1179 _06_ net1 0.0115f
C1180 p[0] b[1] 0.00123f
C1181 VPWR _30_/a_465_297# -4.57e-19
C1182 _30_/a_392_297# net9 9.92e-19
C1183 _21_ net8 0.00656f
C1184 p[9] p[12] 1.4e-19
C1185 _19_ net2 0.101f
C1186 _10_ net14 2.4e-19
C1187 _45_/a_193_297# _22_ 0.0234f
C1188 net5 net1 0.0772f
C1189 net12 p[7] 0.0343f
C1190 net13 _33_/a_209_311# 0.0227f
C1191 _44_/a_250_297# _15_ 0.00517f
C1192 _01_ _55_/a_472_297# 6.28e-19
C1193 input5/a_558_47# _27_/a_27_297# 1.57e-19
C1194 net6 _06_ 0.308f
C1195 input2/a_27_47# net2 0.024f
C1196 net12 _32_/a_27_47# 1.52e-19
C1197 _34_/a_47_47# _48_/a_27_47# 4.45e-21
C1198 net5 _44_/a_93_21# 3.61e-20
C1199 _36_/a_27_47# _18_ 5.46e-20
C1200 net4 net6 0.713f
C1201 _10_ net1 4.34e-19
C1202 _12_ _50_/a_27_47# 0.00354f
C1203 net5 net6 0.722f
C1204 net12 _04_ 0.267f
C1205 _07_ _35_/a_556_47# 0.00128f
C1206 p[10] _27_/a_27_297# 6.35e-19
C1207 _29_/a_29_53# net10 1.77e-19
C1208 net14 _43_/a_297_47# 1.09e-21
C1209 p[9] output19/a_27_47# 0.0852f
C1210 VPWR _33_/a_368_53# -4.26e-19
C1211 input8/a_27_47# _49_/a_201_297# 2.46e-21
C1212 input5/a_62_47# net14 5.28e-20
C1213 _10_ _44_/a_93_21# 2.48e-19
C1214 _13_ _15_ 3.69e-20
C1215 _01_ _31_/a_285_297# 1.92e-19
C1216 _20_ _55_/a_217_297# 0.0013f
C1217 _35_/a_76_199# _06_ 0.00425f
C1218 _10_ net6 0.0965f
C1219 net15 input5/a_558_47# 0.00672f
C1220 _37_/a_27_47# _42_/a_209_311# 1.59e-20
C1221 _35_/a_76_199# net5 3.38e-19
C1222 _00_ _11_ 0.238f
C1223 _12_ _45_/a_193_297# 0.0103f
C1224 net18 _22_ 1.68e-19
C1225 _15_ net19 0.166f
C1226 input5/a_62_47# net1 7.59e-20
C1227 p[10] net15 0.01f
C1228 _10_ _35_/a_76_199# 7.19e-20
C1229 net6 _43_/a_297_47# 8.23e-22
C1230 _52_/a_93_21# _09_ 0.0227f
C1231 input13/a_27_47# _33_/a_209_311# 5.85e-20
C1232 _27_/a_27_297# _04_ 0.0526f
C1233 input5/a_62_47# _44_/a_93_21# 5.05e-20
C1234 _53_/a_111_297# _22_ 4.7e-20
C1235 _36_/a_109_47# _23_ 3.44e-19
C1236 _03_ net11 0.0952f
C1237 input15/a_27_47# _18_ 8.27e-21
C1238 _03_ _23_ 0.0564f
C1239 _31_/a_35_297# net1 0.0111f
C1240 _55_/a_80_21# _22_ 0.00926f
C1241 VPWR b[0] 0.142f
C1242 _37_/a_197_47# net3 0.0028f
C1243 _38_/a_197_47# _06_ 4.32e-19
C1244 net4 _38_/a_197_47# 7.64e-19
C1245 input14/a_27_47# b[3] 0.0211f
C1246 _20_ _40_/a_297_297# 9.18e-21
C1247 input8/a_27_47# _01_ 1.43e-19
C1248 _03_ _35_/a_226_47# 0.028f
C1249 _01_ _05_ 5.03e-19
C1250 _44_/a_346_47# net19 0.00124f
C1251 _40_/a_109_297# net15 0.0016f
C1252 _37_/a_197_47# _17_ 9.19e-21
C1253 net4 _22_ 0.0866f
C1254 _06_ _22_ 0.124f
C1255 _34_/a_47_47# _07_ 0.011f
C1256 _15_ _50_/a_223_47# 0.00698f
C1257 output18/a_27_47# _54_/a_75_212# 2.28e-19
C1258 _37_/a_27_47# _18_ 3.31e-20
C1259 net15 _04_ 0.0569f
C1260 _34_/a_47_47# _05_ 1.26e-20
C1261 _02_ _42_/a_209_311# 9.92e-19
C1262 _12_ net18 8.24e-19
C1263 net5 _22_ 0.405f
C1264 _35_/a_489_413# _08_ 5.56e-19
C1265 net12 _30_/a_465_297# 8.01e-20
C1266 _10_ _38_/a_197_47# 6.29e-19
C1267 _27_/a_205_297# net3 4.37e-19
C1268 _18_ net9 1.51e-19
C1269 _31_/a_35_297# _49_/a_75_199# 6.24e-19
C1270 b[0] _39_/a_129_47# 2.6e-20
C1271 _41_/a_59_75# net15 1.16e-20
C1272 net14 _44_/a_250_297# 4.24e-20
C1273 _10_ _22_ 0.0904f
C1274 _12_ _47_/a_299_297# 0.00805f
C1275 _30_/a_109_53# _05_ 0.033f
C1276 _32_/a_27_47# _50_/a_343_93# 6.48e-20
C1277 input9/a_75_212# net1 0.002f
C1278 p[2] _31_/a_35_297# 0.00264f
C1279 _34_/a_285_47# VPWR -0.00233f
C1280 net3 _42_/a_209_311# 0.029f
C1281 _39_/a_47_47# net6 0.0249f
C1282 _34_/a_285_47# p[6] 8.31e-20
C1283 _42_/a_296_53# net19 2.71e-19
C1284 net4 _50_/a_27_47# 0.0239f
C1285 _12_ _06_ 0.136f
C1286 _06_ _50_/a_27_47# 0.00972f
C1287 net4 _12_ 0.105f
C1288 net12 _33_/a_368_53# 2.63e-19
C1289 input2/a_27_47# b[1] 8.55e-19
C1290 _42_/a_209_311# _17_ 1.22e-19
C1291 _00_ _43_/a_193_413# 0.00721f
C1292 net5 _50_/a_27_47# 0.0169f
C1293 _44_/a_250_297# _44_/a_93_21# -6.97e-22
C1294 net5 _12_ 0.983f
C1295 net11 p[5] 0.0598f
C1296 _02_ _18_ 2.96e-20
C1297 VPWR _54_/a_75_212# 0.0475f
C1298 net17 net2 0.261f
C1299 _03_ _31_/a_285_297# 0.00677f
C1300 _36_/a_27_47# _32_/a_27_47# 0.011f
C1301 _41_/a_59_75# _50_/a_343_93# 6.13e-22
C1302 _49_/a_208_47# _09_ 5.43e-21
C1303 _10_ _50_/a_27_47# 0.0154f
C1304 _00_ net2 0.00732f
C1305 net14 net19 0.148f
C1306 net4 _45_/a_193_297# 7.41e-19
C1307 _06_ _45_/a_193_297# 0.00201f
C1308 _10_ _12_ 0.19f
C1309 _04_ _36_/a_27_47# 0.00169f
C1310 net11 _29_/a_183_297# 3.64e-19
C1311 _14_ _43_/a_369_47# 0.00135f
C1312 net5 _45_/a_193_297# 0.00935f
C1313 _20_ _29_/a_29_53# 0.0111f
C1314 net14 _27_/a_277_297# 5.1e-19
C1315 net11 net10 0.592f
C1316 _09_ _29_/a_29_53# 0.00488f
C1317 net11 net16 4.43e-22
C1318 _52_/a_93_21# _52_/a_346_47# -5.12e-20
C1319 net10 _23_ 7.53e-19
C1320 _13_ net6 0.0106f
C1321 net3 _18_ 7.34e-20
C1322 _04_ _08_ 5.99e-19
C1323 _10_ _45_/a_193_297# 0.0047f
C1324 _21_ _11_ 9.98e-20
C1325 _44_/a_93_21# net19 0.0074f
C1326 p[2] input9/a_75_212# 5.13e-20
C1327 input5/a_664_47# _06_ 3.21e-19
C1328 _01_ _42_/a_209_311# 1.58e-19
C1329 _17_ _18_ 0.271f
C1330 _35_/a_226_47# net10 0.0159f
C1331 net6 net19 0.00352f
C1332 input14/a_27_47# _11_ 1.42e-19
C1333 _49_/a_208_47# _19_ 7.12e-20
C1334 _03_ _07_ 0.0113f
C1335 net5 input5/a_664_47# 0.0536f
C1336 _03_ _05_ 0.135f
C1337 _35_/a_76_199# _13_ 3.01e-21
C1338 net14 _50_/a_223_47# 5.89e-21
C1339 input5/a_558_47# net9 4.42e-19
C1340 VPWR _32_/a_197_47# 0.00146f
C1341 _34_/a_377_297# _07_ 5.8e-19
C1342 _32_/a_109_47# net9 6.44e-19
C1343 _06_ net18 0.0211f
C1344 _02_ _35_/a_489_413# 3.86e-19
C1345 _14_ _15_ 0.148f
C1346 _26_/a_29_53# _15_ 0.00192f
C1347 VPWR _30_/a_215_297# -0.00472f
C1348 VPWR _32_/a_303_47# 6.03e-19
C1349 _30_/a_215_297# p[3] 2.01e-19
C1350 _53_/a_111_297# _06_ 3.82e-19
C1351 net4 _47_/a_299_297# 3.28e-19
C1352 _47_/a_299_297# _06_ 0.0174f
C1353 input5/a_558_47# input7/a_27_47# 1.22e-20
C1354 _48_/a_27_47# net10 8.4e-21
C1355 input5/a_558_47# p[13] 0.00158f
C1356 _14_ _47_/a_81_21# 6.24e-20
C1357 _53_/a_111_297# net4 2.09e-19
C1358 _41_/a_59_75# input15/a_27_47# 3.96e-20
C1359 net5 _47_/a_299_297# 0.00198f
C1360 _34_/a_285_47# net12 8.07e-20
C1361 net6 _50_/a_223_47# 0.0194f
C1362 _55_/a_80_21# _06_ 5.15e-19
C1363 net4 _55_/a_80_21# 1.06e-19
C1364 _01_ _18_ 6.1e-20
C1365 p[7] net9 8.26e-19
C1366 _03_ _30_/a_392_297# 6.33e-19
C1367 _02_ _32_/a_109_47# 3.98e-19
C1368 net5 _55_/a_80_21# 2.78e-19
C1369 _53_/a_29_53# _11_ 2.33e-20
C1370 output18/a_27_47# _25_ 0.072f
C1371 p[10] p[13] 0.124f
C1372 _14_ _44_/a_346_47# 3.76e-19
C1373 _32_/a_27_47# net9 0.0136f
C1374 _10_ _53_/a_111_297# 2.06e-19
C1375 net4 _06_ 0.281f
C1376 _10_ _47_/a_299_297# 0.0134f
C1377 _02_ p[10] 2.17e-19
C1378 VPWR _43_/a_369_47# -3.75e-19
C1379 _13_ _22_ 0.00309f
C1380 net5 _06_ 0.41f
C1381 _39_/a_47_47# _12_ 0.0317f
C1382 net4 net5 0.0447f
C1383 p[4] p[7] 7.8e-20
C1384 _04_ net9 0.0213f
C1385 _31_/a_285_297# net10 1.68e-19
C1386 _42_/a_109_93# _19_ 1.14e-21
C1387 p[11] _15_ 2.93e-19
C1388 _10_ _55_/a_80_21# 5.49e-19
C1389 _20_ _16_ 0.00271f
C1390 _49_/a_544_297# net7 2.72e-19
C1391 _22_ net19 2.17e-19
C1392 net17 b[1] 0.00766f
C1393 _10_ net4 0.183f
C1394 _10_ _06_ 1.14f
C1395 p[13] _32_/a_27_47# 6.49e-20
C1396 _15_ net7 8.4e-20
C1397 input5/a_558_47# net3 0.0137f
C1398 _10_ net5 0.199f
C1399 _39_/a_47_47# _45_/a_193_297# 1.4e-20
C1400 input5/a_558_47# _17_ 2.13e-21
C1401 _03_ _27_/a_205_297# 1.46e-20
C1402 _02_ _32_/a_27_47# 0.00247f
C1403 net11 input10/a_27_47# 0.112f
C1404 p[10] net3 7.98e-19
C1405 VPWR _49_/a_544_297# 0.00569f
C1406 _02_ _04_ 0.0541f
C1407 _43_/a_297_47# _06_ 4.81e-20
C1408 _13_ _50_/a_27_47# 0.00169f
C1409 VPWR _25_ 0.0829f
C1410 VPWR _15_ 0.912f
C1411 _08_ _33_/a_368_53# 5.04e-19
C1412 net16 _38_/a_27_47# 0.114f
C1413 _13_ _12_ 0.462f
C1414 net10 _07_ 0.057f
C1415 net6 _24_ 0.00121f
C1416 _12_ _38_/a_303_47# 0.00153f
C1417 input14/a_27_47# net2 0.0176f
C1418 VPWR _47_/a_384_47# -1.45e-19
C1419 net13 _52_/a_93_21# 7.21e-19
C1420 net10 _05_ 0.457f
C1421 input5/a_62_47# net5 0.00329f
C1422 _50_/a_223_47# _22_ 0.031f
C1423 _31_/a_35_297# _55_/a_80_21# 5.9e-21
C1424 _21_ input12/a_27_47# 2.32e-19
C1425 VPWR _47_/a_81_21# 0.00889f
C1426 net14 _14_ 0.184f
C1427 _10_ _43_/a_297_47# 0.00118f
C1428 _20_ net11 0.00128f
C1429 _40_/a_109_297# net3 3.14e-19
C1430 input14/a_27_47# p[8] 0.0159f
C1431 net11 _09_ 0.0262f
C1432 _02_ _38_/a_109_47# 1.63e-19
C1433 output16/a_27_47# _38_/a_27_47# 9.02e-19
C1434 _09_ _23_ 0.207f
C1435 _40_/a_109_297# _17_ 9.67e-19
C1436 _45_/a_27_47# net6 0.021f
C1437 net12 _30_/a_215_297# 0.00676f
C1438 net3 _04_ 0.113f
C1439 net14 _26_/a_29_53# 1.33e-20
C1440 _31_/a_35_297# net5 2.04e-21
C1441 VPWR _44_/a_346_47# -8.74e-19
C1442 _01_ input5/a_558_47# 3.97e-20
C1443 _30_/a_465_297# net9 0.00138f
C1444 _20_ _35_/a_226_47# 5.19e-20
C1445 _04_ _17_ 4.34e-19
C1446 p[13] output17/a_27_47# 0.00118f
C1447 _49_/a_201_297# _04_ 0.0253f
C1448 _35_/a_226_47# _09_ 0.058f
C1449 _01_ _32_/a_109_47# 0.00129f
C1450 _45_/a_27_47# _35_/a_76_199# 2.04e-21
C1451 _14_ _44_/a_93_21# 0.04f
C1452 _02_ b[2] 2.69e-19
C1453 p[10] _01_ 7.94e-20
C1454 _30_/a_392_297# net10 3.4e-19
C1455 _03_ _18_ 7.25e-23
C1456 _14_ net6 2.11e-19
C1457 _41_/a_59_75# _17_ 0.00149f
C1458 p[0] input1/a_75_212# 0.0172f
C1459 _49_/a_75_199# _49_/a_315_47# 1.78e-33
C1460 _50_/a_27_47# _50_/a_223_47# 5.68e-32
C1461 _12_ _50_/a_223_47# 0.00327f
C1462 net11 _19_ 6.27e-21
C1463 _11_ _43_/a_27_47# 4.27e-19
C1464 _43_/a_469_47# _18_ 1.59e-19
C1465 _26_/a_29_53# net6 0.0032f
C1466 _39_/a_47_47# _06_ 1.44e-19
C1467 input5/a_664_47# net19 1.38e-21
C1468 input14/a_27_47# output19/a_27_47# 0.0101f
C1469 net4 _39_/a_47_47# 0.0202f
C1470 p[2] _49_/a_315_47# 6.65e-20
C1471 _01_ _31_/a_285_47# 3.36e-19
C1472 net14 p[11] 0.00182f
C1473 _28_/a_109_297# _15_ 0.00346f
C1474 input5/a_381_47# net14 0.00479f
C1475 net5 _39_/a_47_47# 0.0352f
C1476 _09_ _48_/a_27_47# 0.00541f
C1477 _49_/a_75_199# _14_ 6.79e-20
C1478 _20_ _55_/a_472_297# 0.00212f
C1479 _24_ _22_ 0.0846f
C1480 _01_ _32_/a_27_47# 0.0266f
C1481 net14 net7 2.23e-19
C1482 VPWR _42_/a_296_53# -6.37e-20
C1483 p[12] _52_/a_250_297# 1.84e-20
C1484 net3 output17/a_27_47# 0.00248f
C1485 _52_/a_93_21# _33_/a_109_93# 2.89e-21
C1486 net10 _33_/a_296_53# 8.22e-20
C1487 net5 _44_/a_250_297# 3.11e-20
C1488 input5/a_381_47# net1 1.27e-19
C1489 _01_ _04_ 0.119f
C1490 _10_ _39_/a_47_47# 0.00824f
C1491 _04_ _34_/a_47_47# 1.17e-20
C1492 _34_/a_285_47# _08_ 0.00414f
C1493 _52_/a_93_21# _21_ 9.4e-19
C1494 _27_/a_109_297# _04_ 7.2e-20
C1495 net7 net1 0.0712f
C1496 net12 _25_ 4.46e-20
C1497 _45_/a_27_47# _22_ 0.0131f
C1498 _53_/a_183_297# _22_ 3.71e-20
C1499 VPWR net14 0.182f
C1500 net17 _42_/a_109_93# 3.1e-21
C1501 _10_ input9/a_75_212# 5.49e-21
C1502 _34_/a_129_47# net11 0.00242f
C1503 _13_ _06_ 0.00188f
C1504 net4 _13_ 0.212f
C1505 _30_/a_109_53# _32_/a_27_47# 1.51e-19
C1506 _55_/a_80_21# net19 0.00423f
C1507 net4 _38_/a_303_47# 5.95e-19
C1508 _11_ net8 1.81e-20
C1509 net13 _29_/a_29_53# 0.00104f
C1510 _03_ _35_/a_489_413# 0.0205f
C1511 net5 _13_ 0.0352f
C1512 _30_/a_109_53# _04_ 9.19e-21
C1513 VPWR net1 1.17f
C1514 _12_ _24_ 1.67e-19
C1515 p[3] net1 6.54e-19
C1516 p[6] net1 3.12e-20
C1517 net4 net19 2.65e-20
C1518 _06_ net19 0.00522f
C1519 net5 net19 0.00124f
C1520 _14_ _22_ 0.00449f
C1521 net14 _37_/a_303_47# 0.00112f
C1522 p[1] net2 5.99e-20
C1523 VPWR _44_/a_93_21# 0.005f
C1524 net14 _42_/a_368_53# 7.39e-19
C1525 _26_/a_29_53# _22_ 0.09f
C1526 _10_ _13_ 0.0621f
C1527 _49_/a_75_199# net7 0.09f
C1528 _35_/a_76_199# net7 1.79e-20
C1529 input5/a_62_47# _44_/a_250_297# 2.45e-20
C1530 _10_ _38_/a_303_47# 7.36e-19
C1531 VPWR net6 0.999f
C1532 _31_/a_285_297# _19_ 1.34e-19
C1533 _27_/a_27_297# _15_ 9.85e-20
C1534 _52_/a_93_21# _52_/a_250_297# -6.97e-22
C1535 _45_/a_27_47# _12_ 0.0866f
C1536 _45_/a_27_47# _50_/a_27_47# 0.109f
C1537 _20_ _07_ 1.28e-21
C1538 _47_/a_299_297# _50_/a_223_47# 2.74e-20
C1539 b[0] _39_/a_285_47# 1.88e-19
C1540 _10_ net19 0.00224f
C1541 _09_ _07_ 0.0405f
C1542 _20_ _05_ 6.79e-19
C1543 net14 _44_/a_256_47# 0.00379f
C1544 _26_/a_111_297# net6 1.12e-19
C1545 _09_ _38_/a_27_47# 0.00195f
C1546 p[2] net7 0.00156f
C1547 _09_ _05_ 0.0683f
C1548 _52_/a_93_21# _53_/a_29_53# 0.00116f
C1549 _00_ _16_ 0.00613f
C1550 VPWR _49_/a_75_199# 0.0177f
C1551 _35_/a_76_199# VPWR -0.00947f
C1552 output18/a_27_47# _22_ 7.51e-19
C1553 input4/a_75_212# _18_ 4.36e-19
C1554 _30_/a_215_297# _36_/a_27_47# 7.13e-20
C1555 _03_ p[10] 8.74e-20
C1556 net10 _18_ 1.47e-21
C1557 net16 _18_ 8.17e-21
C1558 _39_/a_377_297# net6 0.00143f
C1559 _06_ _50_/a_223_47# 0.0481f
C1560 net4 _50_/a_223_47# 0.0107f
C1561 _43_/a_27_47# net2 0.01f
C1562 net15 _15_ 0.156f
C1563 _14_ _12_ 1.98e-20
C1564 _39_/a_129_47# net6 6.91e-19
C1565 net5 _50_/a_223_47# 0.00202f
C1566 p[2] VPWR 0.103f
C1567 p[2] p[3] 0.188f
C1568 _44_/a_256_47# _44_/a_93_21# -6.6e-20
C1569 p[11] _22_ 3.13e-20
C1570 _26_/a_29_53# _50_/a_27_47# 5.56e-19
C1571 _26_/a_29_53# _12_ 0.00243f
C1572 _03_ _31_/a_285_47# 8.54e-19
C1573 b[3] p[14] 0.0645f
C1574 b[3] _11_ 2.37e-20
C1575 _03_ _32_/a_27_47# 1.9e-19
C1576 net7 _22_ 2.73e-20
C1577 net18 _24_ 5.57e-21
C1578 net15 _47_/a_81_21# 0.00106f
C1579 _10_ _50_/a_223_47# 0.0295f
C1580 _04_ _36_/a_109_47# 2.39e-19
C1581 _03_ _04_ 0.586f
C1582 _11_ _40_/a_191_297# 0.00207f
C1583 _34_/a_285_47# _02_ 7.14e-19
C1584 VPWR _38_/a_197_47# -5.24e-19
C1585 _21_ _29_/a_29_53# 0.0775f
C1586 input2/a_27_47# _05_ 1.83e-19
C1587 net11 net17 3.19e-20
C1588 _34_/a_377_297# _04_ 1.7e-20
C1589 _43_/a_193_413# net8 1.62e-20
C1590 _15_ _50_/a_343_93# 0.0098f
C1591 _53_/a_111_297# _24_ 9.08e-21
C1592 VPWR _22_ 1.4f
C1593 _02_ _54_/a_75_212# 6.6e-20
C1594 _26_/a_111_297# _22_ 0.00137f
C1595 net12 net1 1.17e-19
C1596 net2 net8 0.0525f
C1597 _39_/a_47_47# _13_ 0.00117f
C1598 _47_/a_81_21# _50_/a_343_93# 0.00282f
C1599 net4 _24_ 8.65e-20
C1600 _06_ _24_ 0.113f
C1601 net5 _24_ 5.83e-20
C1602 _25_ _36_/a_27_47# 2.34e-20
C1603 net12 net6 0.00643f
C1604 _32_/a_197_47# net9 6.06e-19
C1605 _43_/a_27_47# _55_/a_217_297# 2.18e-19
C1606 net14 _27_/a_27_297# 0.0118f
C1607 _20_ _42_/a_209_311# 1.66e-20
C1608 _26_/a_29_53# net18 2.57e-21
C1609 _03_ output17/a_27_47# 1.95e-19
C1610 p[9] _42_/a_209_311# 5.51e-21
C1611 _45_/a_27_47# net4 0.024f
C1612 _45_/a_27_47# _06_ 0.0021f
C1613 _10_ _24_ 0.00484f
C1614 _44_/a_250_297# net19 0.00592f
C1615 p[5] p[7] 6.77e-20
C1616 _30_/a_215_297# net9 0.0458f
C1617 _32_/a_303_47# net9 0.00218f
C1618 _53_/a_183_297# _06_ 0.00146f
C1619 VPWR _50_/a_27_47# -0.00335f
C1620 _45_/a_27_47# net5 0.0288f
C1621 VPWR _12_ 0.28f
C1622 _35_/a_76_199# net12 0.0132f
C1623 net13 net11 0.093f
C1624 _27_/a_27_297# net1 6.05e-21
C1625 _21_ input5/a_841_47# 1.59e-21
C1626 net13 _23_ 4.11e-19
C1627 _02_ _32_/a_197_47# 3.78e-19
C1628 _14_ _55_/a_80_21# 0.0175f
C1629 _03_ _30_/a_465_297# 7.72e-19
C1630 output18/a_27_47# net18 0.0106f
C1631 _45_/a_27_47# _10_ 0.0143f
C1632 net13 _35_/a_226_47# 0.00709f
C1633 net14 net15 1.07f
C1634 input6/a_27_47# _15_ 5.75e-19
C1635 net4 _14_ 1.54e-20
C1636 _10_ _53_/a_183_297# 2.86e-19
C1637 VPWR _45_/a_193_297# -0.00859f
C1638 input15/a_27_47# _15_ 2.15e-20
C1639 _14_ _06_ 0.0556f
C1640 net5 _14_ 3.89e-19
C1641 _39_/a_377_297# _12_ 6.77e-19
C1642 _02_ _30_/a_215_297# 3.58e-21
C1643 net10 p[7] 4.96e-19
C1644 _02_ _32_/a_303_47# 1.15e-20
C1645 input5/a_664_47# net7 0.00199f
C1646 _39_/a_129_47# _12_ 0.00175f
C1647 net15 net1 7.44e-20
C1648 net11 _36_/a_303_47# 7.63e-20
C1649 net4 _26_/a_29_53# 0.00412f
C1650 _26_/a_29_53# _06_ 0.0135f
C1651 net10 _32_/a_27_47# 2.76e-20
C1652 _04_ _29_/a_183_297# 0.0015f
C1653 net5 _26_/a_29_53# 0.0237f
C1654 b[3] net2 0.311f
C1655 _49_/a_75_199# _27_/a_27_297# 0.011f
C1656 _20_ _18_ 0.0151f
C1657 _06_ _29_/a_111_297# 6.74e-20
C1658 _04_ net10 0.121f
C1659 _10_ _14_ 0.0571f
C1660 input2/a_27_47# _42_/a_209_311# 1e-22
C1661 _09_ _18_ 7.01e-21
C1662 net15 _44_/a_93_21# 0.00573f
C1663 input14/a_27_47# input3/a_27_47# 5.08e-20
C1664 _40_/a_191_297# net2 0.00143f
C1665 _37_/a_27_47# _15_ 1.11e-19
C1666 VPWR input5/a_664_47# 0.00488f
C1667 _10_ _26_/a_29_53# 0.0265f
C1668 net12 _22_ 5.73e-20
C1669 output18/a_27_47# _06_ 0.0114f
C1670 net15 net6 0.0664f
C1671 b[3] p[8] 0.226f
C1672 VPWR input11/a_27_47# 0.0375f
C1673 net14 _50_/a_343_93# 1.07e-20
C1674 _41_/a_59_75# input4/a_75_212# 0.00153f
C1675 p[0] p[10] 8.21e-20
C1676 _14_ _43_/a_297_47# 9.11e-19
C1677 _15_ net9 0.00113f
C1678 _13_ _50_/a_223_47# 8.2e-20
C1679 _12_ _35_/a_226_297# 3.35e-20
C1680 VPWR net18 0.104f
C1681 net16 _38_/a_109_47# 4.17e-19
C1682 _49_/a_75_199# net15 5.13e-20
C1683 net17 _05_ 0.0111f
C1684 input13/a_27_47# _35_/a_226_47# 3.94e-20
C1685 input5/a_381_47# _06_ 1.6e-19
C1686 _55_/a_80_21# net7 0.00163f
C1687 b[3] p[12] 7.54e-20
C1688 net11 _33_/a_109_93# 5.14e-19
C1689 input5/a_381_47# net5 0.0546f
C1690 net13 _31_/a_285_297# 3.85e-20
C1691 _00_ _05_ 5.03e-22
C1692 b[1] net8 0.00195f
C1693 _06_ net7 0.00447f
C1694 _53_/a_111_297# VPWR 1.11e-34
C1695 VPWR _47_/a_299_297# 0.0643f
C1696 _21_ net11 0.586f
C1697 _47_/a_81_21# net9 3.49e-19
C1698 net6 _50_/a_343_93# 0.00214f
C1699 net5 net7 0.195f
C1700 _21_ _23_ 0.0217f
C1701 _10_ _41_/a_145_75# 5.18e-19
C1702 _45_/a_109_297# net6 7.82e-19
C1703 VPWR _55_/a_80_21# 0.0289f
C1704 net10 output17/a_27_47# 1.31e-20
C1705 _35_/a_226_47# _33_/a_109_93# 4.9e-19
C1706 net12 _12_ 7.94e-21
C1707 net12 _50_/a_27_47# 7.99e-21
C1708 _36_/a_27_47# net1 6.99e-20
C1709 _21_ _35_/a_226_47# 9.87e-19
C1710 _02_ _15_ 0.101f
C1711 _02_ _25_ 0.0156f
C1712 _43_/a_369_47# _17_ 5.87e-19
C1713 _01_ _32_/a_197_47# 0.00156f
C1714 output19/a_27_47# b[3] 0.00809f
C1715 VPWR _06_ 1.4f
C1716 VPWR net4 1.07f
C1717 _06_ p[3] 1.59e-20
C1718 p[6] _06_ 2.62e-19
C1719 _10_ net7 6.22e-20
C1720 _35_/a_489_413# _09_ 0.0296f
C1721 _45_/a_27_47# _39_/a_47_47# 1.31e-19
C1722 VPWR net5 0.612f
C1723 b[3] _55_/a_217_297# 3.41e-19
C1724 net6 _36_/a_27_47# 5.1e-19
C1725 _26_/a_111_297# _06_ 9e-19
C1726 _30_/a_465_297# net10 0.00106f
C1727 _02_ _47_/a_81_21# 1.59e-20
C1728 net15 _22_ 2.74e-19
C1729 _01_ _32_/a_303_47# 8.58e-19
C1730 net13 _07_ 0.00686f
C1731 net14 input6/a_27_47# 7.05e-19
C1732 net13 _05_ 0.192f
C1733 input5/a_62_47# p[11] 0.00153f
C1734 _10_ p[3] 1.37e-20
C1735 _11_ _43_/a_193_413# 5.45e-19
C1736 _13_ _24_ 2.47e-19
C1737 _10_ VPWR 0.577f
C1738 net11 _52_/a_250_297# 1.2e-19
C1739 _39_/a_377_297# _06_ 8.76e-20
C1740 net4 _39_/a_377_297# 8.88e-19
C1741 _35_/a_76_199# _36_/a_27_47# 3.22e-19
C1742 _10_ _26_/a_111_297# 7.13e-20
C1743 _52_/a_250_297# _23_ 3.17e-19
C1744 net3 _15_ 0.224f
C1745 input5/a_62_47# net7 2.04e-19
C1746 _21_ _48_/a_27_47# 0.0121f
C1747 net2 p[14] 1.38e-19
C1748 net5 _39_/a_377_297# 0.00234f
C1749 net5 _39_/a_129_47# 0.00344f
C1750 net11 _53_/a_29_53# 8.31e-19
C1751 _15_ _17_ 0.0752f
C1752 _11_ net2 0.234f
C1753 _35_/a_226_47# _52_/a_250_297# 2.63e-20
C1754 _14_ _44_/a_250_297# 4.82e-19
C1755 VPWR _43_/a_297_47# -2.11e-19
C1756 _45_/a_27_47# _13_ 0.0703f
C1757 _49_/a_208_47# net8 1.4e-19
C1758 net10 _33_/a_368_53# 0.00171f
C1759 _47_/a_384_47# _17_ 1.1e-20
C1760 net3 _47_/a_81_21# 6.66e-19
C1761 net14 _37_/a_27_47# 0.0584f
C1762 p[0] output17/a_27_47# 0.00805f
C1763 _35_/a_76_199# _08_ 0.0061f
C1764 _03_ _54_/a_75_212# 5.45e-21
C1765 b[3] b[1] 6.12e-20
C1766 _10_ _39_/a_377_297# 7.42e-19
C1767 _44_/a_93_21# input6/a_27_47# 8.53e-19
C1768 p[14] p[8] 0.226f
C1769 _31_/a_35_297# net7 0.0384f
C1770 input5/a_62_47# VPWR 0.0601f
C1771 _10_ _39_/a_129_47# 2.51e-19
C1772 input6/a_27_47# net6 0.00208f
C1773 _11_ p[8] 7.7e-20
C1774 _50_/a_343_93# _22_ 0.0597f
C1775 _45_/a_109_297# _22_ 0.0425f
C1776 _47_/a_81_21# _17_ 0.0456f
C1777 net6 input15/a_27_47# 0.146f
C1778 net15 _12_ 8.14e-21
C1779 _09_ p[7] 9.25e-21
C1780 net3 _44_/a_346_47# 8.04e-19
C1781 _55_/a_80_21# _28_/a_109_297# 2.05e-20
C1782 _20_ _40_/a_109_297# 2.35e-20
C1783 net17 _42_/a_209_311# 1.04e-21
C1784 net14 net9 7.12e-20
C1785 _06_ _35_/a_226_297# 1.28e-19
C1786 net13 _30_/a_392_297# 6.64e-20
C1787 _20_ _32_/a_27_47# 0.0069f
C1788 _14_ _13_ 1.47e-20
C1789 _44_/a_346_47# _17_ 7.2e-19
C1790 p[12] p[14] 0.00101f
C1791 VPWR _31_/a_35_297# 0.0333f
C1792 _20_ _04_ 0.0677f
C1793 p[12] _11_ 3.51e-21
C1794 input2/a_27_47# input5/a_558_47# 2.04e-20
C1795 input13/a_27_47# _05_ 3.93e-19
C1796 _04_ _09_ 0.0904f
C1797 _37_/a_27_47# _44_/a_93_21# 3.19e-19
C1798 p[10] _19_ 0.00226f
C1799 _01_ _49_/a_544_297# 0.00109f
C1800 _36_/a_27_47# _22_ 2.82e-20
C1801 net9 net1 0.47f
C1802 _37_/a_27_47# net6 4.3e-20
C1803 input5/a_664_47# _27_/a_27_297# 0.0116f
C1804 _14_ net19 0.00714f
C1805 net14 p[13] 1.91e-19
C1806 _01_ _15_ 0.007f
C1807 _53_/a_29_53# _48_/a_27_47# 3.14e-21
C1808 net14 input7/a_27_47# 3.48e-19
C1809 p[9] _41_/a_59_75# 1.02e-19
C1810 _20_ _41_/a_59_75# 1.78e-20
C1811 b[0] net16 0.0306f
C1812 p[10] input2/a_27_47# 0.00924f
C1813 _34_/a_47_47# _25_ 1.08e-19
C1814 _44_/a_250_297# p[11] 1.13e-19
C1815 _16_ _43_/a_27_47# 2.47e-19
C1816 _10_ _28_/a_109_297# 4.34e-19
C1817 _07_ _33_/a_109_93# 3.2e-19
C1818 _02_ net14 0.00952f
C1819 net4 net12 2.57e-20
C1820 net12 _06_ 0.284f
C1821 _52_/a_93_21# _52_/a_256_47# -6.6e-20
C1822 output19/a_27_47# p[14] 0.0932f
C1823 _12_ _50_/a_343_93# 5.63e-20
C1824 net13 _33_/a_296_53# 3.71e-20
C1825 _05_ _33_/a_109_93# 0.0206f
C1826 _45_/a_109_297# _12_ 0.00587f
C1827 _21_ _38_/a_27_47# 3.87e-19
C1828 input7/a_27_47# net1 0.0383f
C1829 p[13] net1 2.13e-19
C1830 _21_ _07_ 0.133f
C1831 net5 net12 0.0674f
C1832 _01_ _47_/a_81_21# 6.05e-21
C1833 _21_ _05_ 0.0104f
C1834 net15 input5/a_664_47# 0.0216f
C1835 _42_/a_296_53# net3 1.81e-19
C1836 b[0] output16/a_27_47# 0.014f
C1837 VPWR _39_/a_47_47# 0.0668f
C1838 _04_ _19_ 0.356f
C1839 _02_ net1 0.00251f
C1840 _49_/a_75_199# net9 0.00382f
C1841 input5/a_841_47# net8 0.025f
C1842 net14 _44_/a_584_47# 7.2e-19
C1843 _50_/a_27_47# _36_/a_27_47# 6.08e-19
C1844 _10_ net12 0.00257f
C1845 _00_ _18_ 0.157f
C1846 _03_ _30_/a_215_297# 0.0393f
C1847 _12_ _36_/a_27_47# 0.00178f
C1848 net6 _45_/a_465_47# 6.06e-20
C1849 _09_ b[2] 4.28e-20
C1850 input9/a_75_212# p[3] 0.0157f
C1851 VPWR input9/a_75_212# 0.0641f
C1852 input2/a_27_47# _04_ 4.5e-21
C1853 VPWR _44_/a_250_297# 0.0231f
C1854 _39_/a_285_47# net6 1.53e-19
C1855 _43_/a_193_413# net2 1.52e-19
C1856 net14 net3 0.689f
C1857 _02_ net6 0.00427f
C1858 p[2] net9 1.4e-20
C1859 p[11] net19 0.00646f
C1860 input5/a_381_47# net19 0.00173f
C1861 _26_/a_29_53# _50_/a_223_47# 0.00124f
C1862 net14 _49_/a_201_297# 1.52e-19
C1863 net5 _27_/a_27_297# 3.48e-19
C1864 _34_/a_285_47# net10 0.0454f
C1865 net14 _17_ 0.104f
C1866 net15 _47_/a_299_297# 1.44e-20
C1867 net3 net1 4.25e-20
C1868 _16_ net8 0.00624f
C1869 _52_/a_250_297# _05_ 8.86e-22
C1870 _02_ _49_/a_75_199# 0.0354f
C1871 net16 _54_/a_75_212# 1.69e-21
C1872 _54_/a_75_212# net10 6.24e-19
C1873 _02_ _35_/a_76_199# 5.73e-19
C1874 _53_/a_29_53# _38_/a_27_47# 1.29e-19
C1875 _11_ _40_/a_297_297# 9.94e-19
C1876 VPWR _13_ 0.0804f
C1877 p[2] input7/a_27_47# 0.0023f
C1878 _49_/a_201_297# net1 0.00304f
C1879 VPWR _38_/a_303_47# -4.83e-19
C1880 net2 p[8] 0.00102f
C1881 net15 _55_/a_80_21# 0.00759f
C1882 _45_/a_27_47# _24_ 4.57e-19
C1883 _44_/a_93_21# net3 0.0102f
C1884 _15_ _50_/a_429_93# 6.82e-19
C1885 net3 net6 0.00152f
C1886 _02_ p[2] 7.08e-19
C1887 _19_ output17/a_27_47# 7.69e-19
C1888 _44_/a_93_21# _17_ 0.0646f
C1889 net4 net15 8.68e-19
C1890 net9 _22_ 0.0023f
C1891 VPWR net19 0.181f
C1892 net15 _06_ 0.033f
C1893 net13 _18_ 1.06e-20
C1894 net5 net15 0.0226f
C1895 net6 _17_ 3.12e-19
C1896 b[3] _42_/a_109_93# 3.29e-19
C1897 input2/a_27_47# output17/a_27_47# 0.107f
C1898 VPWR _27_/a_277_297# -3.63e-19
C1899 _49_/a_75_199# net3 2.01e-19
C1900 net14 _01_ 8.29e-19
C1901 _03_ _49_/a_544_297# 0.00568f
C1902 _25_ _36_/a_109_47# 3.76e-21
C1903 _10_ net15 0.0101f
C1904 _03_ _15_ 7.39e-20
C1905 _03_ _25_ 0.00422f
C1906 _42_/a_368_53# net19 5.12e-19
C1907 _26_/a_29_53# _24_ 2.11e-20
C1908 net14 _27_/a_109_297# 1.32e-19
C1909 input5/a_558_47# net17 2.88e-21
C1910 net11 net8 1.5e-19
C1911 _02_ _22_ 0.552f
C1912 _01_ net1 0.0509f
C1913 net4 _50_/a_343_93# 0.00124f
C1914 _45_/a_109_297# _06_ 0.0023f
C1915 output19/a_27_47# net2 0.00168f
C1916 _06_ _50_/a_343_93# 0.0376f
C1917 _45_/a_109_297# net4 6.43e-20
C1918 net5 _50_/a_343_93# 0.00124f
C1919 VPWR _50_/a_223_47# -0.00601f
C1920 p[2] _49_/a_201_297# 4.58e-20
C1921 _12_ net9 4.39e-22
C1922 _45_/a_109_297# net5 0.0184f
C1923 p[10] net17 0.18f
C1924 _16_ b[3] 2.9e-19
C1925 output19/a_27_47# p[8] 0.0218f
C1926 _30_/a_215_297# net10 0.0512f
C1927 b[3] input3/a_27_47# 0.012f
C1928 _10_ _50_/a_343_93# 0.0284f
C1929 input1/a_75_212# p[1] 0.0023f
C1930 net13 _35_/a_489_413# 7.36e-20
C1931 _06_ _36_/a_27_47# 0.0501f
C1932 net4 _36_/a_27_47# 0.0103f
C1933 _45_/a_109_297# _10_ 0.00202f
C1934 input8/a_27_47# p[1] 5.13e-20
C1935 _30_/a_109_53# net1 0.0297f
C1936 net3 _22_ 9.39e-20
C1937 _12_ _45_/a_465_47# 0.00211f
C1938 net5 _36_/a_27_47# 0.0163f
C1939 _31_/a_285_47# net17 0.00134f
C1940 _35_/a_76_199# _01_ 3.08e-21
C1941 _01_ _49_/a_75_199# 0.009f
C1942 _02_ _50_/a_27_47# 2.09e-19
C1943 _17_ _22_ 0.00334f
C1944 _39_/a_285_47# _12_ 0.0221f
C1945 output19/a_27_47# p[12] 1.78e-19
C1946 _14_ _26_/a_29_53# 3.67e-19
C1947 _49_/a_201_297# _22_ 2.45e-20
C1948 _02_ _12_ 0.265f
C1949 _06_ _08_ 0.0343f
C1950 _04_ net17 0.0218f
C1951 _10_ _36_/a_27_47# 0.00109f
C1952 _00_ _32_/a_27_47# 0.00228f
C1953 p[2] _01_ 0.00164f
C1954 input10/a_27_47# _54_/a_75_212# 1.17e-22
C1955 b[1] net2 0.0191f
C1956 _00_ _04_ 1.98e-20
C1957 _40_/a_297_297# net2 0.00101f
C1958 input5/a_664_47# net9 5.29e-19
C1959 net14 _50_/a_429_93# 6.04e-21
C1960 VPWR _24_ 0.0129f
C1961 _02_ _45_/a_193_297# 0.00988f
C1962 _10_ _08_ 1.51e-19
C1963 input6/a_27_47# _06_ 2.85e-19
C1964 _41_/a_59_75# _00_ 2.43e-20
C1965 input15/a_27_47# _06_ 4.73e-19
C1966 _31_/a_285_297# net8 0.0215f
C1967 _49_/a_315_47# net7 0.00706f
C1968 net3 _12_ 3.09e-20
C1969 _39_/a_47_47# net15 9.44e-22
C1970 p[4] input11/a_27_47# 0.0646f
C1971 input5/a_664_47# input7/a_27_47# 1.08e-21
C1972 input5/a_664_47# p[13] 8.06e-19
C1973 _14_ p[11] 7.85e-20
C1974 input5/a_381_47# _14_ 5.68e-20
C1975 _50_/a_27_47# _17_ 3.93e-20
C1976 _12_ _17_ 0.0109f
C1977 net13 p[7] 0.00809f
C1978 net11 _33_/a_209_311# 2.49e-19
C1979 net15 _44_/a_250_297# 8.86e-20
C1980 _01_ _22_ 0.15f
C1981 _45_/a_27_47# VPWR -0.00418f
C1982 net16 _25_ 1.16e-19
C1983 _03_ net14 1.5e-19
C1984 _02_ input5/a_664_47# 0.00187f
C1985 _14_ net7 0.00251f
C1986 _52_/a_250_297# _18_ 1.77e-19
C1987 _25_ net10 2.02e-19
C1988 _10_ input15/a_27_47# 4.5e-19
C1989 _10_ input6/a_27_47# 4.57e-20
C1990 VPWR _49_/a_315_47# 6.26e-19
C1991 net11 _48_/a_109_47# 1.74e-19
C1992 _34_/a_47_47# _22_ 3.9e-21
C1993 net6 _50_/a_429_93# 6.18e-19
C1994 _37_/a_27_47# _06_ 2.5e-20
C1995 _27_/a_27_297# net19 1.98e-19
C1996 net14 _43_/a_469_47# 1.44e-20
C1997 net17 output17/a_27_47# 0.0149f
C1998 net13 _04_ 0.569f
C1999 _35_/a_226_47# _33_/a_209_311# 1.31e-19
C2000 _37_/a_27_47# net5 1.13e-20
C2001 _03_ net1 0.298f
C2002 _21_ _35_/a_489_413# 0.0448f
C2003 _02_ net18 6.8e-20
C2004 _06_ net9 0.0505f
C2005 net4 net9 1.99e-22
C2006 VPWR _14_ 0.186f
C2007 input8/a_27_47# net8 0.0181f
C2008 _30_/a_109_53# _22_ 3.67e-21
C2009 net8 _05_ 0.0146f
C2010 _16_ _11_ 4.42e-20
C2011 net5 net9 0.0368f
C2012 b[3] _55_/a_472_297# 1.51e-19
C2013 _03_ net6 2.9e-20
C2014 VPWR _26_/a_29_53# 0.0356f
C2015 input5/a_664_47# net3 0.00215f
C2016 _53_/a_111_297# _02_ 9.57e-20
C2017 net15 net19 0.0501f
C2018 VPWR _29_/a_111_297# -5.85e-19
C2019 _43_/a_469_47# net6 4.85e-21
C2020 _10_ net9 0.0438f
C2021 _02_ _55_/a_80_21# 0.164f
C2022 input13/a_27_47# p[7] 0.0167f
C2023 input5/a_381_47# net7 4.91e-19
C2024 _27_/a_277_297# net15 1.93e-19
C2025 _03_ _49_/a_75_199# 0.0849f
C2026 net5 p[13] 0.0069f
C2027 _39_/a_285_47# _06_ 1.23e-20
C2028 _52_/a_256_47# _23_ 6.66e-19
C2029 net4 _39_/a_285_47# 9.71e-19
C2030 _03_ _35_/a_76_199# 0.0733f
C2031 _02_ net4 0.00376f
C2032 VPWR output18/a_27_47# 0.0689f
C2033 _02_ _06_ 0.85f
C2034 net5 _39_/a_285_47# 0.0405f
C2035 _26_/a_183_297# _15_ 4.63e-36
C2036 _13_ _50_/a_343_93# 5.63e-20
C2037 _02_ net5 0.233f
C2038 _20_ _30_/a_215_297# 6.08e-19
C2039 _14_ _44_/a_256_47# 0.00124f
C2040 _20_ _32_/a_303_47# 1.54e-19
C2041 _30_/a_297_297# _30_/a_215_297# -8.88e-34
C2042 _10_ _45_/a_465_47# 3.32e-19
C2043 net3 _47_/a_299_297# 2.55e-19
C2044 _41_/a_145_75# VPWR -2.46e-19
C2045 _31_/a_117_297# net7 0.00472f
C2046 VPWR p[11] 0.247f
C2047 p[7] _33_/a_109_93# 1.15e-19
C2048 input5/a_381_47# VPWR 8.33e-19
C2049 input5/a_62_47# net9 3.12e-19
C2050 _10_ _39_/a_285_47# 0.00289f
C2051 _36_/a_197_47# _25_ 2.37e-21
C2052 _10_ _02_ 0.0537f
C2053 net3 _55_/a_80_21# 2.35e-19
C2054 _11_ _23_ 2e-20
C2055 net13 _30_/a_465_297# 6.36e-20
C2056 VPWR net7 0.784f
C2057 net4 net3 9.28e-21
C2058 _21_ _32_/a_27_47# 8.95e-19
C2059 _04_ _33_/a_109_93# 0.0299f
C2060 _55_/a_80_21# _17_ 7.64e-21
C2061 net3 _06_ 0.0072f
C2062 VPWR _31_/a_117_297# 8.41e-19
C2063 _42_/a_109_93# net2 0.00507f
C2064 _21_ _04_ 0.39f
C2065 _14_ _28_/a_109_297# 5.66e-19
C2066 net6 _45_/a_205_47# 2.59e-20
C2067 net5 net3 0.0365f
C2068 _06_ _17_ 0.0341f
C2069 net4 _17_ 7.52e-21
C2070 input5/a_62_47# p[13] 0.0202f
C2071 _37_/a_303_47# p[11] 1.04e-19
C2072 _10_ _44_/a_584_47# 1.14e-20
C2073 _03_ _22_ 2.55e-20
C2074 net5 _17_ 0.00408f
C2075 input10/a_27_47# _25_ 2.03e-20
C2076 VPWR p[3] 0.0874f
C2077 VPWR p[6] 0.0738f
C2078 VPWR _26_/a_111_297# -5.92e-20
C2079 _10_ net3 3.89e-19
C2080 net10 net1 0.00388f
C2081 _16_ _43_/a_193_413# 0.0261f
C2082 input2/a_27_47# _30_/a_215_297# 3.51e-20
C2083 net13 _33_/a_368_53# 2.1e-20
C2084 _05_ _33_/a_209_311# 0.0311f
C2085 _07_ _33_/a_209_311# 0.00859f
C2086 _10_ _17_ 0.0233f
C2087 _43_/a_27_47# _18_ 0.0201f
C2088 _48_/a_109_47# _07_ 3.01e-19
C2089 _02_ _31_/a_35_297# 0.00316f
C2090 _42_/a_209_311# net8 7.7e-21
C2091 net12 _26_/a_29_53# 6.55e-19
C2092 _49_/a_544_297# _09_ 2.56e-20
C2093 _16_ net2 0.00654f
C2094 _20_ _15_ 0.691f
C2095 VPWR _37_/a_303_47# -3.13e-19
C2096 VPWR _42_/a_368_53# -3.03e-19
C2097 _01_ _55_/a_80_21# 0.0121f
C2098 p[9] _15_ 2.06e-19
C2099 input4/a_75_212# net6 0.0273f
C2100 VPWR _39_/a_129_47# -9.47e-19
C2101 net6 net10 1.35e-20
C2102 net6 net16 8.27e-20
C2103 _09_ _25_ 1.49e-19
C2104 _04_ _52_/a_250_297# 3.98e-21
C2105 net12 _29_/a_111_297# 1.21e-19
C2106 input3/a_27_47# net2 0.0222f
C2107 _50_/a_223_47# _36_/a_27_47# 1.27e-20
C2108 input5/a_62_47# net3 0.00164f
C2109 _43_/a_297_47# _17_ 5.72e-20
C2110 _20_ _47_/a_384_47# 1.72e-19
C2111 VPWR _44_/a_256_47# -7.56e-19
C2112 _01_ _06_ 0.00157f
C2113 _21_ b[2] 2.14e-19
C2114 _03_ _12_ 2.76e-20
C2115 input6/a_27_47# net19 0.00586f
C2116 input15/a_27_47# net19 0.00236f
C2117 input9/a_75_212# net9 0.0247f
C2118 output19/a_27_47# _42_/a_109_93# 1.56e-20
C2119 _01_ net5 0.0779f
C2120 _34_/a_47_47# _06_ 0.0391f
C2121 input3/a_27_47# p[8] 6.2e-19
C2122 _20_ _47_/a_81_21# 0.0457f
C2123 _35_/a_76_199# net10 0.0146f
C2124 net6 output16/a_27_47# 1.5e-19
C2125 _14_ _27_/a_27_297# 1.66e-21
C2126 _02_ _39_/a_47_47# 0.0127f
C2127 _10_ _01_ 2.22e-19
C2128 _03_ _45_/a_193_297# 2.57e-20
C2129 p[0] net1 0.00473f
C2130 _49_/a_201_297# _31_/a_35_297# 5.52e-20
C2131 VPWR _35_/a_226_297# -8.54e-19
C2132 _44_/a_250_297# p[13] 4.09e-20
C2133 _15_ _19_ 1.46e-20
C2134 _37_/a_27_47# net19 0.0105f
C2135 input5/a_558_47# p[1] 1.61e-21
C2136 _30_/a_109_53# _06_ 1.96e-19
C2137 _18_ net8 1.15e-21
C2138 VPWR _28_/a_109_297# -1.71e-19
C2139 net12 net7 1.57e-19
C2140 net5 _30_/a_109_53# 5.84e-22
C2141 input2/a_27_47# _15_ 3.18e-20
C2142 p[10] p[1] 9.52e-20
C2143 b[2] _52_/a_250_297# 1.6e-19
C2144 _14_ net15 0.0538f
C2145 net16 _38_/a_197_47# 5.89e-19
C2146 net15 _26_/a_29_53# 9.06e-21
C2147 b[3] _42_/a_209_311# 3.71e-19
C2148 _11_ _38_/a_27_47# 0.071f
C2149 _13_ _45_/a_465_47# 0.00134f
C2150 _53_/a_29_53# b[2] 6.22e-19
C2151 _39_/a_47_47# net3 1.66e-20
C2152 output19/a_27_47# input3/a_27_47# 4.77e-21
C2153 net11 input12/a_27_47# 0.00246f
C2154 VPWR net12 0.817f
C2155 net16 _22_ 0.00606f
C2156 net12 p[6] 0.0255f
C2157 _04_ _52_/a_584_47# 2.5e-19
C2158 _16_ _55_/a_217_297# 0.0017f
C2159 _39_/a_285_47# _13_ 0.00451f
C2160 input5/a_381_47# _27_/a_27_297# 1.47e-19
C2161 _39_/a_47_47# _17_ 1.47e-20
C2162 _02_ _13_ 0.0676f
C2163 _12_ _45_/a_205_47# 7.46e-19
C2164 net13 _34_/a_285_47# 4.11e-20
C2165 _03_ net18 2.07e-21
C2166 _36_/a_197_47# net6 6.94e-20
C2167 _44_/a_250_297# net3 0.0088f
C2168 _01_ _31_/a_35_297# 4.27e-19
C2169 _27_/a_27_297# net7 1.22e-19
C2170 _44_/a_250_297# _17_ 0.0336f
C2171 _02_ net19 0.0474f
C2172 _06_ _50_/a_429_93# 0.00169f
C2173 _04_ p[1] 1.74e-21
C2174 _14_ _50_/a_343_93# 9.76e-19
C2175 net4 _50_/a_429_93# 4.16e-19
C2176 _50_/a_223_47# net9 2e-19
C2177 _26_/a_29_53# _50_/a_343_93# 2.61e-19
C2178 _20_ net14 8.01e-20
C2179 p[9] net14 1.05e-19
C2180 input5/a_381_47# net15 7.15e-19
C2181 VPWR _27_/a_27_297# 0.0329f
C2182 net15 p[11] 3.83e-19
C2183 _30_/a_215_297# net17 4.69e-20
C2184 net10 _50_/a_27_47# 3.78e-21
C2185 _12_ net10 7.82e-20
C2186 net16 _50_/a_27_47# 2.35e-20
C2187 input4/a_75_212# _12_ 2.09e-20
C2188 _10_ _50_/a_429_93# 0.00167f
C2189 _12_ net16 0.131f
C2190 net15 net7 2.91e-19
C2191 _31_/a_35_297# _30_/a_109_53# 2.89e-20
C2192 _20_ net1 0.363f
C2193 _06_ _36_/a_109_47# 0.00168f
C2194 _03_ _06_ 0.00635f
C2195 input3/a_27_47# b[1] 1.31e-20
C2196 _43_/a_27_47# _32_/a_27_47# 2.01e-20
C2197 net5 _36_/a_109_47# 0.00144f
C2198 _09_ net1 5.26e-20
C2199 _30_/a_297_297# net1 7.34e-20
C2200 _03_ net5 1.04e-19
C2201 net3 net19 0.611f
C2202 _34_/a_377_297# _06_ 0.00427f
C2203 _26_/a_29_53# _36_/a_27_47# 1.6e-19
C2204 input5/a_558_47# net8 0.00357f
C2205 _17_ net19 0.0269f
C2206 _02_ _50_/a_223_47# 2.51e-20
C2207 _32_/a_109_47# net8 0.0011f
C2208 _26_/a_183_297# _22_ 0.00184f
C2209 _27_/a_277_297# net3 2.71e-19
C2210 net16 _45_/a_193_297# 0.00187f
C2211 VPWR net15 0.61f
C2212 _20_ net6 9.69e-20
C2213 p[9] net6 0.14f
C2214 net6 _09_ 5.43e-20
C2215 _03_ _10_ 0.00244f
C2216 p[5] input11/a_27_47# 0.0433f
C2217 net14 _19_ 0.0512f
C2218 p[10] net8 0.0097f
C2219 _52_/a_93_21# net11 2.8e-19
C2220 _52_/a_93_21# _23_ 0.0166f
C2221 p[5] net18 1.98e-19
C2222 _10_ _43_/a_469_47# 0.00124f
C2223 net14 input2/a_27_47# 0.0102f
C2224 _20_ _49_/a_75_199# 0.0233f
C2225 _19_ net1 2.86e-19
C2226 _35_/a_76_199# _20_ 3.21e-20
C2227 _34_/a_285_47# _21_ 6.94e-20
C2228 _52_/a_93_21# _35_/a_226_47# 4.89e-20
C2229 _49_/a_75_199# _09_ 2.93e-19
C2230 _35_/a_76_199# _09_ 0.0374f
C2231 net13 _30_/a_215_297# 0.0246f
C2232 net15 _37_/a_303_47# 0.00118f
C2233 _14_ input6/a_27_47# 3.75e-21
C2234 _14_ input15/a_27_47# 9.48e-21
C2235 _42_/a_209_311# p[14] 3.45e-22
C2236 _31_/a_285_47# net8 0.00129f
C2237 input2/a_27_47# net1 4.81e-19
C2238 net8 _32_/a_27_47# 0.0275f
C2239 net2 _05_ 4.03e-20
C2240 _50_/a_223_47# _17_ 5.24e-20
C2241 VPWR _50_/a_343_93# -0.0126f
C2242 _01_ net19 4.9e-19
C2243 _45_/a_109_297# VPWR -0.011f
C2244 _04_ net8 0.02f
C2245 net16 net18 0.00585f
C2246 _00_ _15_ 0.207f
C2247 net5 _45_/a_205_47# 8.28e-20
C2248 _03_ _31_/a_35_297# 0.00749f
C2249 _02_ _24_ 0.023f
C2250 _37_/a_27_47# _14_ 0.00137f
C2251 _49_/a_75_199# _19_ 0.0206f
C2252 _35_/a_489_413# _33_/a_209_311# 2.77e-20
C2253 _00_ _47_/a_384_47# 5.15e-20
C2254 _08_ net7 9.54e-25
C2255 VPWR _36_/a_27_47# -0.00832f
C2256 _00_ _47_/a_81_21# 0.0258f
C2257 _10_ _45_/a_205_47# 6.19e-20
C2258 _20_ _22_ 0.183f
C2259 _09_ _22_ 0.0279f
C2260 _45_/a_27_47# _02_ 0.00449f
C2261 p[10] b[3] 3.13e-20
C2262 _26_/a_29_53# net9 0.00343f
C2263 _11_ _18_ 0.484f
C2264 _53_/a_183_297# _02_ 4.14e-19
C2265 _02_ _49_/a_315_47# 0.00134f
C2266 net4 net10 8.28e-22
C2267 VPWR _08_ -0.0171f
C2268 _06_ net10 0.184f
C2269 net16 _06_ 0.0511f
C2270 input4/a_75_212# _06_ 0.00205f
C2271 net4 input4/a_75_212# 0.0189f
C2272 net4 net16 0.155f
C2273 p[6] _08_ 1.55e-19
C2274 net5 net16 0.00461f
C2275 net5 net10 0.0316f
C2276 net5 input4/a_75_212# 0.0104f
C2277 net13 _49_/a_544_297# 3.43e-19
C2278 _29_/a_111_297# net9 8.06e-21
C2279 _37_/a_197_47# net2 4.74e-20
C2280 net13 _25_ 0.00297f
C2281 _03_ _39_/a_47_47# 1.47e-19
C2282 net8 output17/a_27_47# 0.0043f
C2283 _10_ _29_/a_183_297# 6.24e-20
C2284 _30_/a_215_297# _33_/a_109_93# 0.00104f
C2285 _37_/a_27_47# p[11] 4.41e-19
C2286 _02_ _14_ 0.0316f
C2287 _10_ net10 4.45e-19
C2288 _10_ net16 0.0338f
C2289 _10_ input4/a_75_212# 0.00372f
C2290 _31_/a_285_297# b[1] 1.12e-19
C2291 _03_ input9/a_75_212# 9.32e-20
C2292 VPWR input6/a_27_47# 0.00162f
C2293 VPWR input15/a_27_47# 0.0113f
C2294 net4 output16/a_27_47# 0.00706f
C2295 net11 _29_/a_29_53# 0.00514f
C2296 _21_ _30_/a_215_297# 1.48e-19
C2297 input3/a_27_47# _42_/a_109_93# 0.00249f
C2298 _02_ _26_/a_29_53# 0.0466f
C2299 _20_ _12_ 3.9e-19
C2300 net5 output16/a_27_47# 4.08e-20
C2301 _09_ _50_/a_27_47# 1.3e-19
C2302 _12_ _09_ 0.00509f
C2303 p[7] _33_/a_209_311# 1.34e-19
C2304 _45_/a_27_47# _17_ 1.16e-20
C2305 input5/a_841_47# _16_ 8.62e-19
C2306 input5/a_381_47# net9 3.4e-19
C2307 _36_/a_303_47# _25_ 2.03e-21
C2308 _35_/a_226_47# _29_/a_29_53# 2.64e-19
C2309 _52_/a_93_21# _05_ 1.12e-20
C2310 net7 net9 0.00233f
C2311 _04_ _33_/a_209_311# 0.00133f
C2312 _03_ _13_ 1.74e-20
C2313 _02_ output18/a_27_47# 3.6e-19
C2314 VPWR _37_/a_27_47# -0.0178f
C2315 net15 _27_/a_27_297# 0.00888f
C2316 _09_ _45_/a_193_297# 0.00961f
C2317 _14_ net3 0.0295f
C2318 _42_/a_209_311# net2 5.1e-19
C2319 input10/a_27_47# input11/a_27_47# 5.3e-19
C2320 input1/a_75_212# b[1] 4.16e-19
C2321 net14 net17 5.43e-19
C2322 input5/a_381_47# p[13] 0.00153f
C2323 _26_/a_29_53# net3 2.83e-21
C2324 p[11] p[13] 0.00897f
C2325 _49_/a_201_297# _14_ 4.76e-21
C2326 _14_ _17_ 0.489f
C2327 net14 _00_ 4.11e-20
C2328 _26_/a_183_297# _06_ 3.16e-19
C2329 b[1] _05_ 5.29e-20
C2330 VPWR net9 0.5f
C2331 input10/a_27_47# net18 4.16e-20
C2332 input7/a_27_47# net7 0.00318f
C2333 p[13] net7 1.91e-19
C2334 _31_/a_35_297# net10 3.95e-20
C2335 p[3] net9 0.0376f
C2336 _34_/a_47_47# _24_ 6.84e-21
C2337 net17 net1 2.89e-19
C2338 net12 _36_/a_27_47# 0.0185f
C2339 _03_ _27_/a_277_297# 2.1e-20
C2340 _36_/a_197_47# _06_ 6.18e-19
C2341 VPWR p[4] 0.112f
C2342 _02_ net7 0.445f
C2343 _00_ net1 9.43e-19
C2344 p[6] p[4] 0.0051f
C2345 _48_/a_181_47# _07_ 5.93e-19
C2346 b[3] output17/a_27_47# 4.01e-20
C2347 net5 _36_/a_197_47# 0.00254f
C2348 _10_ _26_/a_183_297# 5.74e-19
C2349 _43_/a_193_413# _18_ 0.0413f
C2350 VPWR input7/a_27_47# 0.0768f
C2351 _01_ _49_/a_315_47# 1.82e-19
C2352 VPWR p[13] 0.183f
C2353 VPWR _45_/a_465_47# -5.05e-19
C2354 _00_ _44_/a_93_21# 4.54e-20
C2355 _21_ _15_ 1.13e-21
C2356 _21_ _25_ 0.00164f
C2357 net12 _08_ 0.0269f
C2358 _09_ net18 1.97e-21
C2359 _00_ net6 0.00178f
C2360 VPWR _39_/a_285_47# -9.53e-19
C2361 net3 p[11] 0.00406f
C2362 _10_ _36_/a_197_47# 1.54e-19
C2363 _02_ VPWR 0.33f
C2364 _18_ net2 0.00181f
C2365 input5/a_381_47# net3 0.0299f
C2366 input5/a_62_47# p[0] 1.39e-19
C2367 _01_ _14_ 0.0193f
C2368 _03_ _50_/a_223_47# 1.41e-21
C2369 p[11] _17_ 1.93e-19
C2370 _49_/a_75_199# net17 0.00127f
C2371 _39_/a_47_47# net10 4.72e-22
C2372 _20_ _47_/a_299_297# 0.002f
C2373 _39_/a_47_47# input4/a_75_212# 3.1e-19
C2374 _39_/a_47_47# net16 7.7e-20
C2375 net3 net7 7.45e-20
C2376 net13 net14 2.21e-21
C2377 _13_ _45_/a_205_47# 7.51e-20
C2378 input5/a_664_47# _19_ 2.19e-21
C2379 _53_/a_111_297# _09_ 3.4e-19
C2380 _49_/a_201_297# net7 0.00419f
C2381 VPWR _44_/a_584_47# -2.28e-19
C2382 input9/a_75_212# net10 0.00699f
C2383 _11_ _32_/a_27_47# 1.65e-20
C2384 _20_ _55_/a_80_21# 0.0291f
C2385 _40_/a_109_297# _11_ 0.00522f
C2386 net13 net1 3.51e-19
C2387 input2/a_27_47# input5/a_664_47# 4.47e-21
C2388 VPWR _35_/a_556_47# -7.24e-19
C2389 _20_ net4 3.01e-20
C2390 VPWR net3 0.351f
C2391 p[9] _06_ 0.00205f
C2392 _20_ _06_ 0.133f
C2393 _12_ _52_/a_346_47# 3.8e-19
C2394 net4 _09_ 0.00262f
C2395 _09_ _06_ 0.0965f
C2396 _20_ net5 0.0651f
C2397 p[12] _18_ 3.95e-21
C2398 _28_/a_109_297# net9 3.7e-19
C2399 net5 _09_ 5.18e-19
C2400 VPWR _17_ 0.306f
C2401 VPWR _49_/a_201_297# 0.0185f
C2402 _41_/a_59_75# p[14] 5.13e-20
C2403 _29_/a_29_53# _07_ 1.19e-20
C2404 net13 net6 0.00188f
C2405 _53_/a_29_53# _25_ 0.00146f
C2406 _41_/a_59_75# _11_ 8.7e-19
C2407 _29_/a_29_53# _05_ 3.79e-20
C2408 _13_ net10 4.52e-21
C2409 _13_ net16 0.0198f
C2410 _10_ _20_ 0.179f
C2411 net16 _38_/a_303_47# 6.47e-19
C2412 _10_ _30_/a_297_297# 1.25e-20
C2413 _10_ _09_ 0.0222f
C2414 _10_ p[9] 0.00225f
C2415 net3 _37_/a_303_47# 0.00133f
C2416 _42_/a_368_53# net3 3.82e-19
C2417 net12 net9 0.0596f
C2418 net13 _49_/a_75_199# 3.2e-19
C2419 net13 _35_/a_76_199# 0.0337f
C2420 _16_ _55_/a_472_297# 3.71e-19
C2421 _37_/a_303_47# _17_ 1.23e-20
C2422 _01_ net7 0.233f
C2423 _00_ _22_ 0.477f
C2424 _03_ _24_ 9.46e-20
C2425 net11 _23_ 0.0461f
C2426 _44_/a_256_47# net3 0.00101f
C2427 _39_/a_129_47# _17_ 1.38e-20
C2428 _36_/a_303_47# net6 1.25e-19
C2429 _13_ output16/a_27_47# 4.58e-19
C2430 net5 _19_ 6.41e-21
C2431 net12 p[4] 5.33e-19
C2432 _35_/a_226_47# net11 3.21e-19
C2433 input13/a_27_47# net1 1.9e-19
C2434 _35_/a_226_47# _23_ 4.21e-19
C2435 input5/a_558_47# net2 5.99e-21
C2436 _45_/a_27_47# _03_ 2.06e-20
C2437 VPWR _01_ 0.521f
C2438 net15 input6/a_27_47# 0.00115f
C2439 net15 input15/a_27_47# 0.00325f
C2440 _21_ net14 7.17e-21
C2441 _52_/a_93_21# _18_ 1.97e-19
C2442 _03_ _49_/a_315_47# 9.22e-19
C2443 VPWR _34_/a_47_47# 0.0372f
C2444 _02_ net12 2.28e-19
C2445 p[6] _34_/a_47_47# 4.28e-19
C2446 p[10] net2 0.0632f
C2447 VPWR _27_/a_109_297# -2.45e-19
C2448 input14/a_27_47# net14 0.0232f
C2449 _20_ _31_/a_35_297# 1.69e-19
C2450 net16 _50_/a_223_47# 4.77e-21
C2451 _21_ net1 0.0252f
C2452 _00_ _50_/a_27_47# 0.00197f
C2453 _00_ _12_ 0.00396f
C2454 net13 _22_ 4.63e-20
C2455 net11 _48_/a_27_47# 0.0179f
C2456 _37_/a_27_47# net15 0.0541f
C2457 VPWR _30_/a_109_53# 0.0012f
C2458 _34_/a_129_47# _06_ 5.3e-19
C2459 _04_ _43_/a_193_413# 5.67e-21
C2460 _14_ _43_/a_469_47# 0.00259f
C2461 input5/a_62_47# _19_ 0.00159f
C2462 _30_/a_109_53# p[3] 3.23e-20
C2463 _32_/a_197_47# net8 3.39e-20
C2464 _03_ _26_/a_29_53# 7.93e-21
C2465 _27_/a_27_297# input7/a_27_47# 0.00119f
C2466 _21_ net6 2.92e-20
C2467 _40_/a_109_297# net2 0.0011f
C2468 net15 net9 8.49e-20
C2469 _02_ _27_/a_27_297# 0.00179f
C2470 _03_ _29_/a_111_297# 7.48e-19
C2471 _00_ _45_/a_193_297# 4.38e-20
C2472 input12/a_27_47# p[7] 3.2e-20
C2473 _04_ net2 0.158f
C2474 _30_/a_215_297# net8 8.14e-21
C2475 net8 _32_/a_303_47# 2.22e-34
C2476 _06_ _52_/a_346_47# 0.0031f
C2477 _15_ _50_/a_515_93# 0.00147f
C2478 _31_/a_35_297# _19_ 1.47e-19
C2479 _35_/a_76_199# _33_/a_109_93# 3.08e-19
C2480 _20_ _39_/a_47_47# 2.3e-20
C2481 _21_ _49_/a_75_199# 6.64e-19
C2482 _35_/a_76_199# _21_ 0.0175f
C2483 net5 _52_/a_346_47# 7.03e-19
C2484 _39_/a_47_47# _09_ 7.7e-21
C2485 net15 p[13] 1.48e-19
C2486 input2/a_27_47# _31_/a_35_297# 0.00136f
C2487 net15 input7/a_27_47# 1.88e-19
C2488 _15_ _43_/a_27_47# 8.96e-20
C2489 net13 _12_ 0.00632f
C2490 net13 _50_/a_27_47# 7.27e-21
C2491 _02_ net15 0.0806f
C2492 VPWR _50_/a_429_93# -3.61e-19
C2493 net16 _24_ 6.93e-19
C2494 net3 _27_/a_27_297# 0.0166f
C2495 _50_/a_343_93# net9 6.64e-19
C2496 _03_ net7 0.078f
C2497 net6 _52_/a_250_297# 0.00133f
C2498 _27_/a_27_297# _17_ 6.78e-22
C2499 _20_ _13_ 7.38e-21
C2500 _03_ _31_/a_117_297# 5.32e-19
C2501 net11 _38_/a_27_47# 1.68e-20
C2502 net6 _53_/a_29_53# 2.11e-20
C2503 _01_ net12 1.67e-21
C2504 net11 _05_ 2.76e-19
C2505 net11 _07_ 0.0206f
C2506 _13_ _09_ 0.0927f
C2507 _45_/a_27_47# net16 8.68e-19
C2508 _41_/a_59_75# p[12] 0.0547f
C2509 _45_/a_27_47# input4/a_75_212# 2.18e-20
C2510 net2 output17/a_27_47# 0.0285f
C2511 VPWR _36_/a_109_47# -4.66e-19
C2512 _33_/a_109_93# _22_ 1.34e-22
C2513 _07_ _23_ 1.27e-19
C2514 _35_/a_76_199# _52_/a_250_297# 3.4e-21
C2515 _36_/a_27_47# net9 0.00493f
C2516 net12 _34_/a_47_47# 0.0385f
C2517 _00_ _47_/a_299_297# 7.59e-21
C2518 _03_ VPWR 0.845f
C2519 input6/a_27_47# input15/a_27_47# 5.3e-19
C2520 _03_ p[3] 0.00348f
C2521 _20_ net19 1.29e-19
C2522 _21_ _22_ 0.00314f
C2523 net15 net3 0.394f
C2524 p[9] net19 0.0729f
C2525 _35_/a_226_47# _07_ 8.96e-19
C2526 _02_ _50_/a_343_93# 6.94e-19
C2527 VPWR _34_/a_377_297# -0.00192f
C2528 _35_/a_226_47# _05_ 0.0134f
C2529 VPWR _43_/a_469_47# -2.75e-19
C2530 _45_/a_109_297# _02_ 8.44e-19
C2531 _00_ _55_/a_80_21# 5.5e-19
C2532 _34_/a_377_297# p[6] 5.39e-19
C2533 _49_/a_201_297# net15 1.41e-19
C2534 net15 _17_ 0.195f
C2535 _15_ net8 1.79e-19
C2536 p[10] b[1] 0.286f
C2537 net5 net17 4.21e-21
C2538 _08_ net9 7.71e-21
C2539 net4 _00_ 0.0166f
C2540 _00_ _06_ 0.1f
C2541 net12 _30_/a_109_53# 4.25e-20
C2542 _37_/a_27_47# input6/a_27_47# 9.35e-19
C2543 net5 _00_ 0.00954f
C2544 _01_ _27_/a_27_297# 8.04e-19
C2545 net14 p[1] 0.0025f
C2546 _26_/a_29_53# net10 3.48e-22
C2547 _37_/a_27_47# input15/a_27_47# 3.27e-19
C2548 _52_/a_93_21# _04_ 2.35e-19
C2549 _02_ _36_/a_27_47# 9.37e-20
C2550 _47_/a_81_21# net8 2.08e-21
C2551 _30_/a_215_297# _33_/a_209_311# 1.56e-19
C2552 _16_ _42_/a_209_311# 0.00129f
C2553 _12_ _33_/a_109_93# 9.75e-20
C2554 _27_/a_27_297# _27_/a_109_297# -3.68e-20
C2555 _48_/a_27_47# _07_ 0.0524f
C2556 _10_ _00_ 0.301f
C2557 p[1] net1 0.0291f
C2558 net14 _50_/a_515_93# 1.39e-20
C2559 input3/a_27_47# _42_/a_209_311# 1.56e-19
C2560 _20_ _50_/a_223_47# 1.71e-19
C2561 _21_ _50_/a_27_47# 3.38e-21
C2562 _21_ _12_ 7.99e-20
C2563 _52_/a_250_297# _22_ 0.099f
C2564 _11_ _54_/a_75_212# 3.22e-20
C2565 _17_ _50_/a_343_93# 0.0015f
C2566 output18/a_27_47# net16 3.45e-19
C2567 _02_ _08_ 2.26e-20
C2568 _45_/a_109_297# _17_ 4.29e-22
C2569 input2/a_27_47# net19 2.9e-23
C2570 _04_ b[1] 5.79e-19
C2571 _53_/a_29_53# _22_ 0.00749f
C2572 _01_ net15 0.0314f
C2573 _00_ _43_/a_297_47# 1.26e-19
C2574 net14 _43_/a_27_47# 4.87e-20
C2575 VPWR _45_/a_205_47# -1.62e-19
C2576 _03_ _35_/a_226_297# 0.00101f
C2577 input8/a_27_47# _31_/a_285_297# 1.04e-19
C2578 net13 _06_ 0.0766f
C2579 net13 net4 2.48e-19
C2580 p[5] p[6] 0.198f
C2581 VPWR p[5] 0.092f
C2582 _31_/a_285_297# _05_ 6.12e-19
C2583 net13 net5 0.127f
C2584 output18/a_27_47# output16/a_27_47# 7.85e-19
C2585 net6 _50_/a_515_93# 4.7e-19
C2586 _08_ _35_/a_556_47# 7.71e-19
C2587 _26_/a_183_297# _14_ 6.98e-22
C2588 _52_/a_93_21# b[2] 1.63e-19
C2589 _31_/a_35_297# net17 0.0514f
C2590 b[3] _15_ 0.00162f
C2591 net13 _10_ 0.00151f
C2592 _16_ _18_ 0.144f
C2593 _12_ _52_/a_250_297# 0.0139f
C2594 VPWR _29_/a_183_297# -8.13e-19
C2595 _21_ input5/a_664_47# 9.42e-22
C2596 _03_ net12 0.0268f
C2597 _36_/a_303_47# _06_ 5.3e-19
C2598 net6 _43_/a_27_47# 9.07e-20
C2599 _01_ _50_/a_343_93# 0.0131f
C2600 p[2] p[1] 0.188f
C2601 VPWR net10 0.362f
C2602 _12_ _53_/a_29_53# 3.46e-20
C2603 VPWR net16 0.518f
C2604 VPWR input4/a_75_212# 0.06f
C2605 net10 p[3] 8.58e-19
C2606 p[6] net10 0.0023f
C2607 net5 _36_/a_303_47# 0.00256f
C2608 _34_/a_377_297# net12 0.00251f
C2609 b[1] output17/a_27_47# 0.00945f
C2610 p[13] net9 1.72e-19
C2611 _09_ _24_ 0.0202f
C2612 net3 input6/a_27_47# 2.52e-19
C2613 net3 input15/a_27_47# 8.74e-20
C2614 _52_/a_584_47# _22_ 6.24e-19
C2615 _21_ net18 0.00215f
C2616 input8/a_27_47# _05_ 1.58e-19
C2617 net14 net8 0.0516f
C2618 _07_ _05_ 1.21e-19
C2619 input6/a_27_47# _17_ 7.13e-22
C2620 _02_ net9 0.00611f
C2621 _10_ _36_/a_303_47# 4.09e-19
C2622 input15/a_27_47# _17_ 6.14e-19
C2623 input13/a_27_47# _06_ 7.75e-19
C2624 VPWR output16/a_27_47# 0.122f
C2625 _39_/a_47_47# _00_ 1.85e-20
C2626 _45_/a_27_47# _09_ 0.00823f
C2627 _53_/a_111_297# _21_ 4.38e-19
C2628 input5/a_558_47# _42_/a_109_93# 1.75e-19
C2629 net8 net1 0.381f
C2630 _53_/a_183_297# _09_ 4.18e-19
C2631 p[0] net7 1.36e-19
C2632 _03_ _27_/a_27_297# 2.68e-19
C2633 _04_ _29_/a_29_53# 0.0408f
C2634 _37_/a_27_47# net3 0.094f
C2635 _09_ _49_/a_315_47# 1.11e-20
C2636 net13 _31_/a_35_297# 1.86e-20
C2637 _02_ p[13] 7.58e-20
C2638 _06_ _33_/a_109_93# 9.13e-19
C2639 _37_/a_27_47# _17_ 0.00277f
C2640 input5/a_841_47# input5/a_558_47# -4.44e-34
C2641 _00_ _44_/a_250_297# 6.39e-20
C2642 _34_/a_47_47# _08_ 0.00123f
C2643 p[10] _42_/a_109_93# 1.82e-21
C2644 _21_ net4 0.00535f
C2645 _21_ _06_ 0.143f
C2646 _02_ _39_/a_285_47# 0.0019f
C2647 net3 net9 5.09e-20
C2648 p[9] _14_ 2.62e-21
C2649 _20_ _14_ 0.144f
C2650 VPWR p[0] 0.0836f
C2651 _21_ net5 0.00784f
C2652 VPWR _26_/a_183_297# -3.03e-19
C2653 _20_ _26_/a_29_53# 0.00447f
C2654 _17_ net9 2.89e-23
C2655 _03_ net15 4.26e-20
C2656 net10 _35_/a_226_297# 2.48e-19
C2657 _43_/a_27_47# _22_ 0.091f
C2658 _53_/a_29_53# net18 0.0118f
C2659 net12 p[5] 0.00294f
C2660 _49_/a_75_199# net8 0.00214f
C2661 _00_ _13_ 3.77e-20
C2662 _10_ _21_ 0.00421f
C2663 net15 _43_/a_469_47# 7.41e-19
C2664 net3 p[13] 3.65e-19
C2665 _19_ _49_/a_315_47# 1.33e-19
C2666 _09_ _29_/a_111_297# 5.79e-20
C2667 net17 net19 8.84e-23
C2668 VPWR _36_/a_197_47# -5.24e-19
C2669 _04_ _42_/a_109_93# 5.77e-22
C2670 _15_ p[14] 5.32e-19
C2671 p[2] net8 0.00956f
C2672 _02_ net3 9.52e-20
C2673 _39_/a_285_47# _17_ 7.36e-21
C2674 _11_ _25_ 7.05e-19
C2675 net14 b[3] 0.0172f
C2676 _11_ _15_ 0.113f
C2677 net13 input9/a_75_212# 4.4e-19
C2678 _05_ _33_/a_296_53# 4.53e-19
C2679 _14_ _19_ 2.71e-21
C2680 _02_ _17_ 0.00482f
C2681 net4 _52_/a_250_297# 0.00136f
C2682 _06_ _52_/a_250_297# 0.0058f
C2683 _47_/a_384_47# _11_ 7.23e-20
C2684 net12 net10 0.539f
C2685 net5 _52_/a_250_297# 0.018f
C2686 p[9] p[11] 0.114f
C2687 VPWR input10/a_27_47# 0.00986f
C2688 net4 _53_/a_29_53# 3.26e-19
C2689 _53_/a_29_53# _06_ 0.0709f
C2690 _47_/a_81_21# _11_ 0.0454f
C2691 input10/a_27_47# p[6] 0.00214f
C2692 _01_ net9 0.157f
C2693 _12_ _43_/a_27_47# 2.33e-21
C2694 _20_ net7 0.0257f
C2695 _34_/a_47_47# net9 1.41e-20
C2696 _09_ net7 0.00258f
C2697 _44_/a_93_21# b[3] 0.00491f
C2698 _10_ _52_/a_250_297# 0.00368f
C2699 _04_ VGND 0.478f
C2700 _03_ VGND 0.481f
C2701 net10 VGND 0.909f
C2702 _30_/a_465_297# VGND 0.00105f
C2703 _30_/a_392_297# VGND 7.67e-19
C2704 _30_/a_297_297# VGND -4.43e-19
C2705 _30_/a_109_53# VGND 0.152f
C2706 _30_/a_215_297# VGND 0.158f
C2707 _05_ VGND 0.906f
C2708 net8 VGND 0.791f
C2709 _31_/a_285_297# VGND 1.12e-20
C2710 _31_/a_117_297# VGND -0.00177f
C2711 _31_/a_35_297# VGND 0.246f
C2712 _32_/a_303_47# VGND -4.83e-19
C2713 _32_/a_197_47# VGND 8.12e-20
C2714 _32_/a_109_47# VGND 1.05e-19
C2715 _32_/a_27_47# VGND 0.198f
C2716 _50_/a_615_93# VGND -5.19e-19
C2717 _50_/a_515_93# VGND -4.75e-19
C2718 _50_/a_429_93# VGND 4.71e-19
C2719 _50_/a_343_93# VGND 0.171f
C2720 _50_/a_223_47# VGND 0.157f
C2721 _50_/a_27_47# VGND 0.255f
C2722 _07_ VGND 0.483f
C2723 _06_ VGND 1.91f
C2724 net13 VGND 0.524f
C2725 _33_/a_368_53# VGND 2.38e-19
C2726 _33_/a_296_53# VGND -1.43e-19
C2727 _33_/a_209_311# VGND 0.136f
C2728 _33_/a_109_93# VGND 0.145f
C2729 net12 VGND 0.874f
C2730 _34_/a_285_47# VGND 0.0144f
C2731 _34_/a_129_47# VGND -8.76e-20
C2732 _34_/a_377_297# VGND -9.51e-19
C2733 _34_/a_47_47# VGND 0.289f
C2734 _23_ VGND 0.266f
C2735 _09_ VGND 0.544f
C2736 _08_ VGND 0.293f
C2737 _35_/a_556_47# VGND 1.95e-19
C2738 _35_/a_226_297# VGND -4.55e-19
C2739 _35_/a_489_413# VGND 0.0246f
C2740 _35_/a_226_47# VGND 0.151f
C2741 _35_/a_76_199# VGND 0.137f
C2742 p[9] VGND 0.51f
C2743 input15/a_27_47# VGND 0.223f
C2744 _24_ VGND 0.127f
C2745 _12_ VGND 1.2f
C2746 _52_/a_584_47# VGND -0.00112f
C2747 _52_/a_346_47# VGND -0.00175f
C2748 _52_/a_256_47# VGND -0.00161f
C2749 _52_/a_250_297# VGND 0.0246f
C2750 _52_/a_93_21# VGND 0.133f
C2751 _10_ VGND 1.75f
C2752 _36_/a_303_47# VGND 8.14e-19
C2753 _36_/a_197_47# VGND -3.75e-19
C2754 _36_/a_109_47# VGND 3.56e-19
C2755 _36_/a_27_47# VGND 0.196f
C2756 _53_/a_183_297# VGND -4.34e-19
C2757 _53_/a_111_297# VGND -2.89e-19
C2758 _53_/a_29_53# VGND 0.163f
C2759 p[8] VGND 1.26f
C2760 input14/a_27_47# VGND 0.247f
C2761 _11_ VGND 0.358f
C2762 _37_/a_303_47# VGND -1.63e-19
C2763 _37_/a_197_47# VGND -4.58e-19
C2764 _37_/a_109_47# VGND -7.9e-19
C2765 _37_/a_27_47# VGND 0.16f
C2766 p[7] VGND 0.887f
C2767 input13/a_27_47# VGND 0.255f
C2768 net18 VGND 0.463f
C2769 _25_ VGND 0.39f
C2770 _54_/a_75_212# VGND 0.263f
C2771 _38_/a_303_47# VGND 1.78e-19
C2772 _38_/a_197_47# VGND 2.29e-19
C2773 _38_/a_109_47# VGND 2.3e-19
C2774 _38_/a_27_47# VGND 0.183f
C2775 net19 VGND 0.31f
C2776 _22_ VGND 0.256f
C2777 _14_ VGND 0.454f
C2778 _15_ VGND 0.487f
C2779 _55_/a_300_47# VGND -0.00109f
C2780 _55_/a_472_297# VGND -0.00188f
C2781 _55_/a_217_297# VGND -0.00225f
C2782 _55_/a_80_21# VGND 0.213f
C2783 p[6] VGND 0.742f
C2784 input12/a_27_47# VGND 0.248f
C2785 net9 VGND 0.685f
C2786 p[3] VGND 0.825f
C2787 input9/a_75_212# VGND 0.276f
C2788 _39_/a_285_47# VGND 0.0128f
C2789 _39_/a_129_47# VGND -0.00126f
C2790 _39_/a_377_297# VGND -6.28e-19
C2791 _39_/a_47_47# VGND 0.266f
C2792 net11 VGND 1.25f
C2793 p[5] VGND 0.76f
C2794 input11/a_27_47# VGND 0.235f
C2795 p[2] VGND 0.769f
C2796 input8/a_27_47# VGND 0.265f
C2797 p[4] VGND 1.25f
C2798 input10/a_27_47# VGND 0.211f
C2799 net7 VGND 0.881f
C2800 p[1] VGND 0.772f
C2801 input7/a_27_47# VGND 0.265f
C2802 p[14] VGND 0.988f
C2803 input6/a_27_47# VGND 0.205f
C2804 net5 VGND 2.04f
C2805 p[13] VGND 0.557f
C2806 input5/a_841_47# VGND 0.187f
C2807 input5/a_664_47# VGND 0.144f
C2808 input5/a_558_47# VGND 0.163f
C2809 input5/a_381_47# VGND 0.107f
C2810 input5/a_62_47# VGND 0.218f
C2811 p[12] VGND 1.3f
C2812 input4/a_75_212# VGND 0.263f
C2813 p[11] VGND 0.865f
C2814 input3/a_27_47# VGND 0.249f
C2815 net2 VGND 1.5f
C2816 p[10] VGND 0.79f
C2817 input2/a_27_47# VGND 0.194f
C2818 net1 VGND 0.855f
C2819 p[0] VGND 1.01f
C2820 VPWR VGND 40.2f
C2821 input1/a_75_212# VGND 0.268f
C2822 b[3] VGND 0.546f
C2823 output19/a_27_47# VGND 0.534f
C2824 b[2] VGND 0.593f
C2825 output18/a_27_47# VGND 0.601f
C2826 _40_/a_297_297# VGND -5.1e-19
C2827 _40_/a_191_297# VGND -9.29e-19
C2828 _40_/a_109_297# VGND -0.00181f
C2829 b[1] VGND 0.526f
C2830 net17 VGND 0.385f
C2831 output17/a_27_47# VGND 0.545f
C2832 _41_/a_145_75# VGND 3.75e-19
C2833 _41_/a_59_75# VGND 0.191f
C2834 b[0] VGND 0.708f
C2835 output16/a_27_47# VGND 0.616f
C2836 _16_ VGND 0.119f
C2837 _42_/a_368_53# VGND -4.05e-19
C2838 _42_/a_209_311# VGND 0.135f
C2839 _42_/a_109_93# VGND 0.153f
C2840 _17_ VGND 0.563f
C2841 _00_ VGND 0.516f
C2842 _43_/a_369_47# VGND -8.43e-19
C2843 _43_/a_297_47# VGND -1.33e-19
C2844 _43_/a_193_413# VGND 0.122f
C2845 _43_/a_27_47# VGND 0.209f
C2846 net6 VGND 1f
C2847 net4 VGND 0.888f
C2848 _26_/a_183_297# VGND 2.42e-19
C2849 _26_/a_111_297# VGND -2.75e-19
C2850 _26_/a_29_53# VGND 0.218f
C2851 _01_ VGND 0.244f
C2852 net14 VGND 0.958f
C2853 net3 VGND 0.786f
C2854 net15 VGND 0.673f
C2855 _27_/a_277_297# VGND -4.65e-19
C2856 _27_/a_205_297# VGND -3.36e-19
C2857 _27_/a_109_297# VGND -6.15e-19
C2858 _27_/a_27_297# VGND 0.147f
C2859 _18_ VGND 0.159f
C2860 _44_/a_584_47# VGND -0.00145f
C2861 _44_/a_346_47# VGND -0.00198f
C2862 _44_/a_256_47# VGND -0.00184f
C2863 _44_/a_250_297# VGND 0.0219f
C2864 _44_/a_93_21# VGND 0.128f
C2865 net16 VGND 0.375f
C2866 _13_ VGND 0.496f
C2867 _45_/a_465_47# VGND -8.14e-19
C2868 _45_/a_205_47# VGND -2.47e-19
C2869 _45_/a_193_297# VGND -0.00131f
C2870 _45_/a_109_297# VGND -0.00108f
C2871 _45_/a_27_47# VGND 0.187f
C2872 _28_/a_109_297# VGND -9.87e-19
C2873 _29_/a_183_297# VGND 4.41e-19
C2874 _29_/a_111_297# VGND -1.9e-19
C2875 _29_/a_29_53# VGND 0.234f
C2876 _19_ VGND 0.497f
C2877 _47_/a_384_47# VGND -2.05e-19
C2878 _47_/a_299_297# VGND 0.0344f
C2879 _47_/a_81_21# VGND 0.136f
C2880 _48_/a_181_47# VGND 3.03e-19
C2881 _48_/a_109_47# VGND 9.44e-19
C2882 _48_/a_27_47# VGND 0.232f
C2883 _21_ VGND 0.586f
C2884 _20_ VGND 0.709f
C2885 _02_ VGND 2.08f
C2886 _49_/a_315_47# VGND -0.0034f
C2887 _49_/a_208_47# VGND -0.00164f
C2888 _49_/a_544_297# VGND -0.00256f
C2889 _49_/a_201_297# VGND -5.82e-19
C2890 _49_/a_75_199# VGND 0.205f
.ends

.GLOBAL VDD
.GLOBAL GND
.end
