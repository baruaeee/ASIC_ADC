* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : pre_therm1                                   *
* Netlisted  : Wed Dec 11 23:57:00 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733957813110                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733957813110 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3.3e-07 W=8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733957813110

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733957813111                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733957813111 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733957813111

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv12f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv12f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_733957813110 $T=340 555 0 0 $X=-65 $Y=405
X5 VDD Y A pfet_01v8_CDNS_733957813111 $T=385 2785 0 0 $X=-60 $Y=2605
.ends inv12f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733957813112                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733957813112 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=9.5e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733957813112

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733957813113                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733957813113 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733957813113

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv15f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv15f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_733957813112 $T=215 700 0 0 $X=-190 $Y=550
X5 VDD Y A pfet_01v8_CDNS_733957813113 $T=620 2635 0 0 $X=175 $Y=2455
.ends inv15f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733957813114                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733957813114 1 2 3
** N=7 EP=3 FDC=1
M0 2 2 1 3 pfet_01v8 L=1.5e-07 W=1e-06 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733957813114

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733957813115                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733957813115 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 pfet_01v8 L=1.05e-06 W=5.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733957813115

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: div_fixed                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt div_fixed A VSS Y
** N=8 EP=3 FDC=2
X4 Y VSS A pfet_01v8_CDNS_733957813114 $T=470 1900 0 180 $X=-125 $Y=720
X5 A Y VSS A pfet_01v8_CDNS_733957813115 $T=1625 3880 1 270 $X=895 $Y=2385
.ends div_fixed

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733957813116                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733957813116 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6.75e-07 W=4.8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733957813116

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733957813117                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733957813117 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.65e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733957813117

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv14f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv14f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_733957813116 $T=350 675 0 0 $X=-55 $Y=525
X5 VDD Y A pfet_01v8_CDNS_733957813117 $T=445 2705 0 0 $X=0 $Y=2525
.ends inv14f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733957813118                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733957813118 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.6e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733957813118

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv11f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv11f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_733957813112 $T=215 700 0 0 $X=-190 $Y=550
X5 VDD Y A pfet_01v8_CDNS_733957813118 $T=350 2610 0 0 $X=-95 $Y=2430
.ends inv11f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733957813119                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733957813119 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.55e-07 W=9.45e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733957813119

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131110                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131110 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.45e-07 W=8.65e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131110

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv10f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv10f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_733957813119 $T=425 555 0 0 $X=20 $Y=405
X5 VDD Y A pfet_01v8_CDNS_7339578131110 $T=385 2670 0 0 $X=-60 $Y=2490
.ends inv10f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131111                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131111 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=9.9e-07 W=4.9e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131111

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131112                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131112 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.65e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131112

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv08f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv08f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7339578131111 $T=1280 740 0 90 $X=640 $Y=335
X5 VDD Y A pfet_01v8_CDNS_7339578131112 $T=360 2755 0 0 $X=-85 $Y=2575
.ends inv08f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131113                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131113 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=6.95e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131113

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131114                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131114 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=4e-07 W=6.5e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131114

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv05f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv05f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VDD Y A pfet_01v8_CDNS_7339578131113 $T=360 2825 0 0 $X=-85 $Y=2645
X5 VSS Y A nfet_01v8_CDNS_7339578131114 $T=315 630 0 0 $X=-90 $Y=480
.ends inv05f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131115                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131115 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.5e-07 W=8e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131115

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131116                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131116 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=2.85e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131116

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv02f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv02f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VDD Y A pfet_01v8_CDNS_7339578131115 $T=335 2855 0 0 $X=-110 $Y=2675
X5 VSS Y A nfet_01v8_CDNS_7339578131116 $T=315 640 0 0 $X=-90 $Y=490
.ends inv02f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131117                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131117 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3e-07 W=9.8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131117

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131118                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131118 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.55e-07 W=5.7e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131118

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv07f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv07f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7339578131117 $T=315 460 0 0 $X=-90 $Y=310
X5 VDD Y A pfet_01v8_CDNS_7339578131118 $T=360 2950 0 0 $X=-85 $Y=2770
.ends inv07f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131119                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131119 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.9e-07 W=6.2e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131119

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131120                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131120 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6e-07 W=7.05e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131120

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv04f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv04f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VDD Y A pfet_01v8_CDNS_7339578131119 $T=380 2650 0 0 $X=-65 $Y=2470
X5 VSS Y A nfet_01v8_CDNS_7339578131120 $T=280 715 0 0 $X=-125 $Y=565
.ends inv04f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131121                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131121 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=5.5e-07 W=5.4e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131121

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131122                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131122 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.6e-07 W=8.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131122

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv13f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv13f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7339578131121 $T=360 720 0 0 $X=-45 $Y=570
X5 VDD Y A pfet_01v8_CDNS_7339578131122 $T=385 2685 0 0 $X=-60 $Y=2505
.ends inv13f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131123                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131123 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.1e-06 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131123

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131124                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131124 1 2 3
** N=9 EP=3 FDC=2
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.7e-07 $X=0 $Y=0 $dt=8
M1 1 3 2 1 pfet_01v8 L=1.5e-07 W=7.7e-07 $X=430 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131124

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv09f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv09f VDD VSS A Y
** N=9 EP=4 FDC=3
X4 VSS Y A nfet_01v8_CDNS_7339578131123 $T=905 695 0 90 $X=335 $Y=290
X5 VDD Y A pfet_01v8_CDNS_7339578131124 $T=400 2840 0 0 $X=-45 $Y=2660
.ends inv09f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131125                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131125 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=3.2e-07 W=7.25e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131125

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131126                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131126 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=4.35e-07 W=5.6e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131126

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv06f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv06f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7339578131125 $T=395 685 0 0 $X=-10 $Y=535
X5 VDD Y A pfet_01v8_CDNS_7339578131126 $T=335 3005 0 0 $X=-110 $Y=2825
.ends inv06f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131127                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131127 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=3.5e-07 W=6.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131127

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131128                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131128 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=4.5e-07 W=6.4e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131128

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv03f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv03f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VDD Y A pfet_01v8_CDNS_7339578131127 $T=335 3045 0 0 $X=-110 $Y=2865
X5 VSS Y A nfet_01v8_CDNS_7339578131128 $T=290 640 0 0 $X=-115 $Y=490
.ends inv03f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131129                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131129 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6.5e-07 W=4.45e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131129

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131130                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131130 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=6.3e-07 W=7.9e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131130

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv01f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv01f VDD VSS A Y
** N=9 EP=4 FDC=2
X4 VSS Y A nfet_01v8_CDNS_7339578131129 $T=295 475 0 0 $X=-110 $Y=325
X5 VDD Y A pfet_01v8_CDNS_7339578131130 $T=295 2820 0 0 $X=-150 $Y=2640
.ends inv01f

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_7339578131131                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_7339578131131 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 pfet_01v8 L=2.5e-07 W=5.5e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_7339578131131

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131132                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131132 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 nfet_01v8 L=5.5e-07 W=4.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131132

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: preamp1F                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt preamp1F VDD VSS A Y
** N=9 EP=4 FDC=2
X3 Y VSS A VDD pfet_01v8_CDNS_7339578131131 $T=840 2840 0 90 $X=110 $Y=2395
X4 Y VDD A VSS nfet_01v8_CDNS_7339578131132 $T=610 1275 0 270 $X=460 $Y=320
.ends preamp1F

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7339578131133                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7339578131133 1 2 3 4
** N=10 EP=4 FDC=1
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=1.02e-06 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7339578131133

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: preampF                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt preampF VDD VSS A Y
** N=9 EP=4 FDC=2
X3 Y VSS A VDD pfet_01v8_CDNS_733957813115 $T=825 3430 0 270 $X=645 $Y=1935
X6 Y VDD A VSS nfet_01v8_CDNS_7339578131133 $T=430 485 1 180 $X=-125 $Y=335
.ends preampF

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pre_therm1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pre_therm1 IN VDD VSS Y01 Y02 Y03 Y04 Y05 Y06 Y07
+ Y08 Y09 Y10 Y11 Y12 Y13 Y14 Y15
** N=36 EP=18 FDC=37
X43 VDD VSS 9 Y12 inv12f $T=6585 8280 1 0 $X=6405 $Y=3835
X44 VDD VSS 9 Y15 inv15f $T=7525 8280 0 0 $X=7335 $Y=8015
X45 IN VSS 9 div_fixed $T=0 8280 0 0 $X=-180 $Y=8015
X46 VDD VSS 9 Y14 inv14f $T=9405 8280 1 0 $X=9225 $Y=3835
X47 VDD VSS 9 Y11 inv11f $T=5775 8280 0 0 $X=5585 $Y=8015
X48 VDD VSS 9 Y10 inv10f $T=4080 8280 0 0 $X=3900 $Y=8015
X49 VDD VSS IN Y08 inv08f $T=3260 8280 1 0 $X=3080 $Y=3835
X50 VDD VSS 13 Y05 inv05f $T=9405 0 0 0 $X=9225 $Y=-265
X51 VDD VSS 4 Y02 inv02f $T=3260 0 0 0 $X=3080 $Y=-265
X52 VDD VSS IN Y07 inv07f $T=1630 8280 1 0 $X=1450 $Y=3835
X53 VDD VSS 13 Y04 inv04f $T=7900 0 0 0 $X=7720 $Y=-265
X54 VDD VSS 9 Y13 inv13f $T=7965 8280 1 0 $X=7785 $Y=3835
X55 VDD VSS IN Y09 inv09f $T=4955 8280 1 0 $X=4765 $Y=3835
X56 VDD VSS IN Y06 inv06f $T=0 8280 1 0 $X=-180 $Y=3835
X57 VDD VSS 13 Y03 inv03f $T=6270 0 0 0 $X=6090 $Y=-265
X58 VDD VSS 4 Y01 inv01f $T=1630 0 0 0 $X=1450 $Y=-265
X59 VDD VSS IN 13 preamp1F $T=4640 0 0 0 $X=4460 $Y=-265
X60 VDD VSS IN 4 preampF $T=0 0 0 0 $X=-180 $Y=-265
.ends pre_therm1
