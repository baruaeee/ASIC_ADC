magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 364 29 370
rect -29 330 -17 364
rect -29 324 29 330
rect -29 -330 29 -324
rect -29 -364 -17 -330
rect -29 -370 29 -364
<< pwell >>
rect -211 -502 211 502
<< nmos >>
rect -15 -292 15 292
<< ndiff >>
rect -73 280 -15 292
rect -73 -280 -61 280
rect -27 -280 -15 280
rect -73 -292 -15 -280
rect 15 280 73 292
rect 15 -280 27 280
rect 61 -280 73 280
rect 15 -292 73 -280
<< ndiffc >>
rect -61 -280 -27 280
rect 27 -280 61 280
<< psubdiff >>
rect -175 432 -79 466
rect 79 432 175 466
rect -175 370 -141 432
rect 141 370 175 432
rect -175 -432 -141 -370
rect 141 -432 175 -370
rect -175 -466 -79 -432
rect 79 -466 175 -432
<< psubdiffcont >>
rect -79 432 79 466
rect -175 -370 -141 370
rect 141 -370 175 370
rect -79 -466 79 -432
<< poly >>
rect -33 364 33 380
rect -33 330 -17 364
rect 17 330 33 364
rect -33 314 33 330
rect -15 292 15 314
rect -15 -314 15 -292
rect -33 -330 33 -314
rect -33 -364 -17 -330
rect 17 -364 33 -330
rect -33 -380 33 -364
<< polycont >>
rect -17 330 17 364
rect -17 -364 17 -330
<< locali >>
rect -175 432 -79 466
rect 79 432 175 466
rect -175 370 -141 432
rect 141 370 175 432
rect -33 330 -17 364
rect 17 330 33 364
rect -61 280 -27 296
rect -61 -296 -27 -280
rect 27 280 61 296
rect 27 -296 61 -280
rect -33 -364 -17 -330
rect 17 -364 33 -330
rect -175 -432 -141 -370
rect 141 -432 175 -370
rect -175 -466 -79 -432
rect 79 -466 175 -432
<< viali >>
rect -17 330 17 364
rect -61 -280 -27 280
rect 27 -280 61 280
rect -17 -364 17 -330
<< metal1 >>
rect -29 364 29 370
rect -29 330 -17 364
rect 17 330 29 364
rect -29 324 29 330
rect -67 280 -21 292
rect -67 -280 -61 280
rect -27 -280 -21 280
rect -67 -292 -21 -280
rect 21 280 67 292
rect 21 -280 27 280
rect 61 -280 67 280
rect 21 -292 67 -280
rect -29 -330 29 -324
rect -29 -364 -17 -330
rect 17 -364 29 -330
rect -29 -370 29 -364
<< properties >>
string FIXED_BBOX -158 -449 158 449
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.92 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
