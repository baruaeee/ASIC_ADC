** sch_path: /home/exotic/Desktop/ASIC_ADC/xschem/Vth_sch/Pre_layout/th08.sch
**.subckt th08 Vin Vout
*.ipin Vin
*.opin Vout
VDD VDD GND 1.8
Vin Vin GND pulse(0 0.2 0ns 1ns 1ns 5ns 10ns)
V_logic_high V_LH GND 1.25
V_logic_low V_LL GND 0.5
x1 VDD Vout Vin GND th08
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.save all





.dc Vin 0 1.8 0.01
*.tran 1n 30n
.control
run
set color0=white
set color1=black
plot Vin Vout V_LH V_LL
set xbrushwidth=3
.save all
.endc
.end


**** end user architecture code
**.ends

* NGSPICE file created from th08.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_LNCAWD a_n67_n130# a_n125_n42# a_67_n42# a_n227_n216#
X0 a_67_n42# a_n67_n130# a_n125_n42# a_n227_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.67
C0 a_67_n42# a_n125_n42# 0.0322f
C1 a_n67_n130# a_67_n42# 0.0112f
C2 a_n67_n130# a_n125_n42# 0.0112f
C3 a_67_n42# a_n227_n216# 0.0807f
C4 a_n125_n42# a_n227_n216# 0.0807f
C5 a_n67_n130# a_n227_n216# 0.533f
.ends

.subckt sky130_fd_pr__pfet_01v8_M6KFPY a_n73_n67# a_n33_n164# a_15_n67# w_n211_n286#
+ VSUBS
X0 a_15_n67# a_n33_n164# a_n73_n67# w_n211_n286# sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.92 as=0.194 ps=1.92 w=0.67 l=0.15
C0 w_n211_n286# a_15_n67# 0.0616f
C1 a_n73_n67# a_n33_n164# 0.0213f
C2 w_n211_n286# a_n73_n67# 0.0616f
C3 w_n211_n286# a_n33_n164# 0.238f
C4 a_15_n67# a_n73_n67# 0.11f
C5 a_15_n67# a_n33_n164# 0.0213f
C6 a_15_n67# VSUBS 0.0364f
C7 a_n73_n67# VSUBS 0.0364f
C8 a_n33_n164# VSUBS 0.116f
C9 w_n211_n286# VSUBS 1.11f
.ends

.subckt sky130_fd_pr__pfet_01v8_NZD9V2 w_n243_n261# a_47_n42# a_n47_n139# a_n105_n42#
+ VSUBS
X0 a_47_n42# a_n47_n139# a_n105_n42# w_n243_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.47
C0 w_n243_n261# a_47_n42# 0.0499f
C1 a_n105_n42# a_n47_n139# 0.00866f
C2 w_n243_n261# a_n105_n42# 0.0499f
C3 w_n243_n261# a_n47_n139# 0.27f
C4 a_47_n42# a_n105_n42# 0.0406f
C5 a_47_n42# a_n47_n139# 0.00866f
C6 a_47_n42# VSUBS 0.0297f
C7 a_n105_n42# VSUBS 0.0297f
C8 a_n47_n139# VSUBS 0.168f
C9 w_n243_n261# VSUBS 1.17f
.ends

.subckt sky130_fd_pr__nfet_01v8_NCP4B2 a_n73_n47# a_n175_n221# a_n33_n135# a_15_n47#
X0 a_15_n47# a_n33_n135# a_n73_n47# a_n175_n221# sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.52 as=0.136 ps=1.52 w=0.47 l=0.15
C0 a_15_n47# a_n73_n47# 0.0779f
C1 a_n33_n135# a_15_n47# 0.0213f
C2 a_n33_n135# a_n73_n47# 0.0213f
C3 a_15_n47# a_n175_n221# 0.0779f
C4 a_n73_n47# a_n175_n221# 0.0779f
C5 a_n33_n135# a_n175_n221# 0.338f
.ends

.subckt th08 Vp V08 Vin Vn
XXM0 Vin m1_451_n1105# Vn Vn sky130_fd_pr__nfet_01v8_LNCAWD
XXM1 m1_451_n1105# Vin Vp Vp Vn sky130_fd_pr__pfet_01v8_M6KFPY
XXM2 Vp V08 m1_451_n1105# Vp Vn sky130_fd_pr__pfet_01v8_NZD9V2
XXM3 Vn Vn m1_451_n1105# V08 sky130_fd_pr__nfet_01v8_NCP4B2
C0 Vin V08 2.59e-19
C1 V08 Vp 0.0989f
C2 m1_451_n1105# Vin 0.365f
C3 m1_451_n1105# Vp 0.176f
C4 m1_451_n1105# V08 0.175f
C5 Vin Vp 0.125f
C6 m1_451_n1105# Vn 0.838f
C7 Vp Vn 2.37f
C8 V08 Vn 0.403f
C9 Vin Vn 0.981f
.ends


.GLOBAL VDD
.GLOBAL GND
.GLOBAL V_LH
.GLOBAL V_LL
.end
