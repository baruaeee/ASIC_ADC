magic
tech sky130A
magscale 1 2
timestamp 1696186025
<< error_s >>
rect 129 1047 187 1053
rect 129 1013 141 1047
rect 129 1007 187 1013
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 1696184460
transform 1 0 158 0 1 866
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1696186025
transform 1 0 635 0 1 856
box -211 -310 211 310
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 GND
port 3 nsew
<< end >>
