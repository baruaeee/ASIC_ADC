magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_s >>
rect 362 1006 397 1024
rect 362 999 433 1006
rect 363 970 433 999
rect 380 936 451 970
rect 731 963 766 970
rect 731 936 802 963
rect 380 583 450 936
rect 732 927 802 936
rect 749 893 820 927
rect 1100 893 1135 910
rect 562 868 620 874
rect 562 834 574 868
rect 562 828 620 834
rect 562 666 620 672
rect 562 632 574 666
rect 562 626 620 632
rect 380 547 433 583
rect 749 530 819 893
rect 1101 892 1135 893
rect 1101 856 1171 892
rect 931 825 989 831
rect 931 791 943 825
rect 1118 822 1189 856
rect 931 785 989 791
rect 931 613 989 619
rect 931 579 943 613
rect 931 573 989 579
rect 749 494 802 530
rect 1118 477 1188 822
rect 1301 754 1359 760
rect 1301 720 1313 754
rect 1301 714 1359 720
rect 1301 560 1359 566
rect 1301 526 1313 560
rect 1301 520 1359 526
rect 1118 441 1171 477
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_EDPLE3  XM1
timestamp 1703732895
transform 1 0 960 0 1 702
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_VGVEGU  XM3
timestamp 1703732895
transform 1 0 1330 0 1 640
box -212 -252 212 252
use sky130_fd_pr__pfet_01v8_NZD9V2  XM7
timestamp 1703732895
transform 1 0 190 0 1 808
box -243 -261 243 261
use sky130_fd_pr__nfet_01v8_97T34Z  XM10
timestamp 1703732895
transform 1 0 591 0 1 750
box -211 -256 211 256
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
