* NGSPICE file created from analog_therm.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 w_n211_n319# a_n33_n197# 0.246f
C1 a_n73_n100# a_15_n100# 0.162f
C2 a_n33_n197# a_15_n100# 0.0262f
C3 a_n33_n197# a_n73_n100# 0.0281f
C4 w_n211_n319# a_15_n100# 0.0815f
C5 w_n211_n319# a_n73_n100# 0.0813f
C6 a_15_n100# VSUBS 0.0492f
C7 a_n73_n100# VSUBS 0.0487f
C8 a_n33_n197# VSUBS 0.129f
C9 w_n211_n319# VSUBS 1.23f
.ends

.subckt sky130_fd_pr__nfet_01v8_L7T3GD a_n33_n130# a_15_n42# a_n175_n216# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n33_n130# a_n73_n42# 0.0209f
C1 a_n73_n42# a_15_n42# 0.0699f
C2 a_n33_n130# a_15_n42# 0.0209f
C3 a_15_n42# a_n175_n216# 0.0729f
C4 a_n73_n42# a_n175_n216# 0.0729f
C5 a_n33_n130# a_n175_n216# 0.338f
.ends

.subckt sky130_fd_pr__pfet_01v8_QPDSQG a_n87_n42# w_n225_n261# a_n33_n139# a_29_n42#
+ VSUBS
X0 a_29_n42# a_n33_n139# a_n87_n42# w_n225_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.29
C0 w_n225_n261# a_n33_n139# 0.229f
C1 a_n87_n42# a_29_n42# 0.0532f
C2 a_n33_n139# a_29_n42# 0.00625f
C3 a_n33_n139# a_n87_n42# 0.00625f
C4 w_n225_n261# a_29_n42# 0.0499f
C5 w_n225_n261# a_n87_n42# 0.0499f
C6 a_29_n42# VSUBS 0.029f
C7 a_n87_n42# VSUBS 0.029f
C8 a_n33_n139# VSUBS 0.128f
C9 w_n225_n261# VSUBS 1.09f
.ends

.subckt sky130_fd_pr__pfet_01v8_M479BZ a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 w_n211_n261# a_n33_n139# 0.236f
C1 a_n73_n42# a_15_n42# 0.0699f
C2 a_n33_n139# a_15_n42# 0.0192f
C3 a_n33_n139# a_n73_n42# 0.0192f
C4 w_n211_n261# a_15_n42# 0.0463f
C5 w_n211_n261# a_n73_n42# 0.0463f
C6 a_15_n42# VSUBS 0.0263f
C7 a_n73_n42# VSUBS 0.0263f
C8 a_n33_n139# VSUBS 0.115f
C9 w_n211_n261# VSUBS 1.03f
.ends

.subckt th10 V10 Vin m1_718_n418# Vp Vn m1_878_n414#
XXM0 Vn m1_878_n414# Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vin m1_878_n414# Vn m1_718_n418# sky130_fd_pr__nfet_01v8_L7T3GD
XXM2 Vp Vp Vin m1_718_n418# Vn sky130_fd_pr__pfet_01v8_QPDSQG
XXM3 V10 Vp m1_718_n418# Vp Vn sky130_fd_pr__pfet_01v8_M479BZ
XXM4 m1_718_n418# V10 Vn Vn sky130_fd_pr__nfet_01v8_L7T3GD
C0 V10 m1_718_n418# 0.191f
C1 V10 Vin 1.33e-19
C2 Vn m1_718_n418# 0.14f
C3 Vn Vin 0.0481f
C4 Vp m1_878_n414# 0.0409f
C5 V10 m1_878_n414# 9.3e-21
C6 m1_718_n418# Vin 0.308f
C7 Vn m1_878_n414# 0.157f
C8 V10 Vp 0.0825f
C9 Vn Vp 0.468f
C10 V10 Vn 0.0667f
C11 m1_718_n418# m1_878_n414# 0.0145f
C12 Vin m1_878_n414# 0.0391f
C13 Vp m1_718_n418# 0.272f
C14 Vp Vin 0.301f
C15 m1_718_n418# 0 0.567f
C16 V10 0 0.319f
C17 Vn 0 0.208f
C18 Vp 0 3.6f
C19 Vin 0 0.692f
C20 m1_878_n414# 0 0.16f
.ends

.subckt sky130_fd_pr__pfet_01v8_FP437E w_n521_n261# a_n383_n42# a_n325_n139# a_325_n42#
+ VSUBS
X0 a_325_n42# a_n325_n139# a_n383_n42# w_n521_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.25
C0 a_n325_n139# a_n383_n42# 0.0222f
C1 a_325_n42# a_n325_n139# 0.0222f
C2 w_n521_n261# a_n383_n42# 0.0498f
C3 a_325_n42# w_n521_n261# 0.0498f
C4 a_325_n42# a_n383_n42# 0.00865f
C5 w_n521_n261# a_n325_n139# 1.13f
C6 a_325_n42# VSUBS 0.0355f
C7 a_n383_n42# VSUBS 0.0355f
C8 a_n325_n139# VSUBS 0.87f
C9 w_n521_n261# VSUBS 2.3f
.ends

.subckt preamp Vp Vn Vin Vpamp
XXM0 Vpamp Vpamp Vin Vn Vpamp sky130_fd_pr__pfet_01v8_FP437E
XXM1 Vin Vpamp Vpamp Vp sky130_fd_pr__nfet_01v8_L7T3GD
C0 Vp Vin 0.116f
C1 Vpamp Vin 0.665f
C2 Vpamp Vn 0.0667f
C3 Vpamp Vp 0.116f
C4 Vn Vin 0.0405f
C5 Vin 0 1.35f
C6 Vpamp 0 2.29f
C7 Vp 0 0.324f
C8 Vn 0 0.123f
.ends

.subckt sky130_fd_pr__pfet_01v8_NZD9V2 w_n243_n261# a_47_n42# a_n47_n139# a_n105_n42#
+ VSUBS
X0 a_47_n42# a_n47_n139# a_n105_n42# w_n243_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.47
C0 w_n243_n261# a_n47_n139# 0.27f
C1 a_n47_n139# a_n105_n42# 0.00866f
C2 w_n243_n261# a_n105_n42# 0.0499f
C3 a_47_n42# a_n47_n139# 0.00866f
C4 a_47_n42# w_n243_n261# 0.0499f
C5 a_47_n42# a_n105_n42# 0.0406f
C6 a_47_n42# VSUBS 0.0297f
C7 a_n105_n42# VSUBS 0.0297f
C8 a_n47_n139# VSUBS 0.168f
C9 w_n243_n261# VSUBS 1.17f
.ends

.subckt sky130_fd_pr__pfet_01v8_3PDS9J a_n102_n42# a_44_n42# a_n44_n139# w_n240_n261#
+ VSUBS
X0 a_44_n42# a_n44_n139# a_n102_n42# w_n240_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.44
C0 w_n240_n261# a_n44_n139# 0.261f
C1 a_n44_n139# a_n102_n42# 0.00823f
C2 w_n240_n261# a_n102_n42# 0.0499f
C3 a_44_n42# a_n44_n139# 0.00823f
C4 a_44_n42# w_n240_n261# 0.0499f
C5 a_44_n42# a_n102_n42# 0.0423f
C6 a_44_n42# VSUBS 0.0296f
C7 a_n102_n42# VSUBS 0.0296f
C8 a_n44_n139# VSUBS 0.16f
C9 w_n240_n261# VSUBS 1.15f
.ends

.subckt sky130_fd_pr__nfet_01v8_97T34Z a_n73_n46# a_n175_n220# a_n33_n134# a_15_n46#
X0 a_15_n46# a_n33_n134# a_n73_n46# a_n175_n220# sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.5 as=0.133 ps=1.5 w=0.46 l=0.15
C0 a_n33_n134# a_n73_n46# 0.0212f
C1 a_n73_n46# a_15_n46# 0.0763f
C2 a_n33_n134# a_15_n46# 0.0212f
C3 a_15_n46# a_n175_n220# 0.0769f
C4 a_n73_n46# a_n175_n220# 0.0769f
C5 a_n33_n134# a_n175_n220# 0.338f
.ends

.subckt th06 Vp Vin V06 m1_528_n874# Vn
XXM0 Vin m1_528_n874# Vn Vn sky130_fd_pr__nfet_01v8_L7T3GD
XXM1 Vp m1_528_n874# Vin Vp Vn sky130_fd_pr__pfet_01v8_NZD9V2
XXM2 Vp V06 m1_528_n874# Vp Vn sky130_fd_pr__pfet_01v8_3PDS9J
XXM3 Vn Vn m1_528_n874# V06 sky130_fd_pr__nfet_01v8_97T34Z
C0 Vin m1_528_n874# 0.224f
C1 Vin V06 2.39e-21
C2 Vp Vin 0.192f
C3 m1_528_n874# V06 0.135f
C4 Vp m1_528_n874# 0.467f
C5 Vp V06 0.109f
C6 m1_528_n874# Vn 0.971f
C7 V06 Vn 0.353f
C8 Vin Vn 0.726f
C9 Vp Vn 2.62f
.ends

.subckt sky130_fd_pr__pfet_01v8_3QB9EZ a_n296_n139# a_n354_n42# a_296_n42# w_n492_n261#
+ VSUBS
X0 a_296_n42# a_n296_n139# a_n354_n42# w_n492_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.96
C0 w_n492_n261# a_296_n42# 0.0498f
C1 w_n492_n261# a_n354_n42# 0.0498f
C2 a_n296_n139# a_296_n42# 0.0218f
C3 a_n354_n42# a_n296_n139# 0.0218f
C4 w_n492_n261# a_n296_n139# 1.04f
C5 a_n354_n42# a_296_n42# 0.00943f
C6 a_296_n42# VSUBS 0.0352f
C7 a_n354_n42# VSUBS 0.0352f
C8 a_n296_n139# VSUBS 0.797f
C9 w_n492_n261# VSUBS 2.19f
.ends

.subckt sky130_fd_pr__nfet_01v8_J2SMPG a_n33_n398# a_15_n310# a_n175_n484# a_n73_n310#
X0 a_15_n310# a_n33_n398# a_n73_n310# a_n175_n484# sky130_fd_pr__nfet_01v8 ad=0.899 pd=6.78 as=0.899 ps=6.78 w=3.1 l=0.15
C0 a_n33_n398# a_15_n310# 0.0365f
C1 a_15_n310# a_n73_n310# 0.496f
C2 a_n33_n398# a_n73_n310# 0.0365f
C3 a_15_n310# a_n175_n484# 0.345f
C4 a_n73_n310# a_n175_n484# 0.345f
C5 a_n33_n398# a_n175_n484# 0.349f
.ends

.subckt sky130_fd_pr__nfet_01v8_G45C34 a_297_n48# a_n297_n136# a_n457_n222# a_n355_n48#
X0 a_297_n48# a_n297_n136# a_n355_n48# a_n457_n222# sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.54 as=0.139 ps=1.54 w=0.48 l=2.97
C0 a_n297_n136# a_297_n48# 0.0239f
C1 a_297_n48# a_n355_n48# 0.0107f
C2 a_n297_n136# a_n355_n48# 0.0239f
C3 a_297_n48# a_n457_n222# 0.0929f
C4 a_n355_n48# a_n457_n222# 0.0929f
C5 a_n297_n136# a_n457_n222# 1.8f
.ends

.subckt sky130_fd_pr__pfet_01v8_XA2NHL a_15_n310# w_n211_n529# a_n73_n310# a_n33_n407#
+ VSUBS
X0 a_15_n310# a_n33_n407# a_n73_n310# w_n211_n529# sky130_fd_pr__pfet_01v8 ad=0.899 pd=6.78 as=0.899 ps=6.78 w=3.1 l=0.15
C0 w_n211_n529# a_15_n310# 0.21f
C1 w_n211_n529# a_n73_n310# 0.21f
C2 a_n33_n407# a_15_n310# 0.0346f
C3 a_n73_n310# a_n33_n407# 0.0346f
C4 w_n211_n529# a_n33_n407# 0.241f
C5 a_n73_n310# a_15_n310# 0.496f
C6 a_15_n310# VSUBS 0.135f
C7 a_n73_n310# VSUBS 0.135f
C8 a_n33_n407# VSUBS 0.121f
C9 w_n211_n529# VSUBS 1.97f
.ends

.subckt th01 Vin Vout m1_931_n929# Vp Vn
XXM2 Vin Vp m1_931_n929# Vp Vn sky130_fd_pr__pfet_01v8_3QB9EZ
XXM3 Vin m1_931_n929# Vn Vn sky130_fd_pr__nfet_01v8_J2SMPG
XXM4 Vn m1_931_n929# Vn Vout sky130_fd_pr__nfet_01v8_G45C34
XXM5 Vp Vp Vout m1_931_n929# Vn sky130_fd_pr__pfet_01v8_XA2NHL
C0 m1_931_n929# Vout 0.202f
C1 Vp Vout 0.0877f
C2 Vp m1_931_n929# 0.324f
C3 Vin Vout 5.64e-20
C4 m1_931_n929# Vin 0.206f
C5 Vp Vin 0.391f
C6 Vin Vn 1.12f
C7 Vout Vn 0.405f
C8 m1_931_n929# Vn 2.31f
C9 Vp Vn 4.35f
.ends

.subckt sky130_fd_pr__nfet_01v8_VGVEGU a_n74_n42# a_n33_n130# a_n176_n216# a_16_n42#
X0 a_16_n42# a_n33_n130# a_n74_n42# a_n176_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.16
C0 a_16_n42# a_n33_n130# 0.0191f
C1 a_n74_n42# a_n33_n130# 0.0191f
C2 a_n74_n42# a_16_n42# 0.0684f
C3 a_16_n42# a_n176_n216# 0.0737f
C4 a_n74_n42# a_n176_n216# 0.0737f
C5 a_n33_n130# a_n176_n216# 0.338f
.ends

.subckt sky130_fd_pr__pfet_01v8_EDPLE3 a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n42# w_n211_n261# 0.0463f
C1 a_n33_n139# w_n211_n261# 0.236f
C2 a_15_n42# w_n211_n261# 0.0463f
C3 a_n33_n139# a_n73_n42# 0.0192f
C4 a_15_n42# a_n73_n42# 0.0699f
C5 a_n33_n139# a_15_n42# 0.0192f
C6 a_15_n42# VSUBS 0.0263f
C7 a_n73_n42# VSUBS 0.0263f
C8 a_n33_n139# VSUBS 0.115f
C9 w_n211_n261# VSUBS 1.03f
.ends

.subckt th07 Vp Vin V07 m1_400_n1066# Vn
XXM0 m1_400_n1066# Vin Vn Vn sky130_fd_pr__nfet_01v8_VGVEGU
XXM1 m1_400_n1066# Vp Vin Vp Vn sky130_fd_pr__pfet_01v8_EDPLE3
XXM2 Vp V07 m1_400_n1066# Vp Vn sky130_fd_pr__pfet_01v8_NZD9V2
XXM3 Vn Vn m1_400_n1066# V07 sky130_fd_pr__nfet_01v8_97T34Z
C0 Vp V07 0.102f
C1 m1_400_n1066# Vin 0.436f
C2 V07 Vin 6.52e-19
C3 m1_400_n1066# V07 0.167f
C4 Vp Vin 0.212f
C5 Vp m1_400_n1066# 0.32f
C6 Vin Vn 0.75f
C7 m1_400_n1066# Vn 0.943f
C8 V07 Vn 0.395f
C9 Vp Vn 2.43f
.ends

.subckt sky130_fd_pr__nfet_01v8_LNCAWD a_n67_n130# a_n125_n42# a_67_n42# a_n227_n216#
X0 a_67_n42# a_n67_n130# a_n125_n42# a_n227_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.67
C0 a_n125_n42# a_n67_n130# 0.0112f
C1 a_n67_n130# a_67_n42# 0.0112f
C2 a_n125_n42# a_67_n42# 0.0322f
C3 a_67_n42# a_n227_n216# 0.0807f
C4 a_n125_n42# a_n227_n216# 0.0807f
C5 a_n67_n130# a_n227_n216# 0.533f
.ends

.subckt sky130_fd_pr__pfet_01v8_M6KFPY a_n73_n67# a_n33_n164# a_15_n67# w_n211_n286#
+ VSUBS
X0 a_15_n67# a_n33_n164# a_n73_n67# w_n211_n286# sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.92 as=0.194 ps=1.92 w=0.67 l=0.15
C0 a_n33_n164# w_n211_n286# 0.238f
C1 a_n73_n67# a_15_n67# 0.11f
C2 w_n211_n286# a_15_n67# 0.0616f
C3 w_n211_n286# a_n73_n67# 0.0616f
C4 a_n33_n164# a_15_n67# 0.0213f
C5 a_n33_n164# a_n73_n67# 0.0213f
C6 a_15_n67# VSUBS 0.0364f
C7 a_n73_n67# VSUBS 0.0364f
C8 a_n33_n164# VSUBS 0.116f
C9 w_n211_n286# VSUBS 1.11f
.ends

.subckt sky130_fd_pr__nfet_01v8_NCP4B2 a_n73_n47# a_n175_n221# a_n33_n135# a_15_n47#
X0 a_15_n47# a_n33_n135# a_n73_n47# a_n175_n221# sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.52 as=0.136 ps=1.52 w=0.47 l=0.15
C0 a_n73_n47# a_n33_n135# 0.0213f
C1 a_n33_n135# a_15_n47# 0.0213f
C2 a_n73_n47# a_15_n47# 0.0779f
C3 a_15_n47# a_n175_n221# 0.0779f
C4 a_n73_n47# a_n175_n221# 0.0779f
C5 a_n33_n135# a_n175_n221# 0.338f
.ends

.subckt th08 Vp V08 Vin m1_451_n1105# Vn
XXM0 Vin m1_451_n1105# Vn Vn sky130_fd_pr__nfet_01v8_LNCAWD
XXM1 m1_451_n1105# Vin Vp Vp Vn sky130_fd_pr__pfet_01v8_M6KFPY
XXM2 Vp V08 m1_451_n1105# Vp Vn sky130_fd_pr__pfet_01v8_NZD9V2
XXM3 Vn Vn m1_451_n1105# V08 sky130_fd_pr__nfet_01v8_NCP4B2
C0 Vp Vin 0.125f
C1 Vin m1_451_n1105# 0.365f
C2 Vp V08 0.0989f
C3 m1_451_n1105# V08 0.175f
C4 Vin V08 2.59e-19
C5 Vp m1_451_n1105# 0.176f
C6 m1_451_n1105# Vn 0.838f
C7 Vin Vn 0.981f
C8 Vp Vn 2.37f
C9 V08 Vn 0.403f
.ends

.subckt sky130_fd_pr__nfet_01v8_JLSX9N a_n317_n216# a_n157_n130# a_n215_n42# a_157_n42#
X0 a_157_n42# a_n157_n130# a_n215_n42# a_n317_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.57
C0 a_n215_n42# a_n157_n130# 0.0179f
C1 a_157_n42# a_n215_n42# 0.0166f
C2 a_157_n42# a_n157_n130# 0.0179f
C3 a_157_n42# a_n317_n216# 0.0832f
C4 a_n215_n42# a_n317_n216# 0.0832f
C5 a_n157_n130# a_n317_n216# 1.03f
.ends

.subckt sky130_fd_pr__pfet_01v8_XYZSMQ a_n33_n255# a_15_n158# w_n211_n377# a_n73_n158#
+ VSUBS
X0 a_15_n158# a_n33_n255# a_n73_n158# w_n211_n377# sky130_fd_pr__pfet_01v8 ad=0.458 pd=3.74 as=0.458 ps=3.74 w=1.58 l=0.15
C0 a_n33_n255# w_n211_n377# 0.24f
C1 a_15_n158# a_n33_n255# 0.0271f
C2 a_n73_n158# a_n33_n255# 0.0271f
C3 a_15_n158# w_n211_n377# 0.117f
C4 a_n73_n158# w_n211_n377# 0.117f
C5 a_n73_n158# a_15_n158# 0.254f
C6 a_15_n158# VSUBS 0.0732f
C7 a_n73_n158# VSUBS 0.0732f
C8 a_n33_n255# VSUBS 0.118f
C9 w_n211_n377# VSUBS 1.43f
.ends

.subckt sky130_fd_pr__pfet_01v8_AZD9DW w_n353_n261# a_n157_n139# a_n215_n42# a_157_n42#
+ VSUBS
X0 a_157_n42# a_n157_n139# a_n215_n42# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.57
C0 a_n157_n139# w_n353_n261# 0.611f
C1 a_157_n42# a_n157_n139# 0.0179f
C2 a_n215_n42# a_n157_n139# 0.0179f
C3 a_157_n42# w_n353_n261# 0.0498f
C4 a_n215_n42# w_n353_n261# 0.0498f
C5 a_n215_n42# a_157_n42# 0.0166f
C6 a_157_n42# VSUBS 0.0329f
C7 a_n215_n42# VSUBS 0.0329f
C8 a_n157_n139# VSUBS 0.446f
C9 w_n353_n261# VSUBS 1.62f
.ends

.subckt sky130_fd_pr__nfet_01v8_T8HSQ7 a_15_n157# a_n175_n331# a_n33_n245# a_n73_n157#
X0 a_15_n157# a_n33_n245# a_n73_n157# a_n175_n331# sky130_fd_pr__nfet_01v8 ad=0.455 pd=3.72 as=0.455 ps=3.72 w=1.57 l=0.15
C0 a_n73_n157# a_n33_n245# 0.0289f
C1 a_15_n157# a_n73_n157# 0.253f
C2 a_15_n157# a_n33_n245# 0.0289f
C3 a_15_n157# a_n175_n331# 0.19f
C4 a_n73_n157# a_n175_n331# 0.19f
C5 a_n33_n245# a_n175_n331# 0.346f
.ends

.subckt th09 V09 Vin m1_891_n977# Vp m1_1725_85# Vn
XXM0 Vn Vin Vn m1_891_n977# sky130_fd_pr__nfet_01v8_JLSX9N
XXM1 Vin Vp Vp m1_891_n977# Vn sky130_fd_pr__pfet_01v8_XYZSMQ
XXM2 Vp m1_891_n977# Vp m1_1725_85# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM3 Vp m1_891_n977# V09 m1_1725_85# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM4 V09 Vn m1_891_n977# Vn sky130_fd_pr__nfet_01v8_T8HSQ7
C0 Vin Vp 0.162f
C1 Vp m1_1725_85# 0.14f
C2 m1_891_n977# V09 0.291f
C3 Vin m1_1725_85# 9.1e-19
C4 m1_891_n977# Vp 0.469f
C5 Vp V09 0.131f
C6 m1_891_n977# Vin 0.208f
C7 m1_891_n977# m1_1725_85# 0.0672f
C8 Vin V09 0.00135f
C9 V09 m1_1725_85# 0.0153f
C10 Vin Vn 1.36f
C11 m1_891_n977# Vn 1.29f
C12 V09 Vn 0.467f
C13 Vp Vn 4.41f
C14 m1_1725_85# Vn 0.13f
.ends

.subckt sky130_fd_pr__pfet_01v8_P28Q2U a_n33_n232# a_15_n135# w_n211_n354# a_n73_n135#
+ VSUBS
X0 a_15_n135# a_n33_n232# a_n73_n135# w_n211_n354# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.28 as=0.391 ps=3.28 w=1.35 l=0.15
C0 a_n73_n135# w_n211_n354# 0.103f
C1 a_n73_n135# a_15_n135# 0.218f
C2 a_n33_n232# w_n211_n354# 0.24f
C3 a_n33_n232# a_15_n135# 0.0258f
C4 a_n73_n135# a_n33_n232# 0.0258f
C5 w_n211_n354# a_15_n135# 0.103f
C6 a_15_n135# VSUBS 0.0639f
C7 a_n73_n135# VSUBS 0.0639f
C8 a_n33_n232# VSUBS 0.118f
C9 w_n211_n354# VSUBS 1.35f
.ends

.subckt sky130_fd_pr__nfet_01v8_HZA4VB a_n360_n216# a_n200_n130# a_200_n42# a_n258_n42#
X0 a_200_n42# a_n200_n130# a_n258_n42# a_n360_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_200_n42# a_n200_n130# 0.0196f
C1 a_n258_n42# a_n200_n130# 0.0196f
C2 a_200_n42# a_n258_n42# 0.0134f
C3 a_200_n42# a_n360_n216# 0.0841f
C4 a_n258_n42# a_n360_n216# 0.0841f
C5 a_n200_n130# a_n360_n216# 1.26f
.ends

.subckt sky130_fd_pr__pfet_01v8_WV9GCW a_n158_n42# w_n296_n261# a_n100_n139# a_100_n42#
+ VSUBS
X0 a_100_n42# a_n100_n139# a_n158_n42# w_n296_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1
C0 a_n158_n42# w_n296_n261# 0.0499f
C1 a_n158_n42# a_100_n42# 0.024f
C2 a_n100_n139# w_n296_n261# 0.434f
C3 a_n100_n139# a_100_n42# 0.0144f
C4 a_n158_n42# a_n100_n139# 0.0144f
C5 w_n296_n261# a_100_n42# 0.0499f
C6 a_100_n42# VSUBS 0.0315f
C7 a_n158_n42# VSUBS 0.0315f
C8 a_n100_n139# VSUBS 0.302f
C9 w_n296_n261# VSUBS 1.38f
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_15_n100# a_n33_n188# 0.0254f
C1 a_n73_n100# a_n33_n188# 0.0254f
C2 a_15_n100# a_n73_n100# 0.162f
C3 a_15_n100# a_n175_n274# 0.132f
C4 a_n73_n100# a_n175_n274# 0.132f
C5 a_n33_n188# a_n175_n274# 0.343f
.ends

.subckt th12 Vout Vin m1_532_n361# Vp m1_773_n853# Vn
XXM0 Vn m1_773_n853# Vp Vn Vn sky130_fd_pr__pfet_01v8_P28Q2U
XXM1 Vn Vin m1_773_n853# m1_532_n361# sky130_fd_pr__nfet_01v8_HZA4VB
XXM2 m1_532_n361# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM3 Vp Vp m1_532_n361# Vout Vn sky130_fd_pr__pfet_01v8_WV9GCW
XXM4 Vn m1_532_n361# Vout Vn sky130_fd_pr__nfet_01v8_648S5X
C0 Vin m1_532_n361# 0.399f
C1 Vin Vout 4.83e-19
C2 m1_773_n853# m1_532_n361# 0.0208f
C3 m1_773_n853# Vout 0.00284f
C4 Vin Vp 0.434f
C5 Vout m1_532_n361# 0.181f
C6 m1_773_n853# Vp 0.0827f
C7 Vp m1_532_n361# 0.225f
C8 Vin m1_773_n853# 0.102f
C9 Vout Vp 0.0968f
C10 m1_532_n361# Vn 1.04f
C11 Vout Vn 0.478f
C12 Vin Vn 1.62f
C13 Vp Vn 4.59f
C14 m1_773_n853# Vn 0.44f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGAKDL a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
+ VSUBS
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n73_n200# w_n211_n419# 0.143f
C1 a_n73_n200# a_n33_n297# 0.0293f
C2 a_n73_n200# a_15_n200# 0.321f
C3 a_n33_n297# w_n211_n419# 0.24f
C4 w_n211_n419# a_15_n200# 0.143f
C5 a_n33_n297# a_15_n200# 0.0293f
C6 a_15_n200# VSUBS 0.0902f
C7 a_n73_n200# VSUBS 0.0902f
C8 a_n33_n297# VSUBS 0.119f
C9 w_n211_n419# VSUBS 1.58f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFH27D a_50_n42# a_n210_n216# a_n108_n42# a_n50_n130#
X0 a_50_n42# a_n50_n130# a_n108_n42# a_n210_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 a_50_n42# a_n50_n130# 0.00909f
C1 a_50_n42# a_n108_n42# 0.0391f
C2 a_n108_n42# a_n50_n130# 0.00909f
C3 a_50_n42# a_n210_n216# 0.0801f
C4 a_n108_n42# a_n210_n216# 0.0801f
C5 a_n50_n130# a_n210_n216# 0.439f
.ends

.subckt sky130_fd_pr__pfet_01v8_E7ZT25 a_15_n43# w_n211_n262# a_n73_n43# a_n33_n140#
+ VSUBS
X0 a_15_n43# a_n33_n140# a_n73_n43# w_n211_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.15
C0 a_n73_n43# w_n211_n262# 0.0469f
C1 a_n73_n43# a_n33_n140# 0.0193f
C2 a_n73_n43# a_15_n43# 0.0715f
C3 a_n33_n140# w_n211_n262# 0.236f
C4 w_n211_n262# a_15_n43# 0.0469f
C5 a_n33_n140# a_15_n43# 0.0193f
C6 a_15_n43# VSUBS 0.0267f
C7 a_n73_n43# VSUBS 0.0267f
C8 a_n33_n140# VSUBS 0.115f
C9 w_n211_n262# VSUBS 1.03f
.ends

.subckt sky130_fd_pr__pfet_01v8_JM8GTH a_50_n42# w_n246_n261# a_n50_n139# a_n108_n42#
+ VSUBS
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 a_n108_n42# w_n246_n261# 0.0499f
C1 a_n108_n42# a_n50_n139# 0.00909f
C2 a_n108_n42# a_50_n42# 0.0391f
C3 a_n50_n139# w_n246_n261# 0.279f
C4 w_n246_n261# a_50_n42# 0.0499f
C5 a_n50_n139# a_50_n42# 0.00909f
C6 a_50_n42# VSUBS 0.0298f
C7 a_n108_n42# VSUBS 0.0298f
C8 a_n50_n139# VSUBS 0.175f
C9 w_n246_n261# VSUBS 1.18f
.ends

.subckt sky130_fd_pr__nfet_01v8_L9ESAD a_n175_n224# a_n73_n50# a_n33_n138# a_15_n50#
X0 a_15_n50# a_n33_n138# a_n73_n50# a_n175_n224# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_15_n50# a_n33_n138# 0.0216f
C1 a_15_n50# a_n73_n50# 0.0826f
C2 a_n73_n50# a_n33_n138# 0.0216f
C3 a_15_n50# a_n175_n224# 0.081f
C4 a_n73_n50# a_n175_n224# 0.081f
C5 a_n33_n138# a_n175_n224# 0.339f
.ends

.subckt th11 V11 Vin m1_717_301# m1_509_303# Vp Vn
XXM0 m1_717_301# Vp Vn Vn Vn sky130_fd_pr__pfet_01v8_XGAKDL
XXM1 m1_717_301# Vn m1_509_303# Vin sky130_fd_pr__nfet_01v8_ZFH27D
XXM2 m1_509_303# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_E7ZT25
XXM3 V11 Vp m1_509_303# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM4 Vn Vn m1_509_303# V11 sky130_fd_pr__nfet_01v8_L9ESAD
C0 Vin Vp 0.258f
C1 m1_509_303# Vin 0.248f
C2 m1_717_301# V11 1.71e-20
C3 m1_509_303# Vp 0.352f
C4 m1_717_301# Vin 0.0345f
C5 m1_717_301# Vp 0.0487f
C6 m1_717_301# m1_509_303# 0.0301f
C7 Vin V11 0.00112f
C8 V11 Vp 0.0686f
C9 m1_509_303# V11 0.0742f
C10 Vin Vn 0.856f
C11 m1_509_303# Vn 0.717f
C12 V11 Vn 0.485f
C13 Vp Vn 4.47f
C14 m1_717_301# Vn 0.299f
.ends

.subckt sky130_fd_pr__nfet_01v8_L6G859 a_n288_n42# a_230_n42# a_n390_n216# a_n230_n130#
X0 a_230_n42# a_n230_n130# a_n288_n42# a_n390_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.3
C0 a_n230_n130# a_230_n42# 0.0204f
C1 a_n230_n130# a_n288_n42# 0.0204f
C2 a_230_n42# a_n288_n42# 0.0119f
C3 a_230_n42# a_n390_n216# 0.0846f
C4 a_n288_n42# a_n390_n216# 0.0846f
C5 a_n230_n130# a_n390_n216# 1.43f
.ends

.subckt sky130_fd_pr__pfet_01v8_XW9KDL a_n73_n230# a_n33_n327# a_15_n230# w_n211_n449#
+ VSUBS
X0 a_15_n230# a_n33_n327# a_n73_n230# w_n211_n449# sky130_fd_pr__pfet_01v8 ad=0.667 pd=5.18 as=0.667 ps=5.18 w=2.3 l=0.15
C0 a_15_n230# w_n211_n449# 0.161f
C1 w_n211_n449# a_n73_n230# 0.161f
C2 a_15_n230# a_n73_n230# 0.369f
C3 w_n211_n449# a_n33_n327# 0.246f
C4 a_15_n230# a_n33_n327# 0.0338f
C5 a_n73_n230# a_n33_n327# 0.0338f
C6 a_15_n230# VSUBS 0.102f
C7 a_n73_n230# VSUBS 0.102f
C8 a_n33_n327# VSUBS 0.129f
C9 w_n211_n449# VSUBS 1.69f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GC6 a_200_n42# w_n396_n261# a_n200_n139# a_n258_n42#
+ VSUBS
X0 a_200_n42# a_n200_n139# a_n258_n42# w_n396_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_200_n42# w_n396_n261# 0.0498f
C1 w_n396_n261# a_n258_n42# 0.0498f
C2 a_200_n42# a_n258_n42# 0.0134f
C3 w_n396_n261# a_n200_n139# 0.743f
C4 a_200_n42# a_n200_n139# 0.0196f
C5 a_n258_n42# a_n200_n139# 0.0196f
C6 a_200_n42# VSUBS 0.0338f
C7 a_n258_n42# VSUBS 0.0338f
C8 a_n200_n139# VSUBS 0.554f
C9 w_n396_n261# VSUBS 1.79f
.ends

.subckt sky130_fd_pr__nfet_01v8_ATLS57 a_15_n200# a_n175_n374# a_n73_n200# a_n33_n288#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n175_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n33_n288# a_15_n200# 0.0357f
C1 a_n33_n288# a_n73_n200# 0.0336f
C2 a_15_n200# a_n73_n200# 0.321f
C3 a_15_n200# a_n175_n374# 0.232f
C4 a_n73_n200# a_n175_n374# 0.232f
C5 a_n33_n288# a_n175_n374# 0.358f
.ends

.subckt th13 Vout Vin m1_724_n958# m1_546_n454# Vp Vn
XXM0 m1_724_n958# Vn Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 m1_546_n454# m1_724_n958# Vn Vin sky130_fd_pr__nfet_01v8_L6G859
XXM2 m1_546_n454# Vin Vp Vp Vn sky130_fd_pr__pfet_01v8_XW9KDL
XXM3 Vout Vp m1_546_n454# Vp Vn sky130_fd_pr__pfet_01v8_VZ9GC6
XXM4 Vout Vn Vn m1_546_n454# sky130_fd_pr__nfet_01v8_ATLS57
C0 Vp m1_546_n454# 0.574f
C1 m1_724_n958# Vp 0.312f
C2 m1_546_n454# Vin 0.349f
C3 m1_724_n958# Vin 0.14f
C4 m1_724_n958# m1_546_n454# 0.0214f
C5 Vp Vn 0.589f
C6 Vin Vn 0.126f
C7 m1_546_n454# Vn 0.331f
C8 m1_724_n958# Vn 0.0967f
C9 Vp Vout 0.346f
C10 Vout Vin 0.00172f
C11 Vout m1_546_n454# 0.546f
C12 m1_724_n958# Vout 0.00247f
C13 Vout Vn 0.147f
C14 Vp Vin 0.151f
C15 Vout 0 0.513f
C16 Vn 0 0.573f
C17 m1_546_n454# 0 1.54f
C18 Vp 0 4.74f
C19 Vin 0 1.66f
C20 m1_724_n958# 0 0.188f
.ends

.subckt sky130_fd_pr__nfet_01v8_9GNSAK a_n33_n550# a_n125_n550# a_n227_n724# a_63_n550#
+ a_n63_n576#
X0 a_63_n550# a_n63_n576# a_n33_n550# a_n227_n724# sky130_fd_pr__nfet_01v8 ad=1.71 pd=11.6 as=0.908 ps=5.83 w=5.5 l=0.15
X1 a_n33_n550# a_n63_n576# a_n125_n550# a_n227_n724# sky130_fd_pr__nfet_01v8 ad=0.908 pd=5.83 as=1.71 ps=11.6 w=5.5 l=0.15
C0 a_63_n550# a_n63_n576# 0.0319f
C1 a_63_n550# a_n33_n550# 0.809f
C2 a_n63_n576# a_n33_n550# 0.0599f
C3 a_n125_n550# a_n63_n576# 0.0232f
C4 a_n125_n550# a_n33_n550# 0.809f
C5 a_63_n550# a_n227_n724# 0.596f
C6 a_n33_n550# a_n227_n724# 0.0778f
C7 a_n125_n550# a_n227_n724# 0.597f
C8 a_n63_n576# a_n227_n724# 0.3f
.ends

.subckt sky130_fd_pr__pfet_01v8_UTD9YE w_n1296_n261# a_n1158_n42# a_n1100_n139# a_1100_n42#
+ VSUBS
X0 a_1100_n42# a_n1100_n139# a_n1158_n42# w_n1296_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=11
C0 a_1100_n42# w_n1296_n261# 0.0498f
C1 w_n1296_n261# a_n1158_n42# 0.0498f
C2 a_n1100_n139# a_1100_n42# 0.0251f
C3 a_n1100_n139# w_n1296_n261# 3.52f
C4 a_n1100_n139# a_n1158_n42# 0.0251f
C5 a_1100_n42# VSUBS 0.0428f
C6 a_n1158_n42# VSUBS 0.0428f
C7 a_n1100_n139# VSUBS 2.83f
C8 w_n1296_n261# VSUBS 5.47f
.ends

.subckt sky130_fd_pr__nfet_01v8_VZ7MP4 a_n1158_n42# a_n1260_n216# a_n1100_n130# a_1100_n42#
X0 a_1100_n42# a_n1100_n130# a_n1158_n42# a_n1260_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=11
C0 a_n1100_n130# a_1100_n42# 0.0251f
C1 a_n1158_n42# a_n1100_n130# 0.0251f
C2 a_1100_n42# a_n1260_n216# 0.0931f
C3 a_n1158_n42# a_n1260_n216# 0.0931f
C4 a_n1100_n130# a_n1260_n216# 6.21f
.ends

.subckt sky130_fd_pr__pfet_01v8_UGSTRG a_n33_n1197# a_n76_n1100# w_n214_n1319# a_18_n1100#
+ VSUBS
X0 a_18_n1100# a_n33_n1197# a_n76_n1100# w_n214_n1319# sky130_fd_pr__pfet_01v8 ad=3.19 pd=22.6 as=3.19 ps=22.6 w=11 l=0.18
C0 a_18_n1100# w_n214_n1319# 0.693f
C1 a_18_n1100# a_n76_n1100# 1.64f
C2 w_n214_n1319# a_n76_n1100# 0.693f
C3 a_n33_n1197# a_18_n1100# 0.0705f
C4 a_n33_n1197# w_n214_n1319# 0.239f
C5 a_n33_n1197# a_n76_n1100# 0.0705f
C6 a_18_n1100# VSUBS 0.46f
C7 a_n76_n1100# VSUBS 0.46f
C8 a_n33_n1197# VSUBS 0.133f
C9 w_n214_n1319# VSUBS 4.79f
.ends

.subckt th02 Vp Vn m1_4146_502# Vin Vout m1_1199_9#
XXM0 Vn m1_4146_502# Vn m1_4146_502# Vin sky130_fd_pr__nfet_01v8_9GNSAK
XXM1 Vp m1_1199_9# Vin m1_4146_502# Vn sky130_fd_pr__pfet_01v8_UTD9YE
XXM2 m1_1199_9# Vn Vp Vp sky130_fd_pr__nfet_01v8_VZ7MP4
XXM3 m1_4146_502# Vout Vp Vp Vn sky130_fd_pr__pfet_01v8_UGSTRG
XXM4 Vn Vn m1_4146_502# Vout sky130_fd_pr__nfet_01v8_VZ7MP4
C0 Vin m1_1199_9# 0.0993f
C1 Vin m1_4146_502# 0.58f
C2 m1_4146_502# m1_1199_9# 4.98e-19
C3 Vp Vout 0.202f
C4 Vin Vp 0.3f
C5 Vin Vout 0.0111f
C6 Vp m1_1199_9# 0.155f
C7 Vp m1_4146_502# 0.374f
C8 m1_4146_502# Vout 0.328f
C9 m1_4146_502# Vn 9.06f
C10 Vout Vn 0.554f
C11 m1_1199_9# Vn 0.445f
C12 Vp Vn 16.7f
C13 Vin Vn 2.92f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJ7SDL a_15_n450# w_n211_n669# a_n73_n450# a_n33_n547#
+ VSUBS
X0 a_15_n450# a_n33_n547# a_n73_n450# w_n211_n669# sky130_fd_pr__pfet_01v8 ad=1.3 pd=9.58 as=1.3 ps=9.58 w=4.5 l=0.15
C0 a_15_n450# w_n211_n669# 0.295f
C1 a_n73_n450# w_n211_n669# 0.295f
C2 w_n211_n669# a_n33_n547# 0.242f
C3 a_n73_n450# a_15_n450# 0.718f
C4 a_15_n450# a_n33_n547# 0.0407f
C5 a_n73_n450# a_n33_n547# 0.0407f
C6 a_15_n450# VSUBS 0.191f
C7 a_n73_n450# VSUBS 0.191f
C8 a_n33_n547# VSUBS 0.122f
C9 w_n211_n669# VSUBS 2.46f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFMUVB a_n608_n42# a_550_n42# a_n710_n216# a_n550_n130#
X0 a_550_n42# a_n550_n130# a_n608_n42# a_n710_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=5.5
C0 a_550_n42# a_n550_n130# 0.0242f
C1 a_n550_n130# a_n608_n42# 0.0242f
C2 a_550_n42# a_n608_n42# 0.00526f
C3 a_550_n42# a_n710_n216# 0.0873f
C4 a_n608_n42# a_n710_n216# 0.0873f
C5 a_n550_n130# a_n710_n216# 3.19f
.ends

.subckt sky130_fd_pr__pfet_01v8_UJPVTG w_n211_n769# a_n73_n550# a_n33_n647# a_15_n550#
+ VSUBS
X0 a_15_n550# a_n33_n647# a_n73_n550# w_n211_n769# sky130_fd_pr__pfet_01v8 ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.15
C0 a_15_n550# w_n211_n769# 0.356f
C1 a_n73_n550# w_n211_n769# 0.356f
C2 w_n211_n769# a_n33_n647# 0.242f
C3 a_n73_n550# a_15_n550# 0.877f
C4 a_15_n550# a_n33_n647# 0.0449f
C5 a_n73_n550# a_n33_n647# 0.0449f
C6 a_15_n550# VSUBS 0.232f
C7 a_n73_n550# VSUBS 0.232f
C8 a_n33_n647# VSUBS 0.122f
C9 w_n211_n769# VSUBS 2.81f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GTR a_n608_n42# a_550_n42# w_n746_n261# a_n550_n139#
+ VSUBS
X0 a_550_n42# a_n550_n139# a_n608_n42# w_n746_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=5.5
C0 a_550_n42# w_n746_n261# 0.0498f
C1 a_n608_n42# w_n746_n261# 0.0498f
C2 w_n746_n261# a_n550_n139# 1.82f
C3 a_n608_n42# a_550_n42# 0.00526f
C4 a_550_n42# a_n550_n139# 0.0242f
C5 a_n608_n42# a_n550_n139# 0.0242f
C6 a_550_n42# VSUBS 0.037f
C7 a_n608_n42# VSUBS 0.037f
C8 a_n550_n139# VSUBS 1.44f
C9 w_n746_n261# VSUBS 3.22f
.ends

.subckt sky130_fd_pr__nfet_01v8_9GNSAM a_n73_n550# a_n175_n724# a_15_n550# a_n33_n638#
X0 a_15_n550# a_n33_n638# a_n73_n550# a_n175_n724# sky130_fd_pr__nfet_01v8 ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.15
C0 a_15_n550# a_n33_n638# 0.0468f
C1 a_n33_n638# a_n73_n550# 0.0468f
C2 a_15_n550# a_n73_n550# 0.877f
C3 a_15_n550# a_n175_n724# 0.588f
C4 a_n73_n550# a_n175_n724# 0.588f
C5 a_n33_n638# a_n175_n724# 0.352f
.ends

.subckt th14 Vout Vin m1_1594_n962# Vp m1_710_n388# m1_2498_n384# Vn
XXM0 m1_1594_n962# Vp Vn Vn Vn sky130_fd_pr__pfet_01v8_XJ7SDL
XXM1 m1_710_n388# m1_1594_n962# Vn Vin sky130_fd_pr__nfet_01v8_ZFMUVB
XXM2 Vp m1_710_n388# Vin Vp Vn sky130_fd_pr__pfet_01v8_UJPVTG
XXM3 Vp m1_2498_n384# Vp m1_710_n388# Vn sky130_fd_pr__pfet_01v8_VZ9GTR
XXM4 m1_2498_n384# Vout Vp m1_710_n388# Vn sky130_fd_pr__pfet_01v8_VZ9GTR
XXM5 Vn Vn Vout m1_710_n388# sky130_fd_pr__nfet_01v8_9GNSAM
C0 Vp m1_2498_n384# 0.276f
C1 m1_1594_n962# m1_710_n388# 0.00647f
C2 Vout m1_2498_n384# 0.0142f
C3 m1_1594_n962# Vin 0.166f
C4 Vp Vout 0.125f
C5 m1_1594_n962# Vn 0.111f
C6 m1_2498_n384# m1_710_n388# 0.768f
C7 Vin m1_2498_n384# 1.46e-19
C8 Vp m1_710_n388# 0.755f
C9 m1_2498_n384# Vn 3.34e-24
C10 Vin Vp 0.214f
C11 Vp Vn 0.876f
C12 Vout m1_710_n388# 0.191f
C13 Vout Vn 0.0354f
C14 Vin m1_710_n388# 0.365f
C15 m1_1594_n962# Vp 0.237f
C16 m1_710_n388# Vn 0.459f
C17 Vin Vn 0.0583f
C18 Vin 0 3.4f
C19 Vout 0 0.854f
C20 Vn 0 0.831f
C21 m1_710_n388# 0 3.52f
C22 m1_2498_n384# 0 0.297f
C23 Vp 0 11.9f
C24 m1_1594_n962# 0 0.292f
.ends

.subckt sky130_fd_pr__nfet_01v8_8X7S4D a_15_n130# a_n33_n218# a_n73_n130# a_n175_n304#
X0 a_15_n130# a_n33_n218# a_n73_n130# a_n175_n304# sky130_fd_pr__nfet_01v8 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=0.15
C0 a_n33_n218# a_15_n130# 0.0274f
C1 a_n73_n130# a_15_n130# 0.21f
C2 a_n73_n130# a_n33_n218# 0.0274f
C3 a_15_n130# a_n175_n304# 0.162f
C4 a_n73_n130# a_n175_n304# 0.162f
C5 a_n33_n218# a_n175_n304# 0.345f
.ends

.subckt sky130_fd_pr__pfet_01v8_GZD9X3 a_n139_n139# a_139_n42# w_n335_n261# a_n197_n42#
+ VSUBS
X0 a_139_n42# a_n139_n139# a_n197_n42# w_n335_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.39
C0 a_139_n42# w_n335_n261# 0.0498f
C1 w_n335_n261# a_n197_n42# 0.0498f
C2 a_n139_n139# a_139_n42# 0.017f
C3 a_n139_n139# a_n197_n42# 0.017f
C4 a_n139_n139# w_n335_n261# 0.555f
C5 a_139_n42# a_n197_n42# 0.0184f
C6 a_139_n42# VSUBS 0.0325f
C7 a_n197_n42# VSUBS 0.0325f
C8 a_n139_n139# VSUBS 0.4f
C9 w_n335_n261# VSUBS 1.54f
.ends

.subckt sky130_fd_pr__nfet_01v8_LH5FDA a_n310_n216# a_n150_n130# a_n208_n42# a_150_n42#
X0 a_150_n42# a_n150_n130# a_n208_n42# a_n310_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.5
C0 a_n150_n130# a_150_n42# 0.0176f
C1 a_n208_n42# a_150_n42# 0.0172f
C2 a_n208_n42# a_n150_n130# 0.0176f
C3 a_150_n42# a_n310_n216# 0.0831f
C4 a_n208_n42# a_n310_n216# 0.0831f
C5 a_n150_n130# a_n310_n216# 0.99f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJP3BL a_15_n150# w_n211_n369# a_n73_n150# a_n33_n247#
+ VSUBS
X0 a_15_n150# a_n33_n247# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.15
C0 a_15_n150# w_n211_n369# 0.112f
C1 w_n211_n369# a_n73_n150# 0.112f
C2 a_n33_n247# a_15_n150# 0.0267f
C3 a_n33_n247# a_n73_n150# 0.0267f
C4 a_n33_n247# w_n211_n369# 0.24f
C5 a_15_n150# a_n73_n150# 0.242f
C6 a_15_n150# VSUBS 0.07f
C7 a_n73_n150# VSUBS 0.07f
C8 a_n33_n247# VSUBS 0.118f
C9 w_n211_n369# VSUBS 1.41f
.ends

.subckt th03 Vp Vout Vin m1_522_n210# li_1010_10# m1_782_n682# Vn
XXM0 m1_782_n682# Vin Vn Vn sky130_fd_pr__nfet_01v8_8X7S4D
XXM1 Vin m1_782_n682# li_1010_10# m1_522_n210# Vn sky130_fd_pr__pfet_01v8_GZD9X3
XXM2 Vn Vp m1_522_n210# Vp sky130_fd_pr__nfet_01v8_LH5FDA
XXM3 Vout li_1010_10# Vp m1_782_n682# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 Vn m1_782_n682# Vn Vout sky130_fd_pr__nfet_01v8_LH5FDA
C0 m1_522_n210# Vin 0.0482f
C1 m1_522_n210# m1_782_n682# 0.0254f
C2 m1_522_n210# li_1010_10# 0.0635f
C3 Vin m1_782_n682# 0.212f
C4 li_1010_10# Vin 0.0791f
C5 li_1010_10# m1_782_n682# 0.263f
C6 m1_522_n210# Vout 0.00126f
C7 Vin Vout 5.05e-19
C8 m1_782_n682# Vout 0.0652f
C9 li_1010_10# Vout 0.132f
C10 m1_522_n210# Vp 0.041f
C11 Vin Vp 0.0439f
C12 Vp m1_782_n682# 0.143f
C13 li_1010_10# Vp 0.0961f
C14 Vp Vout 3.29e-19
C15 Vout Vn 0.462f
C16 m1_782_n682# Vn 1.57f
C17 Vp Vn 1.26f
C18 m1_522_n210# Vn 0.278f
C19 Vin Vn 0.853f
C20 li_1010_10# Vn 3.06f
.ends

.subckt sky130_fd_pr__pfet_01v8_MYW2PY a_n73_n48# a_n33_n145# a_15_n48# w_n211_n267#
+ VSUBS
X0 a_15_n48# a_n33_n145# a_n73_n48# w_n211_n267# sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.54 as=0.139 ps=1.54 w=0.48 l=0.15
C0 a_n33_n145# w_n211_n267# 0.237f
C1 a_15_n48# w_n211_n267# 0.05f
C2 a_n73_n48# w_n211_n267# 0.05f
C3 a_15_n48# a_n33_n145# 0.0197f
C4 a_n33_n145# a_n73_n48# 0.0197f
C5 a_15_n48# a_n73_n48# 0.0795f
C6 a_15_n48# VSUBS 0.0287f
C7 a_n73_n48# VSUBS 0.0287f
C8 a_n33_n145# VSUBS 0.115f
C9 w_n211_n267# VSUBS 1.05f
.ends

.subckt sky130_fd_pr__nfet_01v8_JRGCPP a_n1108_n42# a_1050_n42# a_n1210_n216# a_n1050_n130#
X0 a_1050_n42# a_n1050_n130# a_n1108_n42# a_n1210_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=10.5
C0 a_n1108_n42# a_n1050_n130# 0.0251f
C1 a_1050_n42# a_n1050_n130# 0.0251f
C2 a_1050_n42# a_n1210_n216# 0.0931f
C3 a_n1108_n42# a_n1210_n216# 0.0931f
C4 a_n1050_n130# a_n1210_n216# 5.94f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJ78MR a_n73_n1050# w_n211_n1269# a_15_n1050# a_n33_n1147#
+ VSUBS
X0 a_15_n1050# a_n33_n1147# a_n73_n1050# w_n211_n1269# sky130_fd_pr__pfet_01v8 ad=3.05 pd=21.6 as=3.05 ps=21.6 w=10.5 l=0.15
C0 a_n33_n1147# w_n211_n1269# 0.242f
C1 a_15_n1050# w_n211_n1269# 0.661f
C2 a_n73_n1050# w_n211_n1269# 0.661f
C3 a_15_n1050# a_n33_n1147# 0.065f
C4 a_n33_n1147# a_n73_n1050# 0.065f
C5 a_15_n1050# a_n73_n1050# 1.67f
C6 a_15_n1050# VSUBS 0.434f
C7 a_n73_n1050# VSUBS 0.434f
C8 a_n33_n1147# VSUBS 0.129f
C9 w_n211_n1269# VSUBS 4.56f
.ends

.subckt sky130_fd_pr__pfet_01v8_6M437L a_n1108_n42# a_1050_n42# a_n1050_n139# w_n1246_n261#
+ VSUBS
X0 a_1050_n42# a_n1050_n139# a_n1108_n42# w_n1246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=10.5
C0 a_n1050_n139# w_n1246_n261# 3.36f
C1 a_1050_n42# w_n1246_n261# 0.0498f
C2 a_n1108_n42# w_n1246_n261# 0.0498f
C3 a_1050_n42# a_n1050_n139# 0.0251f
C4 a_n1050_n139# a_n1108_n42# 0.0251f
C5 a_1050_n42# VSUBS 0.0428f
C6 a_n1108_n42# VSUBS 0.0428f
C7 a_n1050_n139# VSUBS 2.7f
C8 w_n1246_n261# VSUBS 5.27f
.ends

.subckt sky130_fd_pr__nfet_01v8_A5ES5P a_n73_n1000# a_15_n1000# a_n33_n1088# a_n175_n1174#
X0 a_15_n1000# a_n33_n1088# a_n73_n1000# a_n175_n1174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.6 as=2.9 ps=20.6 w=10 l=0.15
C0 a_n73_n1000# a_n33_n1088# 0.0649f
C1 a_15_n1000# a_n33_n1088# 0.0649f
C2 a_n73_n1000# a_15_n1000# 1.59f
C3 a_15_n1000# a_n175_n1174# 1.04f
C4 a_n73_n1000# a_n175_n1174# 1.04f
C5 a_n33_n1088# a_n175_n1174# 0.359f
.ends

.subckt th15 m1_1074_6# m1_915_n714# Vp m1_4024_602# Vin Vout Vn m1_1076_814#
XXM0 m1_915_n714# Vn Vn Vp Vn sky130_fd_pr__pfet_01v8_MYW2PY
XXM1 m1_1074_6# m1_915_n714# Vn Vin sky130_fd_pr__nfet_01v8_JRGCPP
XXM2 m1_1076_814# m1_1074_6# Vn Vin sky130_fd_pr__nfet_01v8_JRGCPP
XXM3 m1_1076_814# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_XJ78MR
XXM4 Vp m1_4024_602# m1_1076_814# Vp Vn sky130_fd_pr__pfet_01v8_6M437L
XXM5 Vn Vout m1_1076_814# Vn sky130_fd_pr__nfet_01v8_A5ES5P
XXM7 m1_4024_602# Vout m1_1076_814# Vp Vn sky130_fd_pr__pfet_01v8_6M437L
C0 m1_1076_814# m1_4024_602# 0.999f
C1 m1_1076_814# m1_1074_6# 0.0103f
C2 m1_4024_602# Vin 1.79e-19
C3 m1_1076_814# Vout 0.214f
C4 m1_915_n714# Vp 0.596f
C5 m1_1074_6# Vin 1.03f
C6 m1_1076_814# Vin 0.6f
C7 m1_4024_602# Vp 0.404f
C8 m1_1074_6# m1_915_n714# 0.0137f
C9 m1_1074_6# Vp 0.0774f
C10 m1_1076_814# m1_915_n714# 3.02e-20
C11 Vout Vp 0.129f
C12 m1_1076_814# Vp 1.22f
C13 Vin m1_915_n714# 0.378f
C14 Vin Vp 0.222f
C15 m1_4024_602# Vout 0.00816f
C16 m1_4024_602# Vn 0.411f
C17 Vout Vn 1.46f
C18 m1_1076_814# Vn 6.13f
C19 Vin Vn 11.5f
C20 Vp Vn 18.4f
C21 m1_1074_6# Vn 0.844f
C22 m1_915_n714# Vn 1.17f
.ends

.subckt sky130_fd_pr__nfet_01v8_42G4RD a_n80_n42# a_n33_n130# a_n182_n216# a_22_n42#
X0 a_22_n42# a_n33_n130# a_n80_n42# a_n182_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_n33_n130# a_22_n42# 0.00866f
C1 a_n33_n130# a_n80_n42# 0.00866f
C2 a_n80_n42# a_22_n42# 0.0604f
C3 a_22_n42# a_n182_n216# 0.0785f
C4 a_n80_n42# a_n182_n216# 0.0785f
C5 a_n33_n130# a_n182_n216# 0.341f
.ends

.subckt sky130_fd_pr__pfet_01v8_DDPLQ8 a_n77_n42# w_n215_n261# a_n33_n139# a_19_n42#
+ VSUBS
X0 a_19_n42# a_n33_n139# a_n77_n42# w_n215_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 w_n215_n261# a_n77_n42# 0.0484f
C1 w_n215_n261# a_19_n42# 0.0484f
C2 a_n77_n42# a_19_n42# 0.0641f
C3 w_n215_n261# a_n33_n139# 0.234f
C4 a_n33_n139# a_n77_n42# 0.0127f
C5 a_n33_n139# a_19_n42# 0.0127f
C6 a_19_n42# VSUBS 0.0275f
C7 a_n77_n42# VSUBS 0.0275f
C8 a_n33_n139# VSUBS 0.119f
C9 w_n215_n261# VSUBS 1.04f
.ends

.subckt sky130_fd_pr__nfet_01v8_VWP3K3 a_n33_n130# a_15_n42# a_n175_n216# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n33_n130# a_15_n42# 0.0209f
C1 a_n33_n130# a_n73_n42# 0.0209f
C2 a_n73_n42# a_15_n42# 0.0699f
C3 a_15_n42# a_n175_n216# 0.0729f
C4 a_n73_n42# a_n175_n216# 0.0729f
C5 a_n33_n130# a_n175_n216# 0.338f
.ends

.subckt sky130_fd_pr__pfet_01v8_LZD9A4 a_n80_n42# a_22_n42# a_n33_n139# w_n218_n261#
+ VSUBS
X0 a_22_n42# a_n33_n139# a_n80_n42# w_n218_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 w_n218_n261# a_n80_n42# 0.0496f
C1 w_n218_n261# a_22_n42# 0.0496f
C2 a_n80_n42# a_22_n42# 0.0604f
C3 w_n218_n261# a_n33_n139# 0.233f
C4 a_n33_n139# a_n80_n42# 0.0084f
C5 a_n33_n139# a_22_n42# 0.0084f
C6 a_22_n42# VSUBS 0.0285f
C7 a_n80_n42# VSUBS 0.0285f
C8 a_n33_n139# VSUBS 0.122f
C9 w_n218_n261# VSUBS 1.06f
.ends

.subckt sky130_fd_pr__nfet_01v8_VRD6K3 a_n77_n42# a_n33_n130# a_19_n42# a_n179_n216#
X0 a_19_n42# a_n33_n130# a_n77_n42# a_n179_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_n33_n130# a_19_n42# 0.0136f
C1 a_n33_n130# a_n77_n42# 0.0136f
C2 a_n77_n42# a_19_n42# 0.0641f
C3 a_19_n42# a_n179_n216# 0.0763f
C4 a_n77_n42# a_n179_n216# 0.0763f
C5 a_n33_n130# a_n179_n216# 0.339f
.ends

.subckt th04 Vp V04 Vin Vn m1_960_n972# m1_397_n357#
XXM0 m1_960_n972# Vin Vn Vn sky130_fd_pr__nfet_01v8_42G4RD
XXM1 m1_397_n357# Vp Vin m1_960_n972# Vn sky130_fd_pr__pfet_01v8_DDPLQ8
XXM2 Vp m1_397_n357# Vn Vp sky130_fd_pr__nfet_01v8_VWP3K3
XXM3 Vp V04 m1_960_n972# Vp Vn sky130_fd_pr__pfet_01v8_LZD9A4
XXM4 V04 m1_960_n972# Vn Vn sky130_fd_pr__nfet_01v8_VRD6K3
C0 V04 Vn 0.181f
C1 Vp m1_960_n972# 0.257f
C2 Vp V04 0.173f
C3 m1_960_n972# V04 0.39f
C4 Vin Vn 0.0911f
C5 m1_397_n357# Vn 0.0588f
C6 Vin Vp 0.103f
C7 Vp m1_397_n357# 0.401f
C8 Vin m1_960_n972# 0.395f
C9 m1_960_n972# m1_397_n357# 0.027f
C10 Vin V04 5.12e-19
C11 V04 m1_397_n357# 0.0695f
C12 Vp Vn 0.228f
C13 Vin m1_397_n357# 0.109f
C14 m1_960_n972# Vn 0.346f
C15 Vin 0 0.599f
C16 Vn 0 0.213f
C17 V04 0 0.324f
C18 m1_960_n972# 0 0.53f
C19 Vp 0 2.61f
C20 m1_397_n357# 0 0.189f
.ends

.subckt sky130_fd_pr__pfet_01v8_PZD9SE a_n112_n139# w_n308_n261# a_112_n42# a_n170_n42#
+ VSUBS
X0 a_112_n42# a_n112_n139# a_n170_n42# w_n308_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.12
C0 a_n112_n139# a_112_n42# 0.0153f
C1 a_n170_n42# a_112_n42# 0.0219f
C2 a_n112_n139# w_n308_n261# 0.472f
C3 a_n170_n42# w_n308_n261# 0.0499f
C4 a_n170_n42# a_n112_n139# 0.0153f
C5 a_112_n42# w_n308_n261# 0.0499f
C6 a_112_n42# VSUBS 0.0318f
C7 a_n170_n42# VSUBS 0.0318f
C8 a_n112_n139# VSUBS 0.332f
C9 w_n308_n261# VSUBS 1.43f
.ends

.subckt sky130_fd_pr__nfet_01v8_UNLS3X a_n33_n200# a_n175_n286# a_n73_n112# a_15_n112#
X0 a_15_n112# a_n33_n200# a_n73_n112# a_n175_n286# sky130_fd_pr__nfet_01v8 ad=0.325 pd=2.82 as=0.325 ps=2.82 w=1.12 l=0.15
C0 a_n73_n112# a_n33_n200# 0.0262f
C1 a_15_n112# a_n33_n200# 0.0262f
C2 a_15_n112# a_n73_n112# 0.181f
C3 a_15_n112# a_n175_n286# 0.144f
C4 a_n73_n112# a_n175_n286# 0.144f
C5 a_n33_n200# a_n175_n286# 0.344f
.ends

.subckt th05 V05 Vin m1_836_n724# Vp Vn
XXM0 m1_836_n724# Vn Vn Vin sky130_fd_pr__nfet_01v8_ATLS57
XXM1 m1_836_n724# Vp Vin Vp Vn sky130_fd_pr__pfet_01v8_VZ9GC6
XXM2 m1_836_n724# Vp V05 Vp Vn sky130_fd_pr__pfet_01v8_PZD9SE
XXM3 m1_836_n724# Vn Vn V05 sky130_fd_pr__nfet_01v8_UNLS3X
C0 Vin m1_836_n724# 0.185f
C1 m1_836_n724# Vp 0.372f
C2 Vin V05 5.09e-20
C3 V05 Vp 0.103f
C4 V05 m1_836_n724# 0.122f
C5 Vin Vp 0.324f
C6 V05 Vn 0.48f
C7 m1_836_n724# Vn 1.23f
C8 Vin Vn 1.06f
C9 Vp Vn 3.53f
.ends

.subckt Analog Vin Vp V1 V2 V3 V4 V5 V6 V7 V8 V10 V11 V12 V13 V14 V15 x28/m1_1594_n962#
+ x29/m1_1074_6# x31/Vp x22/m1_451_n1105# x18/Vin x29/m1_915_n714# x28/m1_710_n388#
+ x28/m1_2498_n384# x21/m1_400_n1066# x27/m1_724_n958# x26/m1_532_n361# x30/Vin x31/m1_931_n929#
+ x25/m1_717_301# th10_0/m1_718_n418# x28/Vin x16/m1_1199_9# x17/m1_522_n210# x26/m1_773_n853#
+ x17/li_1010_10# x25/Vin x16/m1_4146_502# x31/Vin x19/m1_836_n724# x20/m1_528_n874#
+ x23/m1_891_n977# x23/m1_1725_85# x16/Vin x27/m1_546_n454# x28/Vp x25/m1_509_303#
+ x21/Vp x20/Vp x29/Vp x22/Vp x17/m1_782_n682# V9 x29/Vin x22/Vin x18/m1_960_n972#
+ x18/m1_397_n357# Vn x29/m1_1076_814#
Xth10_0 V10 x29/Vin th10_0/m1_718_n418# x29/Vp Vn th10_0/m1_878_n414# th10
Xx30 Vp Vn x30/Vin Vn preamp
Xx20 x20/Vp x29/Vin V6 x20/m1_528_n874# Vn th06
Xx31 x31/Vin V1 x31/m1_931_n929# x31/Vp Vn th01
Xx21 x21/Vp x22/Vin V7 x21/m1_400_n1066# Vn th07
Xx22 x22/Vp V8 x22/Vin x22/m1_451_n1105# Vn th08
Xx23 V9 x29/Vin x23/m1_891_n977# x29/Vp x23/m1_1725_85# Vn th09
Xx26 V12 x29/Vin x26/m1_532_n361# x29/Vp x26/m1_773_n853# Vn th12
Xx25 V11 x25/Vin x25/m1_717_301# x25/m1_509_303# x31/Vp Vn th11
Xx27 V13 x29/Vin x27/m1_724_n958# x27/m1_546_n454# x29/Vp Vn th13
Xx16 x22/Vp Vn x16/m1_4146_502# x16/Vin V2 x16/m1_1199_9# th02
Xx28 V14 x28/Vin x28/m1_1594_n962# x28/Vp x28/m1_710_n388# x28/m1_2498_n384# Vn th14
Xx17 x22/Vp V3 x22/Vin x17/m1_522_n210# x17/li_1010_10# x17/m1_782_n682# Vn th03
Xx29 x29/m1_1074_6# x29/m1_915_n714# x29/Vp x29/m1_4024_602# x29/Vin V15 Vn x29/m1_1076_814#
+ th15
Xx18 x21/Vp V4 x18/Vin Vn x18/m1_960_n972# x18/m1_397_n357# th04
Xx19 V5 x29/Vin x19/m1_836_n724# x21/Vp Vn th05
C0 x22/Vp x16/m1_4146_502# -1.82e-19
C1 x29/Vin x29/m1_1076_814# 0.00331f
C2 x17/li_1010_10# x21/Vp 0.0158f
C3 x17/m1_782_n682# x17/li_1010_10# -1.47e-20
C4 V11 Vp 0.00915f
C5 x31/Vp x22/Vp 0.0045f
C6 x29/Vp th10_0/m1_878_n414# -2.84e-32
C7 x25/m1_717_301# x28/m1_710_n388# 1.28e-19
C8 x25/m1_509_303# V14 1.33e-19
C9 Vp x28/Vin 0.00131f
C10 x29/Vp x23/m1_891_n977# 0.0859f
C11 x18/m1_397_n357# V4 0.022f
C12 V1 x16/m1_1199_9# 1.25e-19
C13 x29/Vp x23/m1_1725_85# 0.0391f
C14 th10_0/m1_718_n418# x29/Vin 0.0103f
C15 x26/m1_532_n361# V10 8.3e-20
C16 x25/Vin x30/Vin 4.83e-19
C17 x23/m1_891_n977# V13 4e-19
C18 x26/m1_532_n361# x28/m1_710_n388# 1.26e-19
C19 x25/Vin x31/Vp 0.026f
C20 V1 x21/Vp 0.0434f
C21 x22/m1_451_n1105# x21/m1_400_n1066# 1.61e-19
C22 x23/m1_1725_85# V13 0.00456f
C23 V12 th10_0/m1_878_n414# 0.00992f
C24 x30/Vin x31/Vin 0.0267f
C25 x30/Vin x28/m1_1594_n962# 2.36e-19
C26 x17/m1_522_n210# x21/Vp 5.03e-19
C27 x31/Vp x31/Vin 3.55e-33
C28 x28/m1_710_n388# Vin 0.129f
C29 x21/m1_400_n1066# x22/Vp 3.67e-19
C30 x29/Vp x29/m1_1076_814# 0.399f
C31 x27/m1_724_n958# x27/m1_546_n454# -1.78e-33
C32 x29/Vin V10 2.18e-19
C33 x22/m1_451_n1105# x22/Vin 0.0151f
C34 x28/m1_710_n388# V14 -0.0187f
C35 x16/Vin x18/Vin 0.0107f
C36 x22/m1_451_n1105# V3 5.41e-20
C37 x25/m1_509_303# x30/Vin 0.00124f
C38 V2 x21/Vp 0.00647f
C39 V2 x17/m1_782_n682# 4.43e-20
C40 x29/Vin x28/m1_710_n388# 5.33e-19
C41 x25/m1_509_303# x31/Vp 0.00104f
C42 x25/m1_717_301# x21/Vp 0.00195f
C43 V13 x29/m1_1076_814# 0.00417f
C44 x16/Vin x31/Vp 1.59e-19
C45 x25/Vin V11 1.83e-21
C46 x29/Vin x20/Vp 0.438f
C47 x22/Vin x22/Vp 0.758f
C48 x22/Vp V3 0.0193f
C49 x21/Vp x16/m1_1199_9# 0.00199f
C50 x25/Vin x31/m1_931_n929# 0.00324f
C51 th10_0/m1_718_n418# x29/Vp -9.36e-19
C52 x26/m1_773_n853# x28/m1_710_n388# 5.73e-19
C53 V12 x28/m1_2498_n384# 0.00326f
C54 x25/Vin x18/m1_960_n972# 5.32e-20
C55 x28/Vp Vp 0.0178f
C56 x17/m1_782_n682# x21/Vp 0.0136f
C57 V14 x16/m1_1199_9# 0.00263f
C58 x18/Vin V1 0.00384f
C59 x16/m1_4146_502# V1 2.15e-20
C60 x20/Vp V8 1.02e-19
C61 x22/m1_451_n1105# x19/m1_836_n724# 8.82e-19
C62 x29/m1_915_n714# V15 0.00975f
C63 x25/m1_509_303# V11 0.00328f
C64 x29/Vp V10 0.00886f
C65 x31/Vp V1 0.0513f
C66 x25/m1_509_303# x31/m1_931_n929# 0.00234f
C67 x31/Vp x28/m1_710_n388# 0.00517f
C68 th10_0/m1_718_n418# V12 0.00398f
C69 x29/Vp x28/m1_710_n388# 0.0173f
C70 x26/m1_532_n361# x29/Vin 0.00817f
C71 x29/Vin x21/Vp 2.17e-20
C72 V9 x29/Vin 0.0119f
C73 x29/Vin x29/m1_1074_6# 2.58e-21
C74 x25/Vin V4 0.0128f
C75 V2 x16/m1_4146_502# 3.84e-19
C76 V14 Vin 0.0451f
C77 x27/m1_724_n958# x29/m1_1076_814# 3.1e-21
C78 x25/m1_717_301# x18/Vin 5.7e-19
C79 x16/Vin x22/Vin 0.321f
C80 V6 x20/Vp 0.177f
C81 x27/m1_546_n454# V15 0.0292f
C82 x30/Vin x25/m1_717_301# 8.88e-22
C83 x31/Vp x25/m1_717_301# 1.95e-21
C84 x22/Vin x17/li_1010_10# 0.138f
C85 V3 x17/li_1010_10# 0.0054f
C86 V12 V10 0.00496f
C87 V11 V1 7.8e-20
C88 V11 x28/m1_710_n388# 0.00221f
C89 V8 x21/Vp 0.00539f
C90 V8 x17/m1_782_n682# 2.02e-20
C91 V12 x28/m1_710_n388# 0.0691f
C92 V15 x29/m1_4024_602# 0.00128f
C93 x31/Vp x16/m1_1199_9# 0.0078f
C94 x31/m1_931_n929# V1 0.00621f
C95 x18/Vin x21/Vp 0.623f
C96 x25/Vin x28/Vp 1.11e-20
C97 x20/m1_528_n874# x20/Vp 0.00483f
C98 x16/m1_4146_502# x21/Vp 0.149f
C99 x16/m1_4146_502# x17/m1_782_n682# 3.69e-20
C100 x16/Vin V4 0.00227f
C101 x28/m1_710_n388# x28/Vin -1.14e-31
C102 x26/m1_773_n853# x29/Vin 4.94e-20
C103 x18/m1_960_n972# V1 0.00115f
C104 x29/Vp x26/m1_532_n361# 0.0456f
C105 x31/Vp x21/Vp 0.0365f
C106 x27/m1_546_n454# x23/m1_891_n977# 0.00379f
C107 x22/Vin V1 0.00133f
C108 x29/Vin V8 0.025f
C109 x29/Vp V9 0.136f
C110 x29/Vp x29/m1_1074_6# 9.16e-21
C111 x27/m1_546_n454# x23/m1_1725_85# 0.0174f
C112 x22/m1_451_n1105# x22/Vp 5.61e-19
C113 V6 x21/Vp 0.00284f
C114 x22/Vin x20/Vp 6.55e-22
C115 x23/m1_891_n977# x29/m1_4024_602# 0.0148f
C116 V7 x21/Vp 0.119f
C117 V7 x17/m1_782_n682# 1.9e-19
C118 x22/Vin x17/m1_522_n210# 0.0362f
C119 x31/Vp V14 5.21e-19
C120 V3 x17/m1_522_n210# 4.11e-20
C121 V5 x21/Vp 0.152f
C122 x25/m1_509_303# x28/Vp 8.44e-19
C123 x23/m1_1725_85# x29/m1_4024_602# 0.00675f
C124 th10_0/m1_718_n418# x29/m1_915_n714# 4.43e-20
C125 x29/Vp x29/Vin 1.43f
C126 x28/Vp th10_0/m1_718_n418# 1.38e-19
C127 x28/m1_1594_n962# Vp 9.76e-21
C128 V2 x22/Vin 0.0874f
C129 V4 V1 0.0394f
C130 x26/m1_532_n361# V12 0.00828f
C131 V11 x21/Vp 7.54e-19
C132 x27/m1_546_n454# x29/m1_1076_814# 0.0017f
C133 x22/Vin x25/m1_717_301# 9.98e-19
C134 V6 x29/Vin 0.0604f
C135 V15 x29/m1_1076_814# 0.141f
C136 x29/Vin V13 -6.2e-24
C137 x21/m1_400_n1066# x21/Vp 0.0408f
C138 x25/m1_509_303# Vp 6.8e-22
C139 x21/m1_400_n1066# x17/m1_782_n682# 6.38e-19
C140 x26/m1_532_n361# x28/Vin 9.23e-19
C141 x31/m1_931_n929# x21/Vp 0.0348f
C142 x29/Vp x26/m1_773_n853# 4.78e-21
C143 x29/Vin V5 2.3e-19
C144 x22/Vin x16/m1_1199_9# 0.00742f
C145 x25/Vin x22/Vp 6.33e-20
C146 x18/Vin x16/m1_4146_502# 0.0268f
C147 V12 Vin 7.02e-20
C148 x18/m1_960_n972# x21/Vp 0.00822f
C149 V10 x29/m1_915_n714# 6.77e-20
C150 V12 V14 3.02e-19
C151 x28/Vp V10 4.43e-19
C152 x20/m1_528_n874# x29/Vin 0.185f
C153 x22/Vin x21/Vp 0.05f
C154 x25/m1_717_301# V4 9.85e-19
C155 V3 x21/Vp 0.00124f
C156 x31/Vp x18/Vin 0.00447f
C157 x22/Vin x17/m1_782_n682# 0.047f
C158 V12 x29/Vin 0.162f
C159 V3 x17/m1_782_n682# 9.85e-20
C160 x28/Vp x28/m1_710_n388# -8.06e-19
C161 x30/Vin x31/Vp 0.0933f
C162 V8 V7 8.93e-20
C163 x23/m1_891_n977# x29/m1_1076_814# 0.0101f
C164 x22/m1_451_n1105# x17/li_1010_10# 4.52e-19
C165 V12 x26/m1_773_n853# 0.00206f
C166 x16/Vin x22/Vp 0.00242f
C167 x22/Vin x29/Vin 2.33e-20
C168 V4 x21/Vp 0.115f
C169 Vp x28/m1_710_n388# 2.22e-19
C170 x26/m1_773_n853# x28/Vin 7.5e-20
C171 x20/m1_528_n874# V8 6.6e-19
C172 x29/Vp V13 0.043f
C173 x22/Vp x17/li_1010_10# 0.0552f
C174 x21/m1_400_n1066# V8 3.49e-19
C175 x27/m1_724_n958# x29/Vin 0.0129f
C176 V11 x30/Vin 1.58e-20
C177 x18/m1_397_n357# x21/Vp 0.0192f
C178 x19/m1_836_n724# x21/Vp 0.0587f
C179 x18/Vin x31/m1_931_n929# 0.0043f
C180 V11 x31/Vp 0.00627f
C181 V7 V5 0.00153f
C182 x25/m1_509_303# x28/m1_2498_n384# 1.35e-20
C183 x29/Vp V12 0.114f
C184 x30/Vin x28/Vin 0.0145f
C185 x18/Vin x18/m1_960_n972# 0.00786f
C186 x18/m1_960_n972# x16/m1_4146_502# 3.43e-21
C187 x22/Vin V8 0.00574f
C188 x28/Vp x26/m1_532_n361# 2.6e-19
C189 x31/Vp x31/m1_931_n929# 0.00777f
C190 x31/Vp x28/Vin 4.25e-20
C191 x20/m1_528_n874# V6 0.0133f
C192 x29/Vp x28/Vin 0.00251f
C193 x22/Vin x18/Vin 0.0834f
C194 th10_0/m1_878_n414# x28/m1_710_n388# 3.97e-19
C195 x22/Vp V1 8.51e-19
C196 x22/Vin x16/m1_4146_502# 0.33f
C197 x31/Vp x18/m1_960_n972# 0.00118f
C198 x19/m1_836_n724# x29/Vin 0.00308f
C199 x20/m1_528_n874# V5 6e-22
C200 x28/Vp Vin 0.0147f
C201 x21/m1_400_n1066# V7 0.00217f
C202 x20/Vp x22/Vp 0.00715f
C203 x31/Vp x22/Vin 0.00882f
C204 x21/m1_400_n1066# V5 0.00268f
C205 x22/Vp x17/m1_522_n210# 0.0741f
C206 x28/Vp V14 -0.00226f
C207 x29/Vin x29/m1_915_n714# 0.114f
C208 x28/Vp x29/Vin 0.009f
C209 x25/Vin V1 0.0347f
C210 x18/Vin V4 0.0762f
C211 V2 x22/Vp 2.75e-19
C212 x16/m1_4146_502# V4 0.0145f
C213 x25/Vin x28/m1_710_n388# 6.17e-21
C214 x29/Vp x27/m1_724_n958# 0.00496f
C215 V11 x31/m1_931_n929# 8.75e-20
C216 x27/m1_546_n454# V9 0.0146f
C217 x22/Vin V7 0.00537f
C218 x25/m1_717_301# x22/Vp 5.8e-21
C219 x22/Vin V5 5.41e-20
C220 V12 x28/Vin 6.97e-21
C221 V15 x29/m1_1074_6# 7.92e-19
C222 x19/m1_836_n724# V8 0.00357f
C223 x31/Vp V4 0.00202f
C224 x18/Vin x18/m1_397_n357# 0.0184f
C225 x31/Vin V1 0.00156f
C226 x22/m1_451_n1105# x21/Vp 0.00105f
C227 x18/m1_397_n357# x16/m1_4146_502# 4.46e-19
C228 x22/m1_451_n1105# x17/m1_782_n682# 6.22e-19
C229 V9 x29/m1_4024_602# 0.00322f
C230 x28/m1_1594_n962# x28/m1_710_n388# -4.44e-34
C231 x18/m1_960_n972# x31/m1_931_n929# 0.00772f
C232 x27/m1_546_n454# x29/Vin -1.44e-19
C233 x26/m1_532_n361# th10_0/m1_878_n414# 0.00271f
C234 x22/Vin x21/m1_400_n1066# 0.0142f
C235 x21/m1_400_n1066# V3 1.89e-20
C236 x22/Vin x31/m1_931_n929# 1.71e-19
C237 x29/Vin V15 0.014f
C238 x25/m1_509_303# V1 4.21e-19
C239 x22/Vp x21/Vp 0.0571f
C240 x22/Vp x17/m1_782_n682# 0.00703f
C241 x25/m1_509_303# x28/m1_710_n388# 0.00174f
C242 x16/Vin V1 0.0131f
C243 th10_0/m1_718_n418# V10 0.00117f
C244 x28/Vp x30/Vin 0.0107f
C245 x25/Vin x16/m1_1199_9# 0.0182f
C246 x23/m1_891_n977# V9 0.00936f
C247 x22/m1_451_n1105# x29/Vin 0.00163f
C248 V6 x19/m1_836_n724# 2.76e-20
C249 th10_0/m1_718_n418# x28/m1_710_n388# 6.85e-19
C250 x28/Vp x31/Vp 0.00232f
C251 x29/Vp x29/m1_915_n714# 0.0172f
C252 x28/Vp x29/Vp 0.0763f
C253 V9 x23/m1_1725_85# 2.2e-19
C254 x22/Vin V3 0.108f
C255 x16/Vin x17/m1_522_n210# 6.18e-20
C256 x19/m1_836_n724# V5 0.00145f
C257 x22/Vp V14 0.00387f
C258 x29/Vin th10_0/m1_878_n414# 8.04e-21
C259 x31/m1_931_n929# V4 0.0179f
C260 x25/Vin x21/Vp 0.038f
C261 x29/Vin x22/Vp 0.0103f
C262 V2 x16/Vin 7.03e-21
C263 x30/Vin Vp 0.00278f
C264 x23/m1_891_n977# x29/Vin 0.0167f
C265 x20/m1_528_n874# x19/m1_836_n724# 4.81e-19
C266 x18/m1_960_n972# V4 1.63e-19
C267 x31/Vp Vp 0.00201f
C268 x23/m1_1725_85# x29/Vin 3.1e-19
C269 x22/m1_451_n1105# V8 0.00689f
C270 V10 x28/m1_710_n388# 2.86e-19
C271 x18/m1_397_n357# x31/m1_931_n929# 1.34e-21
C272 x22/Vin V4 0.00364f
C273 x31/Vin x21/Vp 3.58e-20
C274 x25/Vin V14 4.91e-21
C275 x29/Vp x27/m1_546_n454# 0.102f
C276 x28/Vp V11 5.16e-20
C277 x29/Vp V15 0.162f
C278 x28/Vp V12 0.0719f
C279 V8 x22/Vp 0.0495f
C280 x25/m1_509_303# x21/Vp 0.00381f
C281 x22/Vin x19/m1_836_n724# 8.82e-20
C282 x27/m1_546_n454# V13 0.014f
C283 x16/Vin x21/Vp 0.013f
C284 x28/Vp x28/Vin 5.68e-32
C285 x29/Vp x29/m1_4024_602# 0.0314f
C286 th10_0/m1_718_n418# x26/m1_532_n361# 2.18e-19
C287 V13 V15 0.0168f
C288 Vin Vn 0.2f
C289 V5 Vn 0.441f
C290 x19/m1_836_n724# Vn 1.04f
C291 x29/Vin Vn 25.5f
C292 x18/Vin Vn 1.51f
C293 V4 Vn 0.578f
C294 x18/m1_960_n972# Vn 0.533f
C295 x18/m1_397_n357# Vn 0.192f
C296 x29/m1_4024_602# Vn 0.411f
C297 V15 Vn 2.77f
C298 x29/m1_1076_814# Vn 5.99f
C299 x29/m1_1074_6# Vn 0.643f
C300 x29/m1_915_n714# Vn 0.87f
C301 V3 Vn 0.549f
C302 x17/m1_782_n682# Vn 1.49f
C303 x17/m1_522_n210# Vn 0.24f
C304 x17/li_1010_10# Vn 2.84f
C305 x28/Vin Vn 3.41f
C306 V14 Vn 0.852f
C307 x28/m1_710_n388# Vn 3.65f
C308 x28/m1_2498_n384# Vn 0.3f
C309 x28/Vp Vn 12.2f
C310 x28/m1_1594_n962# Vn 0.294f
C311 x16/m1_4146_502# Vn 8.67f
C312 V2 Vn 0.514f
C313 x16/m1_1199_9# Vn 0.378f
C314 x22/Vp Vn 20.5f
C315 x16/Vin Vn 2.78f
C316 V13 Vn 0.861f
C317 x27/m1_546_n454# Vn 1.65f
C318 x27/m1_724_n958# Vn 0.209f
C319 x25/Vin Vn 0.82f
C320 x25/m1_509_303# Vn 0.638f
C321 V11 Vn 0.53f
C322 x31/Vp Vn 7.94f
C323 x25/m1_717_301# Vn 0.249f
C324 x26/m1_532_n361# Vn 0.839f
C325 V12 Vn 1.36f
C326 x26/m1_773_n853# Vn 0.183f
C327 x23/m1_891_n977# Vn 1.15f
C328 V9 Vn 0.49f
C329 x23/m1_1725_85# Vn 0.13f
C330 x22/m1_451_n1105# Vn 0.686f
C331 V8 Vn 0.645f
C332 x22/Vin Vn 4.96f
C333 x21/m1_400_n1066# Vn 0.751f
C334 V7 Vn 0.341f
C335 x21/Vp Vn 12.4f
C336 x31/Vin Vn 1.04f
C337 V1 Vn 0.463f
C338 x31/m1_931_n929# Vn 2.2f
C339 x20/m1_528_n874# Vn 0.727f
C340 V6 Vn 0.76f
C341 x20/Vp Vn 3.33f
C342 x30/Vin Vn 1.37f
C343 Vp Vn 0.36f
C344 th10_0/m1_718_n418# Vn 0.589f
C345 V10 Vn 0.624f
C346 x29/Vp Vn 35.9f
C347 th10_0/m1_878_n414# Vn 0.169f
.ends

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X a_208_47# a_75_199#
+ a_544_297# a_315_47# a_201_297#
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPB a_75_199# 0.0486f
C1 A2 VPB 0.0376f
C2 C1 a_75_199# 0.0628f
C3 A1 VPB 0.0306f
C4 C1 A1 3.21e-19
C5 a_75_199# B1 0.102f
C6 VPB X 0.0107f
C7 VPB A3 0.0268f
C8 A1 B1 0.0716f
C9 VPB VPWR 0.0749f
C10 VPB a_201_297# 0.00186f
C11 C1 X 5.14e-20
C12 C1 VPWR 0.0146f
C13 C1 a_201_297# 0.00243f
C14 a_544_297# B1 1.13e-19
C15 VPB VGND 0.00772f
C16 X B1 7.79e-20
C17 C1 VGND 0.0181f
C18 VPWR B1 0.0125f
C19 a_201_297# B1 0.00594f
C20 A2 a_75_199# 0.0621f
C21 VGND B1 0.0171f
C22 A1 a_75_199# 0.0696f
C23 A1 A2 0.0689f
C24 a_75_199# a_208_47# 0.0159f
C25 A2 a_208_47# 0.00102f
C26 a_544_297# a_75_199# 0.0176f
C27 X a_75_199# 0.0959f
C28 A2 X 3.01e-19
C29 A3 a_75_199# 0.163f
C30 a_75_199# a_315_47# 0.0202f
C31 A2 A3 0.0747f
C32 A2 a_315_47# 0.00335f
C33 VPWR a_75_199# 0.109f
C34 a_75_199# a_201_297# 0.16f
C35 A2 VPWR 0.0174f
C36 A2 a_201_297# 0.0112f
C37 A1 X 1.2e-19
C38 C1 VPB 0.0394f
C39 A1 a_315_47# 0.00313f
C40 A1 VPWR 0.0151f
C41 X a_208_47# 1.91e-19
C42 A1 a_201_297# 0.011f
C43 A3 a_208_47# 3.65e-19
C44 VPWR a_208_47# 8.35e-19
C45 a_544_297# X 2.35e-19
C46 VGND a_75_199# 0.362f
C47 A2 VGND 0.0119f
C48 VPB B1 0.0292f
C49 a_544_297# VPWR 0.0105f
C50 a_544_297# a_201_297# 0.00702f
C51 A3 X 0.00317f
C52 A1 VGND 0.0113f
C53 C1 B1 0.066f
C54 VPWR X 0.0676f
C55 X a_201_297# 0.0131f
C56 VPWR A3 0.0181f
C57 VPWR a_315_47# 0.00154f
C58 A3 a_201_297# 0.00642f
C59 VGND a_208_47# 0.00302f
C60 VPWR a_201_297# 0.211f
C61 a_544_297# VGND 0.00256f
C62 VGND X 0.0609f
C63 VGND A3 0.0161f
C64 VGND a_315_47# 0.00427f
C65 VGND VPWR 0.0735f
C66 VGND a_201_297# 0.00403f
C67 VGND VNB 0.437f
C68 VPWR VNB 0.365f
C69 X VNB 0.0906f
C70 C1 VNB 0.148f
C71 B1 VNB 0.0947f
C72 A1 VNB 0.101f
C73 A2 VNB 0.11f
C74 A3 VNB 0.0908f
C75 VPB VNB 0.782f
C76 a_201_297# VNB 0.00345f
C77 a_75_199# VNB 0.205f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_181_47# a_109_47# a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VGND C 0.0703f
C1 C a_181_47# 0.00151f
C2 X VPB 0.0121f
C3 X B 0.00111f
C4 a_27_47# VGND 0.134f
C5 a_27_47# a_181_47# 0.00401f
C6 a_109_47# VGND 0.00123f
C7 X VPWR 0.0766f
C8 a_27_47# C 0.186f
C9 VGND VPB 0.00604f
C10 A VGND 0.0154f
C11 VGND B 0.00714f
C12 VPB C 0.0347f
C13 B C 0.0746f
C14 VGND VPWR 0.0475f
C15 VPWR a_181_47# 3.97e-19
C16 a_109_47# a_27_47# 0.00517f
C17 VPWR C 0.00464f
C18 a_27_47# VPB 0.0501f
C19 A a_27_47# 0.157f
C20 a_27_47# B 0.0625f
C21 VGND X 0.0708f
C22 a_109_47# A 6.45e-19
C23 X C 0.0149f
C24 a_27_47# VPWR 0.145f
C25 a_109_47# VPWR 3.29e-19
C26 A VPB 0.0426f
C27 B VPB 0.0836f
C28 A B 0.0869f
C29 VGND a_181_47# 0.00261f
C30 VPWR VPB 0.0795f
C31 a_27_47# X 0.087f
C32 A VPWR 0.0185f
C33 VPWR B 0.128f
C34 VGND VNB 0.3f
C35 X VNB 0.0923f
C36 C VNB 0.12f
C37 A VNB 0.174f
C38 VPWR VNB 0.274f
C39 B VNB 0.102f
C40 VPB VNB 0.516f
C41 a_27_47# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
C0 VPWR VPB 0.0625f
C1 VGND VPB 0.0797f
C2 VPWR VGND 0.353f
C3 VPWR VNB 0.47f
C4 VGND VNB 0.427f
C5 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VPWR VPB 0.0787f
C1 VGND VPB 0.116f
C2 VPWR VGND 0.546f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_384_47# a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
C0 a_384_47# a_81_21# 0.00138f
C1 a_81_21# B1 0.148f
C2 VGND A2 0.0495f
C3 VPB a_81_21# 0.0593f
C4 VPWR A2 0.0201f
C5 a_384_47# A1 0.00884f
C6 B1 A1 0.0817f
C7 VPWR VGND 0.0579f
C8 VPB A1 0.0264f
C9 a_81_21# A1 0.0568f
C10 VGND X 0.0512f
C11 VPWR X 0.0847f
C12 a_299_297# A2 0.0468f
C13 a_299_297# VGND 0.00772f
C14 a_299_297# VPWR 0.202f
C15 VPB A2 0.0373f
C16 a_384_47# VGND 0.00366f
C17 a_384_47# VPWR 4.08e-19
C18 VGND B1 0.0181f
C19 VPWR B1 0.0196f
C20 VPB VGND 0.00713f
C21 VPB VPWR 0.068f
C22 A2 a_81_21# 7.47e-19
C23 VGND a_81_21# 0.173f
C24 VPWR a_81_21# 0.146f
C25 A2 A1 0.0921f
C26 X B1 3.04e-20
C27 VPB X 0.0108f
C28 VGND A1 0.0786f
C29 VPWR A1 0.0209f
C30 a_384_47# a_299_297# 1.48e-19
C31 a_299_297# B1 0.00863f
C32 a_81_21# X 0.112f
C33 VPB a_299_297# 0.0111f
C34 a_299_297# a_81_21# 0.0821f
C35 a_299_297# A1 0.0585f
C36 VPB B1 0.0387f
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 VGND A 0.0638f
C1 VGND VPB 0.00649f
C2 VPB A 0.0742f
C3 VPWR VGND 0.0423f
C4 VPWR A 0.0631f
C5 VPWR VPB 0.0521f
C6 Y VGND 0.155f
C7 Y A 0.0894f
C8 Y VPB 0.0061f
C9 VPWR Y 0.209f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X a_29_53# a_183_297# a_111_297#
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 VPWR VGND 0.0459f
C1 VPB B 0.0962f
C2 a_183_297# VGND 5.75e-19
C3 a_111_297# VGND 3.96e-19
C4 VPWR a_183_297# 8.13e-19
C5 A a_29_53# 0.242f
C6 VPWR a_111_297# 5.94e-19
C7 X A 0.00127f
C8 a_29_53# VGND 0.217f
C9 X VGND 0.036f
C10 VPWR a_29_53# 0.0833f
C11 VPWR X 0.0885f
C12 a_183_297# a_29_53# 0.00868f
C13 a_111_297# a_29_53# 0.005f
C14 A C 0.0343f
C15 X a_29_53# 0.0991f
C16 C VGND 0.0161f
C17 VPWR C 0.00457f
C18 VPB A 0.0377f
C19 A B 0.0787f
C20 VPB VGND 0.00724f
C21 a_29_53# C 0.0857f
C22 VPB VPWR 0.0649f
C23 VGND B 0.0152f
C24 VPWR B 0.147f
C25 VPB a_29_53# 0.0491f
C26 VPB X 0.0109f
C27 a_29_53# B 0.121f
C28 X B 6.52e-19
C29 VPB C 0.0396f
C30 C B 0.0802f
C31 A VGND 0.0187f
C32 VPWR A 0.00936f
C33 a_183_297# A 0.00239f
C34 a_111_297# A 0.00223f
C35 VGND VNB 0.306f
C36 X VNB 0.0882f
C37 A VNB 0.117f
C38 C VNB 0.16f
C39 B VNB 0.117f
C40 VPWR VNB 0.253f
C41 VPB VNB 0.516f
C42 a_29_53# VNB 0.18f
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
C0 VPB VGND 0.161f
C1 VPWR VGND 0.903f
C2 VPB VPWR 0.0858f
C3 VPWR VNB 0.867f
C4 VGND VNB 0.761f
C5 VPB VNB 0.605f
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 Y VPB 0.0139f
C1 VPWR B 0.0148f
C2 A B 0.0584f
C3 VGND B 0.0451f
C4 B VPB 0.0367f
C5 Y B 0.0877f
C6 VPWR A 0.0528f
C7 VPWR a_109_297# 0.00638f
C8 VGND VPWR 0.0314f
C9 VPWR VPB 0.0449f
C10 VPWR Y 0.0995f
C11 VGND A 0.0486f
C12 A VPB 0.0415f
C13 VGND a_109_297# 0.00128f
C14 Y A 0.0471f
C15 VGND VPB 0.00456f
C16 Y a_109_297# 0.0113f
C17 VGND Y 0.154f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X a_193_297# a_465_47#
+ a_205_47# a_109_297# a_27_47#
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
C0 A2 VGND 0.0168f
C1 a_109_297# B1 0.00736f
C2 B2 a_193_297# 0.00126f
C3 B2 X 6.77e-20
C4 VPB C1 0.0367f
C5 VPWR B2 0.00842f
C6 A1 VGND 0.0126f
C7 a_193_297# VGND 0.00438f
C8 X VGND 0.061f
C9 VPWR VGND 0.0722f
C10 a_205_47# a_27_47# 0.00762f
C11 A2 a_27_47# 0.153f
C12 B2 VGND 0.0174f
C13 a_27_47# A1 0.0984f
C14 a_27_47# a_193_297# 0.144f
C15 a_27_47# X 0.0921f
C16 B1 C1 6.46e-19
C17 VPWR a_27_47# 0.099f
C18 a_109_297# A1 1.05e-19
C19 a_109_297# a_193_297# 0.0927f
C20 a_109_297# X 3.99e-19
C21 B1 VPB 0.0321f
C22 a_109_297# VPWR 0.15f
C23 a_27_47# B2 0.0959f
C24 a_109_297# B2 0.0133f
C25 a_27_47# VGND 0.395f
C26 A1 a_465_47# 7.06e-19
C27 a_465_47# X 1.56e-19
C28 A2 C1 9.03e-21
C29 a_109_297# VGND 0.00284f
C30 VPWR a_465_47# 5.05e-19
C31 A2 VPB 0.027f
C32 A1 C1 1.77e-20
C33 C1 X 5.03e-20
C34 VPWR C1 0.0139f
C35 A1 VPB 0.0343f
C36 a_465_47# VGND 0.00257f
C37 VPB a_193_297# 0.00774f
C38 VPB X 0.0113f
C39 a_109_297# a_27_47# 0.0961f
C40 VPWR VPB 0.0799f
C41 C1 B2 0.0726f
C42 VPB B2 0.0256f
C43 C1 VGND 0.0196f
C44 a_27_47# a_465_47# 0.013f
C45 VPB VGND 0.00844f
C46 A1 B1 0.0609f
C47 B1 a_193_297# 0.00869f
C48 B1 X 9.58e-20
C49 VPWR B1 0.00982f
C50 a_27_47# C1 0.0792f
C51 B1 B2 0.0784f
C52 a_27_47# VPB 0.0512f
C53 a_109_297# C1 0.00739f
C54 a_109_297# VPB 0.00421f
C55 B1 VGND 0.0133f
C56 A2 A1 0.0692f
C57 A2 a_193_297# 0.00683f
C58 A2 X 0.00157f
C59 a_205_47# VPWR 1.62e-19
C60 A2 VPWR 0.0209f
C61 A1 a_193_297# 0.0109f
C62 A1 X 2.77e-19
C63 a_193_297# X 0.00367f
C64 VPWR A1 0.0161f
C65 a_27_47# B1 0.112f
C66 VPWR a_193_297# 0.169f
C67 VPWR X 0.0897f
C68 a_205_47# VGND 0.00156f
C69 VGND VNB 0.437f
C70 X VNB 0.0919f
C71 VPWR VNB 0.364f
C72 A2 VNB 0.0896f
C73 A1 VNB 0.106f
C74 B1 VNB 0.108f
C75 B2 VNB 0.0887f
C76 C1 VNB 0.139f
C77 VPB VNB 0.782f
C78 a_193_297# VNB 0.0011f
C79 a_109_297# VNB 7.11e-19
C80 a_27_47# VNB 0.216f
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X a_256_47# a_584_47#
+ a_93_21# a_250_297# a_346_47#
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
C0 a_256_47# VGND 0.00394f
C1 a_256_47# a_93_21# 0.0114f
C2 X VGND 0.06f
C3 X a_93_21# 0.0841f
C4 a_584_47# VGND 0.00683f
C5 a_584_47# a_93_21# 0.00278f
C6 VPWR B1 0.01f
C7 VPWR A1 0.016f
C8 X VPB 0.0108f
C9 A1 B1 0.0965f
C10 a_93_21# VGND 0.251f
C11 VGND VPB 0.00788f
C12 a_93_21# VPB 0.0485f
C13 VPWR A2 0.0133f
C14 B1 A2 1.44e-20
C15 B2 VPWR 0.0108f
C16 A1 A2 0.0971f
C17 B2 B1 0.0823f
C18 B2 A1 3.14e-19
C19 VPWR a_250_297# 0.313f
C20 a_250_297# B1 0.0125f
C21 a_250_297# A1 0.0129f
C22 B2 A2 1.46e-19
C23 VPWR A3 0.0158f
C24 a_250_297# A2 0.0129f
C25 B1 A3 7.88e-22
C26 B2 a_250_297# 0.0344f
C27 a_346_47# VPWR 0.00109f
C28 a_346_47# B1 5.39e-20
C29 a_346_47# A1 0.00465f
C30 VPWR a_256_47# 9.47e-19
C31 A2 A3 0.0788f
C32 X VPWR 0.0849f
C33 a_256_47# B1 2.07e-20
C34 VPWR a_584_47# 9.47e-19
C35 B2 A3 9.12e-20
C36 X B1 3.83e-20
C37 X A1 6.03e-20
C38 a_346_47# A2 0.00252f
C39 a_584_47# B1 0.00143f
C40 VPWR VGND 0.076f
C41 VPWR a_93_21# 0.0907f
C42 a_250_297# A3 0.00602f
C43 B1 VGND 0.0344f
C44 A1 VGND 0.0133f
C45 B1 a_93_21# 0.0774f
C46 A1 a_93_21# 0.0641f
C47 a_256_47# A2 0.00256f
C48 X A2 1.19e-19
C49 VPWR VPB 0.0756f
C50 B1 VPB 0.0276f
C51 A1 VPB 0.0296f
C52 A2 VGND 0.0114f
C53 a_93_21# A2 0.0747f
C54 X a_250_297# 5.42e-19
C55 B2 VGND 0.0469f
C56 a_584_47# a_250_297# 2.43e-19
C57 B2 a_93_21# 0.0147f
C58 A2 VPB 0.0287f
C59 a_250_297# VGND 0.0072f
C60 a_250_297# a_93_21# 0.188f
C61 B2 VPB 0.0355f
C62 a_256_47# A3 4.42e-19
C63 X A3 2.45e-19
C64 a_250_297# VPB 0.00616f
C65 A3 VGND 0.00974f
C66 a_93_21# A3 0.124f
C67 a_346_47# VGND 0.00514f
C68 a_346_47# a_93_21# 0.0119f
C69 A3 VPB 0.0291f
C70 VGND VNB 0.465f
C71 VPWR VNB 0.365f
C72 X VNB 0.0937f
C73 B2 VNB 0.14f
C74 B1 VNB 0.101f
C75 A1 VNB 0.0951f
C76 A2 VNB 0.0921f
C77 A3 VNB 0.0929f
C78 VPB VNB 0.782f
C79 a_250_297# VNB 0.0278f
C80 a_93_21# VNB 0.151f
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X a_277_297# a_205_297# a_27_297#
+ a_109_297#
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 C VGND 0.0191f
C1 a_277_297# VGND 4.65e-19
C2 VPB A 0.033f
C3 D a_27_297# 0.054f
C4 C D 0.0954f
C5 B a_27_297# 0.159f
C6 B C 0.0917f
C7 a_277_297# B 2.29e-19
C8 a_27_297# A 0.163f
C9 VGND X 0.0354f
C10 C A 0.028f
C11 a_277_297# A 2.28e-19
C12 VPB a_27_297# 0.0517f
C13 VPB C 0.0338f
C14 a_205_297# a_27_297# 0.00412f
C15 a_109_297# a_27_297# 0.00695f
C16 C a_205_297# 0.00261f
C17 C a_109_297# 0.00356f
C18 B X 6.42e-19
C19 X A 0.00133f
C20 C a_27_297# 0.158f
C21 a_277_297# a_27_297# 0.00876f
C22 VPB X 0.0109f
C23 a_277_297# C 5.54e-19
C24 VGND VPWR 0.0546f
C25 D VPWR 0.00503f
C26 a_27_297# X 0.0991f
C27 B VPWR 0.193f
C28 a_277_297# X 6.43e-20
C29 A VPWR 0.00769f
C30 VPB VPWR 0.075f
C31 a_205_297# VPWR 5.16e-19
C32 a_109_297# VPWR 9.23e-19
C33 a_27_297# VPWR 0.084f
C34 C VPWR 0.00723f
C35 a_277_297# VPWR 7.48e-19
C36 D VGND 0.0517f
C37 B VGND 0.0159f
C38 VGND A 0.016f
C39 VPB VGND 0.00796f
C40 B D 0.00287f
C41 X VPWR 0.0878f
C42 a_205_297# VGND 3.36e-19
C43 a_109_297# VGND 7.58e-19
C44 D A 2.13e-19
C45 B A 0.0639f
C46 VPB D 0.0405f
C47 B VPB 0.106f
C48 VGND a_27_297# 0.235f
C49 VGND VNB 0.367f
C50 X VNB 0.0883f
C51 A VNB 0.109f
C52 C VNB 0.105f
C53 D VNB 0.175f
C54 B VNB 0.115f
C55 VPWR VNB 0.29f
C56 VPB VNB 0.605f
C57 a_27_297# VNB 0.163f
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
C0 VPB VGND 0.35f
C1 VPWR VGND 1.57f
C2 VPB VPWR 0.137f
C3 VPWR VNB 1.67f
C4 VGND VNB 1.47f
C5 VPB VNB 1.14f
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X a_369_47# a_469_47#
+ a_297_47# a_193_413# a_27_47#
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_193_413# a_469_47# 0.00109f
C1 B a_369_47# 0.00129f
C2 a_193_413# X 0.108f
C3 a_193_413# a_27_47# 0.125f
C4 VPWR VPB 0.0818f
C5 C a_369_47# 0.00448f
C6 a_193_413# VGND 0.0915f
C7 VPWR B 0.0186f
C8 a_193_413# a_297_47# 0.00137f
C9 VPWR C 0.0182f
C10 a_193_413# A_N 0.00151f
C11 VPB D 0.0763f
C12 VPWR a_469_47# 7.77e-19
C13 VGND a_369_47# 0.00505f
C14 C D 0.183f
C15 VPWR X 0.0586f
C16 VPWR a_27_47# 0.106f
C17 a_469_47# D 0.00183f
C18 VPWR VGND 0.0727f
C19 VPWR a_297_47# 2.82e-19
C20 VPWR A_N 0.02f
C21 X D 0.0168f
C22 VGND D 0.0372f
C23 B VPB 0.089f
C24 a_193_413# a_369_47# 0.00181f
C25 C VPB 0.0742f
C26 C B 0.164f
C27 VPWR a_193_413# 0.281f
C28 C a_469_47# 0.00202f
C29 VPB X 0.0108f
C30 a_193_413# D 0.155f
C31 VPB a_27_47# 0.092f
C32 B a_27_47# 0.0794f
C33 VPB VGND 0.0123f
C34 B VGND 0.037f
C35 VPWR a_369_47# 6.65e-19
C36 C X 0.00479f
C37 VPB A_N 0.0832f
C38 B a_297_47# 0.00353f
C39 C VGND 0.0395f
C40 a_469_47# X 0.001f
C41 VGND a_469_47# 0.00551f
C42 VPWR D 0.0186f
C43 VGND X 0.0588f
C44 VGND a_27_47# 0.103f
C45 a_193_413# VPB 0.0644f
C46 a_193_413# B 0.144f
C47 a_27_47# A_N 0.237f
C48 VGND a_297_47# 0.00183f
C49 VGND A_N 0.0205f
C50 C a_193_413# 0.0389f
C51 VGND VNB 0.456f
C52 X VNB 0.0934f
C53 VPWR VNB 0.368f
C54 D VNB 0.123f
C55 C VNB 0.108f
C56 B VNB 0.12f
C57 A_N VNB 0.198f
C58 VPB VNB 0.782f
C59 a_193_413# VNB 0.136f
C60 a_27_47# VNB 0.224f
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X a_109_93# a_368_53# a_209_311#
+ a_296_53#
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
C0 a_209_311# C 0.19f
C1 X B 0.00119f
C2 a_109_93# VPWR 0.0984f
C3 VGND a_109_93# 0.0784f
C4 a_209_311# VPWR 0.155f
C5 a_368_53# a_209_311# 0.0026f
C6 C VPB 0.0339f
C7 VGND a_209_311# 0.131f
C8 a_109_93# a_296_53# 1.84e-19
C9 a_209_311# X 0.0877f
C10 a_209_311# a_296_53# 0.0049f
C11 C A_N 7.6e-19
C12 VPB VPWR 0.104f
C13 a_109_93# B 0.0802f
C14 VGND VPB 0.00909f
C15 a_209_311# B 0.0609f
C16 A_N VPWR 0.0513f
C17 X VPB 0.0119f
C18 VGND A_N 0.045f
C19 VPB B 0.0914f
C20 X A_N 1.44e-19
C21 a_209_311# a_109_93# 0.168f
C22 C VPWR 0.005f
C23 a_368_53# C 0.00415f
C24 A_N B 2.03e-19
C25 VGND C 0.0678f
C26 a_109_93# VPB 0.0652f
C27 X C 0.0176f
C28 a_368_53# VPWR 4.26e-19
C29 a_209_311# VPB 0.0515f
C30 VGND VPWR 0.0657f
C31 a_368_53# VGND 0.0031f
C32 C B 0.0671f
C33 a_109_93# A_N 0.117f
C34 X VPWR 0.0732f
C35 VPWR a_296_53# 1.15e-19
C36 a_209_311# A_N 0.00515f
C37 VGND X 0.0647f
C38 VGND a_296_53# 6.07e-19
C39 B VPWR 0.131f
C40 VGND B 0.00796f
C41 a_109_93# C 3.91e-20
C42 A_N VPB 0.111f
C43 VGND VNB 0.44f
C44 X VNB 0.0925f
C45 C VNB 0.114f
C46 B VNB 0.101f
C47 VPWR VNB 0.342f
C48 A_N VNB 0.197f
C49 VPB VNB 0.693f
C50 a_209_311# VNB 0.143f
C51 a_109_93# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
C0 A VGND 0.0431f
C1 VPB a_27_47# 0.139f
C2 a_27_47# X 0.328f
C3 VPWR a_27_47# 0.219f
C4 VPB VGND 0.00583f
C5 X VGND 0.216f
C6 VPWR VGND 0.057f
C7 a_27_47# VGND 0.148f
C8 A VPB 0.0321f
C9 A X 0.014f
C10 A VPWR 0.022f
C11 VPB X 0.0122f
C12 A a_27_47# 0.195f
C13 VPWR VPB 0.0632f
C14 VPWR X 0.317f
C15 VGND VNB 0.358f
C16 X VNB 0.067f
C17 VPWR VNB 0.308f
C18 A VNB 0.148f
C19 VPB VNB 0.605f
C20 a_27_47# VNB 0.543f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
C0 VPB B 0.0629f
C1 a_59_75# A 0.0809f
C2 VPWR a_59_75# 0.15f
C3 A B 0.0971f
C4 X VGND 0.0993f
C5 VPWR B 0.0117f
C6 a_59_75# B 0.143f
C7 X a_145_75# 5.76e-19
C8 VPB X 0.0127f
C9 a_145_75# VGND 0.00468f
C10 X A 1.68e-19
C11 X VPWR 0.111f
C12 X a_59_75# 0.109f
C13 VPB VGND 0.008f
C14 X B 0.00276f
C15 VGND A 0.0147f
C16 VPWR VGND 0.0461f
C17 a_59_75# VGND 0.116f
C18 VPWR a_145_75# 6.31e-19
C19 VGND B 0.0115f
C20 a_145_75# a_59_75# 0.00658f
C21 VPB A 0.0806f
C22 VPB VPWR 0.0729f
C23 VPB a_59_75# 0.0563f
C24 VPWR A 0.0362f
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y a_297_297# a_191_297#
+ a_109_297#
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
C0 D VPWR 0.0128f
C1 VPB C 0.0299f
C2 a_297_297# VPWR 0.00317f
C3 a_191_297# VPWR 0.0049f
C4 a_297_297# B 0.0132f
C5 a_191_297# B 0.00223f
C6 Y A 0.0175f
C7 a_109_297# VPWR 0.00576f
C8 Y VPWR 0.0561f
C9 Y B 0.0403f
C10 D Y 0.108f
C11 Y a_297_297# 1.24e-19
C12 Y a_191_297# 0.00142f
C13 A VGND 0.0526f
C14 VGND VPWR 0.0492f
C15 Y a_109_297# 0.0122f
C16 B VGND 0.0191f
C17 D VGND 0.0456f
C18 a_297_297# VGND 8.1e-19
C19 a_191_297# VGND 9.29e-19
C20 VPB A 0.041f
C21 A C 0.00268f
C22 a_109_297# VGND 0.00181f
C23 VPB VPWR 0.0524f
C24 VPB B 0.0304f
C25 Y VGND 0.151f
C26 VPB D 0.0376f
C27 VPWR C 0.0509f
C28 B C 0.173f
C29 D C 0.0523f
C30 a_191_297# C 0.0195f
C31 VPB Y 0.0127f
C32 a_109_297# C 0.0062f
C33 Y C 0.125f
C34 VPB VGND 0.0048f
C35 VGND C 0.0184f
C36 A VPWR 0.0483f
C37 A B 0.11f
C38 a_297_297# A 3.16e-19
C39 B VPWR 0.0887f
C40 VGND VNB 0.322f
C41 VPWR VNB 0.276f
C42 Y VNB 0.0645f
C43 A VNB 0.174f
C44 B VNB 0.0968f
C45 C VNB 0.0911f
C46 D VNB 0.159f
C47 VPB VNB 0.516f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X a_75_212#
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 VPWR VPB 0.0355f
C1 VGND A 0.0184f
C2 X A 8.48e-19
C3 a_75_212# A 0.178f
C4 A VPB 0.0525f
C5 VPWR A 0.0217f
C6 VGND X 0.0545f
C7 VGND a_75_212# 0.105f
C8 VGND VPB 0.00507f
C9 a_75_212# X 0.107f
C10 VGND VPWR 0.0289f
C11 X VPB 0.0128f
C12 VPWR X 0.0896f
C13 a_75_212# VPB 0.0571f
C14 VPWR a_75_212# 0.134f
C15 VGND VNB 0.207f
C16 VPWR VNB 0.176f
C17 X VNB 0.0942f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_75_212# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 X VPB 0.0128f
C1 VGND A 0.0184f
C2 VPWR A 0.0215f
C3 a_27_47# A 0.181f
C4 A VPB 0.0524f
C5 X A 8.48e-19
C6 VGND VPWR 0.029f
C7 VGND a_27_47# 0.105f
C8 VGND VPB 0.00505f
C9 a_27_47# VPWR 0.135f
C10 VGND X 0.0546f
C11 VPWR VPB 0.0355f
C12 X VPWR 0.0897f
C13 a_27_47# VPB 0.0592f
C14 X a_27_47# 0.107f
C15 VGND VNB 0.207f
C16 X VNB 0.0941f
C17 VPWR VNB 0.175f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_27_47# VNB 0.208f
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X a_664_47# a_841_47#
+ a_381_47# a_62_47# a_558_47#
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPB a_664_47# 0.043f
C1 X a_664_47# 6.67e-19
C2 VPB A 0.105f
C3 X A 0.0142f
C4 VPWR a_664_47# 0.131f
C5 VPWR A 0.0174f
C6 a_841_47# a_664_47# 0.134f
C7 a_381_47# a_558_47# 0.16f
C8 VPB VGND 0.008f
C9 X VGND 0.106f
C10 VPWR VGND 0.0902f
C11 a_62_47# A 0.244f
C12 a_664_47# a_558_47# 0.314f
C13 a_841_47# VGND 0.0585f
C14 a_62_47# VGND 0.144f
C15 VGND a_558_47# 0.0816f
C16 X VPB 0.126f
C17 VPWR VPB 0.103f
C18 a_381_47# A 5.42e-19
C19 VPWR X 0.108f
C20 VPB a_841_47# 0.0108f
C21 VPWR a_841_47# 0.0614f
C22 a_381_47# VGND 0.125f
C23 VPB a_62_47# 0.0515f
C24 X a_62_47# 0.156f
C25 VPWR a_62_47# 0.149f
C26 VPB a_558_47# 0.115f
C27 X a_558_47# 0.0144f
C28 VPWR a_558_47# 0.084f
C29 a_664_47# VGND 0.125f
C30 a_841_47# a_558_47# 0.00368f
C31 A VGND 0.0176f
C32 a_381_47# VPB 0.0447f
C33 a_381_47# X 0.318f
C34 VPWR a_381_47# 0.134f
C35 VGND VNB 0.537f
C36 VPWR VNB 0.439f
C37 X VNB 0.163f
C38 A VNB 0.198f
C39 VPB VNB 0.959f
C40 a_841_47# VNB 0.0929f
C41 a_664_47# VNB 0.13f
C42 a_558_47# VNB 0.164f
C43 a_381_47# VNB 0.11f
C44 a_62_47# VNB 0.169f
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y a_129_47# a_47_47# a_285_47#
+ a_377_297#
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 a_377_297# Y 0.00188f
C1 VGND VPWR 0.0665f
C2 VPWR a_129_47# 9.47e-19
C3 a_285_47# a_47_47# 0.0175f
C4 A Y 0.00181f
C5 Y VPB 0.00878f
C6 a_47_47# VGND 0.104f
C7 a_47_47# a_129_47# 0.00369f
C8 a_377_297# VGND 0.00125f
C9 Y B 0.00334f
C10 a_47_47# VPWR 0.273f
C11 a_285_47# A 0.0353f
C12 a_285_47# VPB 5.53e-19
C13 a_377_297# VPWR 0.00559f
C14 A VGND 0.0635f
C15 VGND VPB 0.00568f
C16 a_285_47# B 0.067f
C17 A VPWR 0.0349f
C18 VPB VPWR 0.0718f
C19 VGND B 0.0389f
C20 B a_129_47# 0.00236f
C21 a_377_297# a_47_47# 0.00899f
C22 a_285_47# Y 0.0439f
C23 B VPWR 0.0408f
C24 A a_47_47# 0.0307f
C25 a_47_47# VPB 0.0444f
C26 VGND Y 0.0381f
C27 Y VPWR 0.107f
C28 a_47_47# B 0.356f
C29 a_285_47# VGND 0.211f
C30 a_377_297# B 0.00254f
C31 A VPB 0.0822f
C32 a_285_47# VPWR 0.00255f
C33 VGND a_129_47# 0.00547f
C34 a_47_47# Y 0.143f
C35 A B 0.236f
C36 B VPB 0.0643f
C37 VGND VNB 0.4f
C38 Y VNB 0.0783f
C39 VPWR VNB 0.352f
C40 A VNB 0.217f
C41 B VNB 0.212f
C42 VPB VNB 0.693f
C43 a_285_47# VNB 0.0174f
C44 a_47_47# VNB 0.199f
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X a_472_297# a_80_21#
+ a_300_47# a_217_297#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
C0 a_472_297# a_80_21# 0.0164f
C1 a_80_21# VPB 0.0661f
C2 VGND a_80_21# 0.293f
C3 X A1 3.62e-19
C4 VPB A2 0.0384f
C5 VGND A2 0.0191f
C6 C1 X 7.15e-20
C7 A1 B1 0.0834f
C8 a_80_21# A2 0.128f
C9 VPWR A1 0.0149f
C10 X B1 1.18e-19
C11 C1 B1 0.0846f
C12 VPWR X 0.0884f
C13 VPWR C1 0.0137f
C14 a_217_297# A1 0.0124f
C15 a_217_297# X 0.00271f
C16 a_217_297# C1 0.00262f
C17 VPWR B1 0.0129f
C18 a_217_297# B1 0.00651f
C19 a_300_47# A1 5.95e-19
C20 VPWR a_217_297# 0.197f
C21 a_300_47# X 5.31e-19
C22 A1 VPB 0.0266f
C23 VGND A1 0.0147f
C24 a_472_297# X 2.6e-19
C25 X VPB 0.0118f
C26 VGND X 0.0654f
C27 C1 VPB 0.0379f
C28 VGND C1 0.0176f
C29 A1 a_80_21# 0.111f
C30 a_300_47# VPWR 8.53e-19
C31 X a_80_21# 0.118f
C32 C1 a_80_21# 0.079f
C33 a_472_297# B1 1.87e-19
C34 A1 A2 0.0881f
C35 B1 VPB 0.0267f
C36 VGND B1 0.0175f
C37 VPWR a_472_297# 0.00703f
C38 VPWR VPB 0.0754f
C39 X A2 6.82e-19
C40 VPWR VGND 0.0665f
C41 a_472_297# a_217_297# 0.00517f
C42 a_217_297# VPB 0.00494f
C43 a_80_21# B1 0.0964f
C44 VGND a_217_297# 0.00342f
C45 VPWR a_80_21# 0.119f
C46 a_217_297# a_80_21# 0.127f
C47 VPWR A2 0.0161f
C48 a_217_297# A2 0.0135f
C49 a_300_47# VGND 0.00536f
C50 VGND a_472_297# 0.00188f
C51 a_300_47# a_80_21# 0.00997f
C52 VGND VPB 0.00775f
C53 VGND VNB 0.385f
C54 VPWR VNB 0.325f
C55 X VNB 0.0899f
C56 C1 VNB 0.144f
C57 B1 VNB 0.0899f
C58 A1 VNB 0.0905f
C59 A2 VNB 0.108f
C60 VPB VNB 0.693f
C61 a_217_297# VNB 0.00117f
C62 a_80_21# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
C0 D VGND 0.0898f
C1 a_303_47# VGND 0.00381f
C2 VPB VPWR 0.077f
C3 a_197_47# VPWR 5.24e-19
C4 a_109_47# VPWR 4.66e-19
C5 C a_27_47# 0.0516f
C6 D C 0.18f
C7 a_303_47# C 0.00527f
C8 a_27_47# VPWR 0.326f
C9 VGND X 0.0903f
C10 D VPWR 0.0207f
C11 a_303_47# VPWR 4.83e-19
C12 VPB a_27_47# 0.082f
C13 VGND B 0.0453f
C14 VPB D 0.0782f
C15 a_197_47# a_27_47# 0.00167f
C16 a_109_47# a_27_47# 0.00578f
C17 C B 0.161f
C18 X VPWR 0.0945f
C19 D a_27_47# 0.107f
C20 a_303_47# a_27_47# 0.00119f
C21 B VPWR 0.0231f
C22 a_303_47# D 0.00119f
C23 VPB X 0.0111f
C24 VPB B 0.0643f
C25 VGND A 0.0151f
C26 a_197_47# B 0.00623f
C27 a_109_47# B 0.00153f
C28 a_27_47# X 0.0754f
C29 D X 0.00746f
C30 a_27_47# B 0.13f
C31 VPWR A 0.044f
C32 VPB A 0.0907f
C33 a_27_47# A 0.153f
C34 C VGND 0.0408f
C35 VGND VPWR 0.0662f
C36 VPB VGND 0.00852f
C37 a_197_47# VGND 0.00387f
C38 a_109_47# VGND 0.00223f
C39 B A 0.0839f
C40 C VPWR 0.021f
C41 VPB C 0.0609f
C42 a_197_47# C 0.00123f
C43 a_109_47# C 1.72e-20
C44 VGND a_27_47# 0.132f
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X a_489_413# a_226_47#
+ a_556_47# a_226_297# a_76_199#
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_226_47# A2_N 0.141f
C1 a_226_47# a_76_199# 0.188f
C2 A1_N VPB 0.0339f
C3 B2 a_226_47# 0.0975f
C4 a_226_47# VGND 0.149f
C5 a_226_47# a_489_413# 0.00579f
C6 A1_N X 0.00211f
C7 VPB VPWR 0.0951f
C8 B1 VPWR 0.0188f
C9 a_76_199# a_226_297# 0.00354f
C10 VGND a_226_297# 5.63e-19
C11 X VPWR 0.0589f
C12 A1_N A2_N 0.11f
C13 A1_N a_76_199# 0.119f
C14 a_556_47# VPWR 7.24e-19
C15 A1_N VGND 0.0261f
C16 A2_N VPWR 0.00449f
C17 a_76_199# VPWR 0.2f
C18 B2 VPWR 0.0161f
C19 VGND VPWR 0.0743f
C20 VPWR a_489_413# 0.143f
C21 B1 VPB 0.0803f
C22 a_226_47# a_226_297# 0.00128f
C23 X VPB 0.0113f
C24 A1_N a_226_47# 0.0209f
C25 VPB A2_N 0.0327f
C26 a_226_47# VPWR 0.0187f
C27 VPB a_76_199# 0.0817f
C28 B1 a_76_199# 0.00185f
C29 B2 VPB 0.0645f
C30 VPB VGND 0.0128f
C31 B2 B1 0.182f
C32 B1 VGND 0.0471f
C33 A1_N a_226_297# 0.00184f
C34 X A2_N 2.55e-19
C35 X a_76_199# 0.0995f
C36 VPB a_489_413# 0.015f
C37 B1 a_489_413# 0.0382f
C38 X VGND 0.0627f
C39 a_76_199# a_556_47# 0.0017f
C40 B2 a_556_47# 0.00291f
C41 VGND a_556_47# 0.00639f
C42 a_226_297# VPWR 8.54e-19
C43 a_76_199# A2_N 0.0125f
C44 A1_N VPWR 0.00672f
C45 VGND A2_N 0.0174f
C46 B2 a_76_199# 0.0626f
C47 VGND a_76_199# 0.108f
C48 B2 VGND 0.0335f
C49 a_226_47# VPB 0.111f
C50 a_76_199# a_489_413# 0.0473f
C51 B2 a_489_413# 0.0541f
C52 VGND a_489_413# 0.0058f
C53 X a_226_47# 0.0108f
C54 VGND VNB 0.462f
C55 A2_N VNB 0.103f
C56 A1_N VNB 0.111f
C57 VPWR VNB 0.369f
C58 X VNB 0.0975f
C59 B1 VNB 0.206f
C60 B2 VNB 0.106f
C61 VPB VNB 0.782f
C62 a_489_413# VNB 0.0254f
C63 a_226_47# VNB 0.162f
C64 a_76_199# VNB 0.141f
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X a_515_93# a_223_47#
+ a_615_93# a_343_93# a_429_93# a_27_47#
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
C0 D VGND 0.0414f
C1 a_223_47# B_N 0.0431f
C2 VPWR A_N 0.0318f
C3 C VGND 0.025f
C4 a_343_93# VGND 0.0548f
C5 X VGND 0.0609f
C6 VPWR VGND 0.0906f
C7 a_429_93# a_223_47# 0.00492f
C8 A_N VGND 0.0146f
C9 D a_223_47# 4.03e-19
C10 a_27_47# a_343_93# 0.0406f
C11 B_N VPB 0.0646f
C12 VPWR a_27_47# 0.0897f
C13 a_223_47# C 0.151f
C14 a_223_47# a_343_93# 0.269f
C15 a_223_47# VPWR 0.114f
C16 a_27_47# A_N 0.0906f
C17 D a_615_93# 0.00564f
C18 a_223_47# A_N 0.00833f
C19 a_27_47# VGND 0.0715f
C20 C a_515_93# 0.00389f
C21 a_515_93# a_343_93# 0.00115f
C22 D VPB 0.081f
C23 a_223_47# VGND 0.199f
C24 VPWR a_515_93# 7.86e-19
C25 C a_615_93# 0.00407f
C26 a_615_93# a_343_93# 0.00103f
C27 VPWR a_615_93# 8.49e-19
C28 C VPB 0.0686f
C29 VPB a_343_93# 0.0857f
C30 VPB X 0.0103f
C31 VPWR VPB 0.106f
C32 a_515_93# VGND 0.00408f
C33 a_223_47# a_27_47# 0.267f
C34 a_615_93# VGND 0.0044f
C35 VPB A_N 0.0848f
C36 VPB VGND 0.0167f
C37 D B_N 6.67e-20
C38 C B_N 9.56e-20
C39 a_223_47# a_515_93# 0.00482f
C40 B_N a_343_93# 0.00112f
C41 B_N X 4.64e-20
C42 VPWR B_N 0.0168f
C43 a_27_47# VPB 0.154f
C44 B_N A_N 0.117f
C45 a_223_47# VPB 0.0799f
C46 B_N VGND 0.0427f
C47 a_429_93# a_343_93# 0.00484f
C48 D C 0.163f
C49 D a_343_93# 0.114f
C50 D X 0.0193f
C51 a_429_93# VPWR 5.19e-19
C52 D VPWR 0.0143f
C53 C a_343_93# 0.0397f
C54 a_343_93# X 0.126f
C55 VPWR C 0.012f
C56 a_27_47# B_N 0.138f
C57 VPWR a_343_93# 0.255f
C58 VPWR X 0.0582f
C59 a_429_93# VGND 0.00122f
C60 VGND VNB 0.553f
C61 X VNB 0.0908f
C62 VPWR VNB 0.453f
C63 D VNB 0.124f
C64 C VNB 0.107f
C65 B_N VNB 0.134f
C66 A_N VNB 0.144f
C67 VPB VNB 0.959f
C68 a_343_93# VNB 0.172f
C69 a_223_47# VNB 0.141f
C70 a_27_47# VNB 0.259f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 a_285_47# B 3.98e-19
C1 a_285_297# a_35_297# 0.025f
C2 a_35_297# VPB 0.0699f
C3 a_285_297# B 0.0553f
C4 VPB B 0.0697f
C5 X VGND 0.173f
C6 a_35_297# B 0.203f
C7 VGND VPWR 0.0643f
C8 X VPWR 0.0537f
C9 a_117_297# VGND 0.00177f
C10 a_117_297# X 2.25e-19
C11 a_117_297# VPWR 0.00852f
C12 VGND A 0.0325f
C13 X A 0.00166f
C14 a_285_47# VGND 0.00552f
C15 a_285_47# X 0.00206f
C16 VPWR A 0.0348f
C17 a_285_297# VGND 0.00394f
C18 a_285_297# X 0.0712f
C19 VGND VPB 0.00696f
C20 X VPB 0.0154f
C21 a_285_47# VPWR 8.6e-19
C22 VGND a_35_297# 0.177f
C23 X a_35_297# 0.166f
C24 a_285_297# VPWR 0.246f
C25 VPWR VPB 0.0689f
C26 VGND B 0.0304f
C27 X B 0.0149f
C28 a_35_297# VPWR 0.096f
C29 VPWR B 0.0703f
C30 a_117_297# a_35_297# 0.00641f
C31 a_285_297# A 0.00749f
C32 A VPB 0.051f
C33 a_117_297# B 0.00777f
C34 a_35_297# A 0.0633f
C35 a_285_297# VPB 0.0133f
C36 a_285_47# a_35_297# 0.00723f
C37 A B 0.221f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X a_465_297# a_297_297#
+ a_215_297# a_392_297# a_109_53#
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 VGND C 0.0202f
C1 a_297_297# C 0.00375f
C2 a_109_53# C 0.0984f
C3 B a_215_297# 0.159f
C4 a_297_297# VGND 6.5e-19
C5 a_109_53# VGND 0.118f
C6 VPWR a_215_297# 0.0871f
C7 a_109_53# a_297_297# 7.06e-21
C8 VPWR D_N 0.0412f
C9 a_392_297# VPWR 5.29e-19
C10 a_215_297# C 0.161f
C11 X A 0.00127f
C12 a_392_297# C 0.00267f
C13 VGND a_215_297# 0.237f
C14 a_297_297# a_215_297# 0.00659f
C15 a_109_53# a_215_297# 0.0807f
C16 D_N VGND 0.0531f
C17 a_392_297# VGND 3.44e-19
C18 D_N a_109_53# 0.0889f
C19 B A 0.0666f
C20 VPWR A 0.0073f
C21 A C 0.0281f
C22 D_N a_215_297# 3.19e-19
C23 a_392_297# a_215_297# 0.00419f
C24 VGND A 0.0158f
C25 a_109_53# A 1.19e-19
C26 X VPB 0.011f
C27 VPWR a_465_297# 7.08e-19
C28 B VPB 0.116f
C29 a_215_297# A 0.157f
C30 a_465_297# C 6.89e-19
C31 VPWR VPB 0.122f
C32 a_465_297# VGND 5.02e-19
C33 C VPB 0.0337f
C34 VGND VPB 0.0115f
C35 a_109_53# VPB 0.0547f
C36 a_465_297# a_215_297# 0.00827f
C37 a_215_297# VPB 0.0508f
C38 D_N VPB 0.0461f
C39 B X 6.65e-19
C40 VPWR X 0.0885f
C41 a_465_297# A 5.42e-19
C42 VPWR B 0.255f
C43 A VPB 0.0325f
C44 VGND X 0.0359f
C45 B C 0.0893f
C46 VPWR C 0.00753f
C47 VGND B 0.0161f
C48 a_109_53# B 0.0246f
C49 VPWR VGND 0.075f
C50 X a_215_297# 0.0991f
C51 VPWR a_297_297# 8.59e-19
C52 VPWR a_109_53# 0.0418f
C53 VGND VNB 0.469f
C54 X VNB 0.0884f
C55 A VNB 0.108f
C56 C VNB 0.101f
C57 D_N VNB 0.185f
C58 B VNB 0.101f
C59 VPWR VNB 0.399f
C60 VPB VNB 0.782f
C61 a_109_53# VNB 0.159f
C62 a_215_297# VNB 0.142f
.ends

.subckt therm b[0] b[2] p[11] p[12] p[13] p[14] p[2] p[5] p[8] input3/a_27_47# _35_/a_226_47#
+ input4/a_75_212# _50_/a_27_47# _45_/a_465_47# net7 input13/a_27_47# _45_/a_205_47#
+ _30_/a_215_297# output19/a_27_47# net19 _45_/a_27_47# input10/a_27_47# _18_ _10_
+ _31_/a_285_47# _31_/a_35_297# _50_/a_429_93# _07_ input7/a_27_47# _04_ output16/a_27_47#
+ input9/a_75_212# _30_/a_109_53# _39_/a_129_47# b[1] _27_/a_27_297# input1/a_75_212#
+ _41_/a_59_75# input5/a_62_47# net3 input14/a_27_47# b[3] _31_/a_285_297# _11_ net2
+ _47_/a_81_21# _49_/a_208_47# p[0] _09_ net14 _13_ _34_/a_47_47# _19_ input11/a_27_47#
+ net12 _34_/a_285_47# _49_/a_75_199# net4 _47_/a_384_47# net8 net6 _17_ input8/a_27_47#
+ _33_/a_209_311# _41_/a_145_75# output17/a_27_47# p[7] _01_ _37_/a_27_47# _38_/a_109_47#
+ _47_/a_299_297# _44_/a_93_21# _44_/a_250_297# p[9] net13 _02_ input15/a_27_47# _39_/a_47_47#
+ _43_/a_27_47# p[1] _50_/a_223_47# _50_/a_515_93# input2/a_27_47# _38_/a_197_47#
+ _15_ _50_/a_615_93# _14_ input12/a_27_47# p[3] _20_ net1 _38_/a_27_47# VPWR _34_/a_129_47#
+ net11 _03_ _06_ _49_/a_315_47# net16 net10 output18/a_27_47# _08_ _16_ _34_/a_377_297#
+ _12_ net9 _00_ _05_ p[4] input6/a_27_47# _39_/a_285_47# net17 _31_/a_117_297# m1_7039_1799#
+ _50_/a_343_93# net5 p[10] _39_/a_377_297# net15 VGND p[6]
X_49_ net7 _02_ _19_ _20_ _21_ VGND VGND VPWR VPWR net17 _49_/a_208_47# _49_/a_75_199#
+ _49_/a_544_297# _49_/a_315_47# _49_/a_201_297# sky130_fd_sc_hd__a311o_1
X_48_ net11 _02_ _07_ VGND VGND VPWR VPWR _21_ _48_/a_181_47# _48_/a_109_47# _48_/a_27_47#
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ net5 _12_ _17_ VGND VGND VPWR VPWR _20_ _47_/a_384_47# _47_/a_81_21# _47_/a_299_297#
+ sky130_fd_sc_hd__a21o_1
X_46_ _04_ VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__inv_2
X_29_ net11 net13 net12 VGND VGND VPWR VPWR _03_ _29_/a_29_53# _29_/a_183_297# _29_/a_111_297#
+ sky130_fd_sc_hd__or3_1
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28_ _00_ _01_ VGND VGND VPWR VPWR _02_ _28_/a_109_297# sky130_fd_sc_hd__nor2_1
X_45_ _02_ _09_ _12_ _13_ _18_ VGND VGND VPWR VPWR net16 _45_/a_193_297# _45_/a_465_47#
+ _45_/a_205_47# _45_/a_109_297# _45_/a_27_47# sky130_fd_sc_hd__a221o_1
X_44_ net14 _14_ _15_ _17_ net2 VGND VGND VPWR VPWR _18_ _44_/a_256_47# _44_/a_584_47#
+ _44_/a_93_21# _44_/a_250_297# _44_/a_346_47# sky130_fd_sc_hd__a32o_1
X_27_ net14 net15 net3 net2 VGND VGND VPWR VPWR _01_ _27_/a_277_297# _27_/a_205_297#
+ _27_/a_27_297# _27_/a_109_297# sky130_fd_sc_hd__or4_1
XFILLER_0_7_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_26_ net5 net4 net6 VGND VGND VPWR VPWR _00_ _26_/a_29_53# _26_/a_183_297# _26_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_43_ _00_ _06_ _10_ _16_ VGND VGND VPWR VPWR _17_ _43_/a_369_47# _43_/a_469_47# _43_/a_297_47#
+ _43_/a_193_413# _43_/a_27_47# sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_42_ net3 net15 net14 VGND VGND VPWR VPWR _16_ _42_/a_109_93# _42_/a_368_53# _42_/a_209_311#
+ _42_/a_296_53# sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_3_Left_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND VPWR VPWR b[0] output16/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_41_ _06_ _10_ VGND VGND VPWR VPWR _15_ _41_/a_145_75# _41_/a_59_75# sky130_fd_sc_hd__and2_1
Xoutput17 net17 VGND VGND VPWR VPWR b[1] output17/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_40_ net15 net3 net2 _00_ VGND VGND VPWR VPWR _14_ _40_/a_297_297# _40_/a_191_297#
+ _40_/a_109_297# sky130_fd_sc_hd__nor4_1
Xoutput18 net18 VGND VGND VPWR VPWR b[2] output18/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR b[3] output19/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_7_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 p[0] VGND VGND VPWR VPWR net1 input1/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput2 p[10] VGND VGND VPWR VPWR net2 input2/a_27_47# sky130_fd_sc_hd__buf_1
Xinput3 p[11] VGND VGND VPWR VPWR net3 input3/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 p[12] VGND VGND VPWR VPWR net4 input4/a_75_212# sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 p[13] VGND VGND VPWR VPWR net5 input5/a_664_47# input5/a_841_47# input5/a_381_47#
+ input5/a_62_47# input5/a_558_47# sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_1_Left_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 p[14] VGND VGND VPWR VPWR net6 input6/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 p[1] VGND VGND VPWR VPWR net7 input7/a_27_47# sky130_fd_sc_hd__buf_1
Xinput10 p[4] VGND VGND VPWR VPWR net10 input10/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 p[2] VGND VGND VPWR VPWR net8 input8/a_27_47# sky130_fd_sc_hd__buf_1
Xinput11 p[5] VGND VGND VPWR VPWR net11 input11/a_27_47# sky130_fd_sc_hd__buf_1
X_39_ net5 net6 VGND VGND VPWR VPWR _13_ _39_/a_129_47# _39_/a_47_47# _39_/a_285_47#
+ _39_/a_377_297# sky130_fd_sc_hd__xnor2_1
Xinput9 p[3] VGND VGND VPWR VPWR net9 input9/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput12 p[6] VGND VGND VPWR VPWR net12 input12/a_27_47# sky130_fd_sc_hd__buf_1
X_55_ _14_ _15_ _20_ _22_ VGND VGND VPWR VPWR net19 _55_/a_472_297# _55_/a_80_21#
+ _55_/a_300_47# _55_/a_217_297# sky130_fd_sc_hd__a211o_1
X_38_ net4 _06_ _10_ _11_ VGND VGND VPWR VPWR _12_ _38_/a_109_47# _38_/a_197_47# _38_/a_303_47#
+ _38_/a_27_47# sky130_fd_sc_hd__and4_1
X_54_ _25_ VGND VGND VPWR VPWR net18 _54_/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput13 p[7] VGND VGND VPWR VPWR net13 input13/a_27_47# sky130_fd_sc_hd__buf_1
X_37_ net14 net15 net3 net2 VGND VGND VPWR VPWR _11_ _37_/a_109_47# _37_/a_197_47#
+ _37_/a_303_47# _37_/a_27_47# sky130_fd_sc_hd__and4_1
X_53_ _21_ _22_ _24_ VGND VGND VPWR VPWR _25_ _53_/a_29_53# _53_/a_183_297# _53_/a_111_297#
+ sky130_fd_sc_hd__or3_1
Xinput14 p[8] VGND VGND VPWR VPWR net14 input14/a_27_47# sky130_fd_sc_hd__buf_1
X_36_ net11 net10 net13 net12 VGND VGND VPWR VPWR _10_ _36_/a_109_47# _36_/a_197_47#
+ _36_/a_303_47# _36_/a_27_47# sky130_fd_sc_hd__and4_1
X_52_ _02_ _06_ _23_ _12_ net5 VGND VGND VPWR VPWR _24_ _52_/a_256_47# _52_/a_584_47#
+ _52_/a_93_21# _52_/a_250_297# _52_/a_346_47# sky130_fd_sc_hd__a32o_1
X_35_ _04_ _05_ _07_ _08_ VGND VGND VPWR VPWR _09_ _35_/a_489_413# _35_/a_226_47#
+ _35_/a_556_47# _35_/a_226_297# _35_/a_76_199# sky130_fd_sc_hd__a2bb2o_1
Xinput15 p[9] VGND VGND VPWR VPWR net15 input15/a_27_47# sky130_fd_sc_hd__buf_1
X_51_ _03_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__inv_2
X_34_ net11 net12 VGND VGND VPWR VPWR _08_ _34_/a_129_47# _34_/a_47_47# _34_/a_285_47#
+ _34_/a_377_297# sky130_fd_sc_hd__xnor2_1
X_33_ net13 _06_ net10 VGND VGND VPWR VPWR _07_ _33_/a_109_93# _33_/a_368_53# _33_/a_209_311#
+ _33_/a_296_53# sky130_fd_sc_hd__and3b_1
X_50_ net5 net6 _15_ _11_ VGND VGND VPWR VPWR _22_ _50_/a_515_93# _50_/a_223_47# _50_/a_615_93#
+ _50_/a_343_93# _50_/a_429_93# _50_/a_27_47# sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ net7 net1 net9 net8 VGND VGND VPWR VPWR _06_ _32_/a_109_47# _32_/a_197_47# _32_/a_303_47#
+ _32_/a_27_47# sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_5_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31_ net7 net8 VGND VGND VPWR VPWR _05_ _31_/a_117_297# _31_/a_285_297# _31_/a_285_47#
+ _31_/a_35_297# sky130_fd_sc_hd__xor2_1
X_30_ net9 net10 _03_ net1 VGND VGND VPWR VPWR _04_ _30_/a_465_297# _30_/a_297_297#
+ _30_/a_215_297# _30_/a_392_297# _30_/a_109_53# sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
C0 net2 net3 0.518f
C1 b[1] input3/a_27_47# 1.31e-20
C2 _16_ input15/a_27_47# 7.13e-19
C3 _10_ _55_/a_472_297# 7.35e-21
C4 _24_ _22_ 0.0846f
C5 _06_ _45_/a_193_297# 0.00201f
C6 VGND _40_/a_191_297# -9.29e-19
C7 _30_/a_109_53# _22_ 3.67e-21
C8 _42_/a_209_311# net3 0.029f
C9 _35_/a_76_199# _33_/a_109_93# 3.08e-19
C10 net10 _13_ 4.52e-21
C11 _45_/a_27_47# _18_ 0.00347f
C12 _19_ _27_/a_109_297# 7.54e-21
C13 _17_ _20_ 0.102f
C14 VGND net12 0.345f
C15 VGND _05_ 0.754f
C16 _50_/a_615_93# net6 1.43e-19
C17 _28_/a_109_297# b[3] 7.49e-20
C18 _01_ net1 0.0509f
C19 _34_/a_47_47# _04_ 1.17e-20
C20 _39_/a_47_47# p[12] 0.00185f
C21 net19 p[12] 6.8e-20
C22 VPWR p[11] 0.194f
C23 net10 _09_ 0.037f
C24 net7 input5/a_558_47# 0.00358f
C25 net18 _21_ 0.00215f
C26 net9 _29_/a_183_297# 3.51e-19
C27 p[4] p[5] 0.332f
C28 net5 _14_ 3.89e-19
C29 _36_/a_27_47# net1 6.99e-20
C30 p[2] input7/a_27_47# 0.0023f
C31 net13 _49_/a_75_199# 3.2e-19
C32 net1 _22_ 0.0129f
C33 _19_ p[10] 0.00289f
C34 _15_ net7 8.4e-20
C35 _52_/a_93_21# net18 8.21e-21
C36 _01_ _21_ 7.94e-19
C37 _40_/a_109_297# net15 0.0016f
C38 _01_ net8 0.0802f
C39 _11_ b[3] 2.37e-20
C40 net11 _13_ 2.34e-19
C41 _36_/a_27_47# _21_ 0.0276f
C42 _06_ _40_/a_191_297# 5.84e-19
C43 VGND _44_/a_250_297# -0.00591f
C44 _22_ _21_ 0.00314f
C45 _36_/a_27_47# net8 1.52e-19
C46 _31_/a_35_297# _49_/a_75_199# 6.24e-19
C47 VPWR _35_/a_489_413# -0.00725f
C48 net8 _22_ 3.3e-20
C49 _23_ net6 2.13e-19
C50 _36_/a_197_47# net13 1.06e-19
C51 net1 input5/a_62_47# 7.59e-20
C52 _07_ _35_/a_556_47# 0.00128f
C53 _34_/a_129_47# _08_ 3.29e-19
C54 _06_ net12 0.284f
C55 net11 _09_ 0.0262f
C56 _04_ input5/a_664_47# 6.73e-21
C57 net16 _25_ 1.16e-19
C58 _52_/a_93_21# _22_ 0.0347f
C59 _06_ _05_ 0.00724f
C60 p[8] input6/a_27_47# 0.00805f
C61 b[2] _09_ 4.28e-20
C62 net9 _32_/a_27_47# 0.0136f
C63 _11_ net4 0.0858f
C64 _31_/a_285_297# _01_ 1.92e-19
C65 input13/a_27_47# _09_ 1.27e-21
C66 output19/a_27_47# p[12] 1.78e-19
C67 _19_ _49_/a_208_47# 7.12e-20
C68 _45_/a_27_47# net6 0.021f
C69 p[8] _37_/a_303_47# 6.41e-20
C70 net2 net19 0.599f
C71 net8 input5/a_62_47# 2.05e-19
C72 _48_/a_27_47# net12 0.0126f
C73 _11_ _45_/a_193_297# 0.0292f
C74 _18_ net7 2.58e-20
C75 _10_ _47_/a_81_21# 0.0061f
C76 VPWR net17 0.0371f
C77 _37_/a_197_47# net14 6.99e-19
C78 _33_/a_109_93# _09_ 7.36e-20
C79 _49_/a_544_297# _09_ 2.56e-20
C80 _23_ _03_ 0.0564f
C81 _42_/a_209_311# net19 0.0766f
C82 _17_ _00_ 0.0851f
C83 _07_ b[1] 1.59e-19
C84 _14_ _44_/a_93_21# 0.04f
C85 _10_ _39_/a_285_47# 0.00289f
C86 VPWR net15 0.61f
C87 _35_/a_226_47# _22_ 1.39e-20
C88 net2 input5/a_381_47# 0.0138f
C89 _29_/a_29_53# net10 1.77e-19
C90 p[8] b[3] 0.237f
C91 net9 _20_ 0.328f
C92 VGND net18 0.255f
C93 _04_ input9/a_75_212# 7.69e-22
C94 _45_/a_27_47# _03_ 2.06e-20
C95 _32_/a_109_47# _02_ 3.98e-19
C96 p[3] _09_ 1.47e-21
C97 _42_/a_209_311# input5/a_381_47# 3.88e-19
C98 _42_/a_109_93# input5/a_558_47# 1.75e-19
C99 p[4] p[6] 0.382f
C100 VPWR net10 0.375f
C101 _10_ net14 2.4e-19
C102 VGND _52_/a_584_47# -0.00112f
C103 VGND _01_ 0.0939f
C104 _01_ _43_/a_193_413# 8.16e-19
C105 _07_ _03_ 0.0113f
C106 _25_ output18/a_27_47# 0.072f
C107 output17/a_27_47# b[3] 0.00196f
C108 _42_/a_109_93# _15_ 0.00367f
C109 input15/a_27_47# _14_ 9.48e-21
C110 net2 output19/a_27_47# 0.00168f
C111 _23_ _08_ 1.81e-19
C112 _17_ _04_ 4.34e-19
C113 VGND _36_/a_27_47# 0.0211f
C114 _11_ _40_/a_191_297# 0.00207f
C115 VGND _22_ 0.0404f
C116 _40_/a_109_297# net3 3.14e-19
C117 _17_ _50_/a_223_47# 5.24e-20
C118 _14_ _43_/a_369_47# 0.00135f
C119 _22_ _43_/a_193_413# 0.00133f
C120 _23_ _02_ 0.0648f
C121 _00_ _26_/a_111_297# 3.7e-19
C122 net13 _18_ 1.06e-20
C123 _29_/a_29_53# net11 0.00514f
C124 VPWR _40_/a_297_297# -5.42e-19
C125 _11_ net12 3.82e-21
C126 b[0] net6 2.52e-19
C127 b[0] b[1] 0.156f
C128 p[13] b[3] 0.128f
C129 VPWR input2/a_27_47# 0.00872f
C130 b[1] net7 0.00382f
C131 VPWR net11 0.996f
C132 net5 _47_/a_81_21# 4.59e-19
C133 _49_/a_315_47# _09_ 1.11e-20
C134 _30_/a_109_53# net17 4.18e-20
C135 _06_ net18 0.0211f
C136 VPWR b[2] 0.26f
C137 VGND input5/a_62_47# 0.0489f
C138 input1/a_75_212# p[0] 0.0172f
C139 _10_ net5 0.199f
C140 input7/a_27_47# input5/a_664_47# 1.08e-21
C141 _16_ b[3] 3.71e-19
C142 _45_/a_27_47# _02_ 0.00449f
C143 _07_ _08_ 0.348f
C144 VPWR input13/a_27_47# 0.0696f
C145 b[1] _38_/a_109_47# 5.74e-20
C146 _39_/a_47_47# _13_ 0.00117f
C147 net5 _39_/a_285_47# 0.05f
C148 _06_ _52_/a_584_47# 0.00218f
C149 _41_/a_59_75# _20_ 1.78e-20
C150 _01_ _06_ 0.00157f
C151 _35_/a_489_413# _21_ 0.0448f
C152 VGND _45_/a_205_47# -2.47e-19
C153 _27_/a_27_297# b[3] 4.34e-19
C154 _07_ _02_ 0.0083f
C155 _29_/a_29_53# net3 1.68e-20
C156 _36_/a_27_47# _06_ 0.0501f
C157 _06_ _22_ 0.124f
C158 _30_/a_215_297# _20_ 6.08e-19
C159 _39_/a_47_47# _09_ 7.7e-21
C160 VPWR _33_/a_109_93# -0.00817f
C161 VPWR _49_/a_544_297# 0.00569f
C162 _16_ net4 2.73e-20
C163 net1 net17 2.89e-19
C164 net9 _00_ 0.00501f
C165 _03_ net7 0.078f
C166 VPWR net3 0.341f
C167 _30_/a_109_53# net10 5.6e-20
C168 _50_/a_27_47# _00_ 0.00197f
C169 p[5] b[3] 0.295f
C170 net5 net14 0.0263f
C171 p[8] _40_/a_191_297# 2.5e-19
C172 net1 net15 7.44e-20
C173 _29_/a_29_53# p[3] 2.07e-19
C174 net13 _26_/a_29_53# 2.23e-20
C175 _50_/a_27_47# _38_/a_27_47# 2.37e-20
C176 _27_/a_277_297# net15 1.93e-19
C177 net17 net8 0.18f
C178 net13 net6 0.00188f
C179 _55_/a_300_47# _14_ 8.09e-19
C180 VPWR p[3] 0.0933f
C181 _52_/a_250_297# net4 0.00136f
C182 net13 b[1] 1.69e-19
C183 _42_/a_368_53# b[3] 4.8e-20
C184 net8 net15 0.2f
C185 net10 net1 0.00388f
C186 input11/a_27_47# b[1] 0.00155f
C187 _19_ _20_ 0.00734f
C188 _12_ _38_/a_197_47# 0.00173f
C189 _10_ _44_/a_93_21# 2.48e-19
C190 _24_ b[2] 1.85e-19
C191 net9 _04_ 0.0213f
C192 _08_ net7 9.54e-25
C193 VGND p[11] 0.148f
C194 _30_/a_109_53# input2/a_27_47# 1.54e-20
C195 _30_/a_297_297# net12 7.14e-21
C196 _20_ _55_/a_217_297# 0.0013f
C197 _50_/a_27_47# _04_ 2.07e-21
C198 _50_/a_223_47# net9 2e-19
C199 output17/a_27_47# _05_ 1.12e-19
C200 _31_/a_35_297# b[1] 1.56e-19
C201 net16 net4 0.155f
C202 _12_ p[12] 0.00639f
C203 net10 _21_ 0.0275f
C204 _02_ net7 0.445f
C205 p[2] net7 0.00156f
C206 _04_ _27_/a_109_297# 7.2e-20
C207 _44_/a_250_297# p[8] 6.66e-20
C208 net10 net8 2.05e-21
C209 net13 _03_ 0.271f
C210 _38_/a_109_47# _02_ 1.63e-19
C211 net16 _45_/a_193_297# 0.00187f
C212 _52_/a_93_21# net10 7.84e-20
C213 _41_/a_59_75# _00_ 2.43e-20
C214 VPWR _49_/a_315_47# 6.26e-19
C215 input6/a_27_47# _14_ 3.75e-21
C216 _43_/a_27_47# net7 6.31e-19
C217 net1 input2/a_27_47# 4.81e-19
C218 VGND _35_/a_489_413# -8.78e-19
C219 net14 _44_/a_93_21# 0.0646f
C220 net11 net1 1.13e-19
C221 _12_ _45_/a_109_297# 0.00587f
C222 _10_ input15/a_27_47# 4.5e-19
C223 _04_ p[10] 0.00265f
C224 p[7] _09_ 9.25e-21
C225 _11_ _22_ 0.15f
C226 input13/a_27_47# net1 1.9e-19
C227 _10_ _43_/a_369_47# 0.00199f
C228 _37_/a_27_47# net2 0.0692f
C229 input5/a_841_47# _02_ 0.00591f
C230 _31_/a_285_297# net10 1.68e-19
C231 _31_/a_35_297# _03_ 0.00749f
C232 _07_ _34_/a_47_47# 0.011f
C233 net12 _29_/a_111_297# 1.21e-19
C234 VPWR _36_/a_109_47# -4.66e-19
C235 net11 _21_ 0.586f
C236 VPWR _39_/a_47_47# 0.0668f
C237 VPWR net19 0.181f
C238 b[2] _21_ 2.14e-19
C239 input2/a_27_47# net8 0.0207f
C240 net11 net8 1.5e-19
C241 _10_ _25_ 0.0109f
C242 _42_/a_209_311# _37_/a_27_47# 1.59e-20
C243 _30_/a_109_53# p[3] 1.81e-20
C244 p[6] b[3] 0.184f
C245 net13 _08_ 1.82e-19
C246 _49_/a_544_297# net1 0.00175f
C247 _52_/a_93_21# net11 2.8e-19
C248 VGND net17 0.212f
C249 p[13] _44_/a_250_297# 4.09e-20
C250 _52_/a_250_297# _05_ 8.86e-22
C251 _52_/a_93_21# b[2] 1.63e-19
C252 _35_/a_226_47# net10 0.018f
C253 net1 net3 4.25e-20
C254 p[8] _43_/a_469_47# 2.83e-20
C255 net17 p[1] 6.65e-20
C256 _12_ net2 1.02e-20
C257 _32_/a_27_47# _20_ 0.0069f
C258 net12 p[5] 0.00302f
C259 net13 _02_ 0.00154f
C260 b[3] _14_ 1.92e-19
C261 net5 _44_/a_93_21# 3.61e-20
C262 p[2] net13 2.24e-19
C263 _44_/a_250_297# _16_ 3.25e-19
C264 _30_/a_215_297# _04_ 0.00225f
C265 _20_ _49_/a_201_297# 5.24e-21
C266 VGND net15 0.222f
C267 net15 _43_/a_193_413# 0.00169f
C268 net14 _43_/a_369_47# 6.79e-21
C269 VPWR input5/a_381_47# 8.33e-19
C270 _33_/a_109_93# _21_ 1.62e-20
C271 p[1] net15 6.22e-20
C272 _27_/a_277_297# net3 2.71e-19
C273 _06_ _35_/a_489_413# 9.22e-19
C274 _35_/a_226_297# _09_ 4.98e-19
C275 _31_/a_285_47# _05_ 5.61e-19
C276 p[2] input11/a_27_47# 1.02e-20
C277 _55_/a_80_21# net7 0.00163f
C278 net13 _33_/a_296_53# 3.71e-20
C279 p[3] net1 6.54e-19
C280 input12/a_27_47# b[1] 5.49e-19
C281 net8 net3 9.23e-19
C282 p[9] input14/a_27_47# 6.51e-20
C283 _52_/a_93_21# _33_/a_109_93# 2.89e-21
C284 _35_/a_76_199# _12_ 6.84e-20
C285 _31_/a_35_297# _02_ 0.00316f
C286 p[2] _31_/a_35_297# 0.00264f
C287 output16/a_27_47# _38_/a_27_47# 9.02e-19
C288 _14_ net4 1.54e-20
C289 VGND net10 0.456f
C290 VPWR output19/a_27_47# 0.0229f
C291 _35_/a_226_47# net11 3.21e-19
C292 p[3] _21_ 3.95e-21
C293 p[3] net8 0.0015f
C294 _55_/a_472_297# b[3] 1.51e-19
C295 _34_/a_285_47# b[1] 8.85e-20
C296 input13/a_27_47# _35_/a_226_47# 3.94e-20
C297 _04_ _19_ 0.356f
C298 _06_ net15 0.033f
C299 VGND _40_/a_297_297# -5.1e-19
C300 _42_/a_296_53# net3 1.81e-19
C301 net5 _25_ 6.42e-19
C302 p[8] input5/a_62_47# 1.15e-19
C303 _35_/a_226_47# _33_/a_109_93# 4.9e-19
C304 _35_/a_76_199# _33_/a_209_311# 9.95e-21
C305 _15_ _26_/a_183_297# 4.63e-36
C306 VPWR p[7] 0.023f
C307 VGND input2/a_27_47# -0.0137f
C308 VGND net11 0.475f
C309 p[1] input2/a_27_47# 0.0118f
C310 input7/a_27_47# p[10] 0.00138f
C311 VGND b[2] 0.0779f
C312 p[13] _01_ 2.02e-20
C313 net5 _52_/a_346_47# 7.03e-19
C314 _45_/a_27_47# _17_ 1.16e-20
C315 _34_/a_377_297# _04_ 1.7e-20
C316 _39_/a_377_297# p[12] 4.23e-19
C317 _06_ net10 0.184f
C318 VGND input13/a_27_47# 0.0471f
C319 net7 input5/a_664_47# 0.00199f
C320 _04_ _29_/a_183_297# 0.0015f
C321 _47_/a_384_47# VPWR -1.45e-19
C322 _32_/a_27_47# _00_ 0.00228f
C323 _01_ _16_ 3.24e-19
C324 output17/a_27_47# input5/a_62_47# 1.02e-19
C325 _12_ _13_ 0.462f
C326 net12 p[6] 0.0277f
C327 _16_ _22_ 3.8e-19
C328 _10_ input6/a_27_47# 4.57e-20
C329 _01_ _27_/a_27_297# 8.04e-19
C330 _40_/a_191_297# _14_ 2.4e-19
C331 _48_/a_27_47# net10 0.00377f
C332 _50_/a_343_93# p[12] 5.88e-21
C333 VGND _33_/a_109_93# -0.013f
C334 _31_/a_35_297# _55_/a_80_21# 5.9e-21
C335 net13 _34_/a_47_47# 1.68e-19
C336 VGND _49_/a_544_297# -0.00256f
C337 net18 p[5] 1.98e-19
C338 VGND net3 0.322f
C339 input12/a_27_47# _02_ 1.88e-19
C340 net3 _43_/a_193_413# 5.65e-20
C341 _06_ _40_/a_297_297# 1.64e-19
C342 p[2] input12/a_27_47# 1.02e-20
C343 _12_ _09_ 0.00526f
C344 VPWR _35_/a_226_297# -8.54e-19
C345 net8 net19 1.15e-19
C346 p[13] input5/a_62_47# 0.0215f
C347 _36_/a_303_47# net13 5.5e-20
C348 net1 input5/a_381_47# 1.27e-19
C349 VPWR input1/a_75_212# 0.0786f
C350 _15_ p[12] 0.0163f
C351 _34_/a_285_47# _08_ 0.00414f
C352 _06_ net11 0.546f
C353 net16 net18 0.00585f
C354 _52_/a_93_21# _39_/a_47_47# 1.44e-20
C355 _52_/a_250_297# _22_ 0.0996f
C356 _06_ b[2] 0.0116f
C357 _04_ _32_/a_27_47# 1.43e-19
C358 net9 _32_/a_109_47# 6.44e-19
C359 VGND p[3] 0.219f
C360 input13/a_27_47# _06_ 7.75e-19
C361 _31_/a_285_47# _01_ 3.36e-19
C362 p[3] p[1] 0.0145f
C363 _20_ _00_ 0.271f
C364 _04_ _49_/a_201_297# 0.0253f
C365 _34_/a_285_47# _02_ 7.14e-19
C366 input6/a_27_47# net14 7.05e-19
C367 p[8] p[11] 0.00173f
C368 _48_/a_27_47# net11 0.0179f
C369 net8 input5/a_381_47# 7.48e-19
C370 _10_ b[3] 3.27e-20
C371 _11_ net15 0.145f
C372 _44_/a_250_297# _14_ 4.82e-19
C373 net16 _22_ 0.00606f
C374 _37_/a_303_47# net14 0.00112f
C375 _06_ _33_/a_109_93# 9.13e-19
C376 _33_/a_209_311# _09_ 3.79e-20
C377 _23_ net9 1.21e-19
C378 _42_/a_296_53# net19 2.71e-19
C379 _06_ net3 0.0072f
C380 net3 _27_/a_205_297# 4.37e-19
C381 _19_ input7/a_27_47# 3.12e-21
C382 _50_/a_343_93# net2 1.25e-20
C383 _47_/a_299_297# p[12] 1.8e-19
C384 _45_/a_27_47# input4/a_75_212# 2.18e-20
C385 net2 input5/a_558_47# 5.99e-21
C386 _10_ net4 0.183f
C387 _18_ p[12] 1.89e-19
C388 input8/a_27_47# b[3] 1.21e-19
C389 _04_ _20_ 0.0677f
C390 VGND _49_/a_315_47# -0.0034f
C391 _39_/a_285_47# net4 9.71e-19
C392 _50_/a_223_47# _20_ 1.71e-19
C393 _06_ p[3] 1.59e-20
C394 b[3] net14 0.0194f
C395 _32_/a_197_47# _02_ 3.78e-19
C396 p[7] net1 7.5e-20
C397 net2 _15_ 9.8e-19
C398 _42_/a_209_311# input5/a_558_47# 7.85e-20
C399 _10_ _45_/a_193_297# 0.0047f
C400 VPWR _37_/a_27_47# -0.0178f
C401 _45_/a_27_47# _50_/a_27_47# 0.109f
C402 p[13] p[11] 0.023f
C403 _07_ net9 1.39e-20
C404 p[9] p[12] 1.4e-19
C405 net18 output18/a_27_47# 0.0106f
C406 _42_/a_209_311# _15_ 0.0521f
C407 VGND _36_/a_109_47# 3.56e-19
C408 _11_ _40_/a_297_297# 9.94e-19
C409 net13 input9/a_75_212# 4.4e-19
C410 VGND _39_/a_47_47# 0.0665f
C411 VGND net19 0.133f
C412 net19 _43_/a_193_413# 3.31e-19
C413 _14_ _43_/a_469_47# 0.00259f
C414 net14 net4 2.21e-21
C415 _34_/a_47_47# input12/a_27_47# 2.17e-19
C416 VPWR _12_ 0.28f
C417 _10_ _45_/a_465_47# 3.32e-19
C418 p[8] net15 0.0122f
C419 _22_ output18/a_27_47# 7.51e-19
C420 net5 b[3] 0.00347f
C421 _49_/a_75_199# _09_ 2.93e-19
C422 net2 _47_/a_299_297# 1.18e-19
C423 output17/a_27_47# net17 0.0149f
C424 VGND input5/a_381_47# -0.0034f
C425 input1/a_75_212# net1 0.00208f
C426 _01_ _14_ 0.0193f
C427 net2 _18_ 0.00181f
C428 b[1] _38_/a_197_47# 7.64e-20
C429 _14_ _22_ 0.00449f
C430 net6 p[12] 0.1f
C431 input6/a_27_47# _44_/a_93_21# 8.53e-19
C432 _42_/a_209_311# _18_ 3.21e-19
C433 _36_/a_109_47# _06_ 0.00168f
C434 net5 net4 0.0447f
C435 _11_ net3 0.165f
C436 _39_/a_47_47# _06_ 1.44e-19
C437 _06_ net19 0.00522f
C438 _37_/a_109_47# net3 0.00212f
C439 VPWR _33_/a_209_311# -0.0131f
C440 _10_ net12 0.00257f
C441 _10_ _05_ 9.25e-21
C442 _50_/a_343_93# _13_ 5.63e-20
C443 p[9] net2 0.00156f
C444 VGND output19/a_27_47# -0.00902f
C445 _42_/a_109_93# _17_ 7.83e-20
C446 _35_/a_226_47# p[7] 2.82e-19
C447 _35_/a_76_199# _18_ 6.82e-21
C448 p[0] b[1] 0.0562f
C449 net9 net7 0.00233f
C450 _04_ _00_ 1.98e-20
C451 _30_/a_297_297# net10 1.68e-19
C452 net5 _45_/a_193_297# 0.00935f
C453 net10 output17/a_27_47# 1.31e-20
C454 _50_/a_223_47# _00_ 0.00738f
C455 _45_/a_109_297# net6 7.82e-19
C456 p[13] net15 8.62e-19
C457 p[8] _40_/a_297_297# 1.12e-19
C458 _42_/a_209_311# p[9] 5.51e-21
C459 _01_ _55_/a_472_297# 6.28e-19
C460 _16_ net15 0.214f
C461 _15_ _13_ 3.69e-20
C462 _27_/a_27_297# net17 0.00181f
C463 _06_ input5/a_381_47# 1.6e-19
C464 input15/a_27_47# input6/a_27_47# 5.3e-19
C465 input8/a_27_47# _05_ 1.58e-19
C466 _24_ _12_ 1.67e-19
C467 _27_/a_27_297# net15 0.00888f
C468 b[3] _44_/a_93_21# 0.00491f
C469 input5/a_841_47# net9 2.7e-19
C470 VGND p[7] 0.198f
C471 p[10] net7 0.00546f
C472 _12_ _38_/a_303_47# 0.00153f
C473 _30_/a_392_297# net12 2.19e-20
C474 output17/a_27_47# input2/a_27_47# 0.107f
C475 net2 net6 0.00139f
C476 VGND _47_/a_384_47# -2.05e-19
C477 _06_ output19/a_27_47# 1.53e-19
C478 _50_/a_223_47# _04_ 7.89e-22
C479 _31_/a_285_47# net17 0.00134f
C480 b[1] net2 0.0189f
C481 _31_/a_117_297# b[1] 1.45e-19
C482 _29_/a_29_53# _49_/a_75_199# 1.28e-19
C483 p[8] net3 0.00454f
C484 _37_/a_27_47# net8 6.66e-21
C485 _42_/a_209_311# net6 1.32e-20
C486 net13 net9 0.035f
C487 VPWR _49_/a_75_199# 0.0177f
C488 _44_/a_250_297# net14 4.24e-20
C489 _52_/a_250_297# net10 2.86e-21
C490 _13_ _18_ 0.019f
C491 input15/a_27_47# b[3] 1.77e-19
C492 _50_/a_27_47# net13 7.27e-21
C493 _35_/a_76_199# net6 4.6e-21
C494 p[4] b[3] 0.0504f
C495 net5 net12 0.0674f
C496 _35_/a_76_199# b[1] 5.2e-21
C497 net10 p[5] 0.00814f
C498 VGND _35_/a_226_297# -4.55e-19
C499 _02_ p[12] 0.00185f
C500 output17/a_27_47# net3 0.00248f
C501 VGND input1/a_75_212# 0.0581f
C502 _12_ _21_ 7.99e-20
C503 _49_/a_208_47# net7 0.00312f
C504 _06_ p[7] 0.00874f
C505 _09_ _18_ 7.01e-21
C506 _11_ net19 2.19e-19
C507 _39_/a_47_47# _11_ 3.9e-19
C508 input1/a_75_212# p[1] 0.0023f
C509 _31_/a_117_297# _03_ 5.32e-19
C510 _03_ net2 1.89e-19
C511 _10_ _43_/a_469_47# 0.00124f
C512 _37_/a_109_47# net19 1.16e-20
C513 _07_ _34_/a_377_297# 5.8e-19
C514 net11 _29_/a_111_297# 8.27e-19
C515 _25_ b[3] 5.83e-19
C516 _27_/a_27_297# input2/a_27_47# 1.16e-19
C517 VPWR _36_/a_197_47# -5.24e-19
C518 _27_/a_27_297# net11 1.58e-20
C519 _52_/a_93_21# _12_ 0.0157f
C520 _30_/a_297_297# p[3] 1.74e-20
C521 _45_/a_109_297# _02_ 8.44e-19
C522 _50_/a_615_93# _20_ 8.8e-19
C523 _01_ _47_/a_81_21# 6.05e-21
C524 _52_/a_250_297# net11 1.2e-19
C525 net5 _44_/a_250_297# 3.11e-20
C526 p[13] net3 8.64e-19
C527 _35_/a_76_199# _03_ 0.0733f
C528 _52_/a_250_297# b[2] 1.6e-19
C529 _10_ _01_ 2.22e-19
C530 VPWR _50_/a_343_93# -0.0126f
C531 net11 p[5] 0.0857f
C532 _16_ net3 1.77e-19
C533 _22_ _47_/a_81_21# 7.25e-19
C534 net14 _43_/a_469_47# 1.44e-20
C535 _10_ _36_/a_27_47# 0.00109f
C536 VPWR input5/a_558_47# 0.0083f
C537 b[0] output16/a_27_47# 0.0228f
C538 _10_ _22_ 0.0904f
C539 _06_ _35_/a_226_297# 1.28e-19
C540 input13/a_27_47# p[5] 3.09e-19
C541 _35_/a_556_47# _09_ 0.00122f
C542 _31_/a_35_297# p[10] 2.29e-19
C543 _19_ net7 0.0458f
C544 _27_/a_27_297# net3 0.0133f
C545 _55_/a_217_297# net7 1.04e-19
C546 net13 _33_/a_368_53# 2.1e-20
C547 net16 net11 4.43e-22
C548 VPWR _15_ 0.912f
C549 _52_/a_250_297# _33_/a_109_93# 5.17e-22
C550 _42_/a_109_93# p[10] 1.82e-21
C551 _35_/a_226_47# _12_ 8.38e-20
C552 net6 _13_ 0.0106f
C553 input8/a_27_47# _01_ 1.43e-19
C554 _30_/a_215_297# net13 0.0246f
C555 b[1] _13_ 2.71e-21
C556 VGND _37_/a_27_47# -0.0147f
C557 _37_/a_27_47# _43_/a_193_413# 0.0102f
C558 input11/a_27_47# input10/a_27_47# 5.3e-19
C559 net17 _14_ 2.4e-20
C560 _01_ net14 8.29e-19
C561 p[8] net19 0.0358f
C562 _35_/a_76_199# _08_ 0.0061f
C563 _42_/a_209_311# _02_ 9.92e-19
C564 net6 _09_ 5.43e-20
C565 net2 _43_/a_27_47# 0.01f
C566 _14_ net15 0.0538f
C567 _22_ net14 2.23e-19
C568 _35_/a_76_199# _02_ 5.73e-19
C569 _31_/a_35_297# _30_/a_215_297# 6.37e-19
C570 _10_ _45_/a_205_47# 6.19e-20
C571 net10 p[6] 0.00668f
C572 VGND _12_ 0.816f
C573 _52_/a_256_47# net10 8.13e-20
C574 net1 _49_/a_75_199# 0.00799f
C575 _12_ _43_/a_193_413# 7.94e-22
C576 _42_/a_368_53# net3 3.82e-19
C577 VPWR _47_/a_299_297# 0.0643f
C578 _44_/a_250_297# _44_/a_93_21# -6.97e-22
C579 _03_ _13_ 1.74e-20
C580 _35_/a_226_47# _33_/a_209_311# 1.31e-19
C581 _07_ _20_ 1.28e-21
C582 p[4] net12 6.15e-19
C583 VPWR _18_ 0.0721f
C584 net14 input5/a_62_47# 5.28e-20
C585 _47_/a_384_47# _11_ 7.23e-20
C586 net13 _19_ 4.45e-20
C587 net5 _52_/a_584_47# 0.0022f
C588 net5 _01_ 0.0779f
C589 _49_/a_75_199# _21_ 6.64e-19
C590 _03_ _09_ 0.326f
C591 _06_ _37_/a_27_47# 2.5e-20
C592 _44_/a_346_47# _17_ 7.2e-19
C593 net8 _49_/a_75_199# 0.00214f
C594 _04_ input3/a_27_47# 3.55e-19
C595 _40_/a_109_297# net6 2.53e-20
C596 net5 _36_/a_27_47# 0.0163f
C597 _32_/a_27_47# net7 0.00559f
C598 output17/a_27_47# input5/a_381_47# 6.6e-20
C599 _25_ net12 4.46e-20
C600 net5 _22_ 0.405f
C601 input6/a_27_47# b[3] 4.02e-19
C602 net11 output18/a_27_47# 6.84e-20
C603 p[8] output19/a_27_47# 0.035f
C604 _49_/a_201_297# net7 0.00419f
C605 b[2] output18/a_27_47# 0.0141f
C606 VPWR p[9] 0.41f
C607 net11 p[6] 0.0126f
C608 _16_ net19 0.206f
C609 _31_/a_35_297# _19_ 1.47e-19
C610 _40_/a_297_297# _14_ 1.58e-19
C611 _50_/a_429_93# p[12] 3.96e-20
C612 VGND _33_/a_209_311# -0.00669f
C613 input13/a_27_47# p[6] 1.07e-19
C614 _27_/a_27_297# net19 1.98e-19
C615 _06_ _12_ 0.136f
C616 _42_/a_109_93# _19_ 1.14e-21
C617 VPWR _35_/a_556_47# -7.24e-19
C618 net5 input5/a_62_47# 0.00329f
C619 p[13] input5/a_381_47# 0.00214f
C620 _42_/a_209_311# _55_/a_80_21# 0.0175f
C621 net1 input5/a_558_47# 1.1e-19
C622 _02_ _13_ 0.0676f
C623 _53_/a_29_53# _13_ 9.05e-19
C624 _29_/a_29_53# _26_/a_29_53# 0.00121f
C625 _08_ _09_ 0.106f
C626 net9 _32_/a_197_47# 6.06e-19
C627 input12/a_27_47# input10/a_27_47# 0.0154f
C628 net5 _45_/a_205_47# 8.28e-20
C629 _29_/a_29_53# net6 1.4e-20
C630 _20_ net7 0.0257f
C631 _50_/a_343_93# net8 7.25e-19
C632 _02_ _09_ 0.297f
C633 VPWR _26_/a_29_53# 0.0356f
C634 _29_/a_29_53# b[1] 1.49e-21
C635 _53_/a_29_53# _09_ 0.00642f
C636 _27_/a_27_297# input5/a_381_47# 1.47e-19
C637 _35_/a_226_47# _49_/a_75_199# 8.73e-20
C638 _43_/a_27_47# _13_ 1.66e-20
C639 _45_/a_27_47# _00_ 4.84e-20
C640 net8 input5/a_558_47# 0.00357f
C641 _47_/a_384_47# p[8] 1.34e-20
C642 _10_ _35_/a_489_413# 3.41e-19
C643 VPWR net6 0.999f
C644 p[11] net14 1.32e-19
C645 VPWR b[1] 0.621f
C646 _14_ net3 0.0295f
C647 net16 _39_/a_47_47# 7.7e-20
C648 _15_ _21_ 1.13e-21
C649 _37_/a_197_47# net15 1.78e-19
C650 _06_ _33_/a_209_311# 0.0187f
C651 net8 _15_ 1.79e-19
C652 VPWR _54_/a_75_212# 0.0475f
C653 net13 _49_/a_201_297# 3.31e-19
C654 _42_/a_368_53# net19 5.12e-19
C655 net2 input5/a_664_47# 8.11e-20
C656 _29_/a_29_53# _03_ 0.0414f
C657 VGND _49_/a_75_199# 5.87e-20
C658 _31_/a_35_297# _32_/a_27_47# 9.17e-20
C659 _11_ _37_/a_27_47# 0.0018f
C660 m1_7039_1799# p[5] 4.89e-20
C661 _31_/a_35_297# _49_/a_201_297# 5.52e-20
C662 _32_/a_303_47# _02_ 1.15e-20
C663 _42_/a_209_311# input5/a_664_47# 0.0124f
C664 net15 _47_/a_81_21# 0.00106f
C665 VPWR _03_ 0.845f
C666 _44_/a_93_21# input5/a_62_47# 5.05e-20
C667 _10_ net15 0.0101f
C668 _25_ net18 0.0594f
C669 _07_ _04_ 9.74e-20
C670 _42_/a_296_53# _15_ 1.28e-19
C671 net13 _20_ 5.95e-19
C672 VGND _36_/a_197_47# -3.75e-19
C673 input1/a_75_212# output17/a_27_47# 0.0101f
C674 _11_ _12_ 0.195f
C675 VGND _39_/a_377_297# -6.28e-19
C676 _48_/a_109_47# net11 1.74e-19
C677 _45_/a_193_297# net4 7.41e-19
C678 net8 _18_ 1.15e-21
C679 _17_ _45_/a_109_297# 4.29e-22
C680 _24_ _26_/a_29_53# 2.11e-20
C681 _10_ net10 4.45e-19
C682 net17 net14 5.43e-19
C683 _36_/a_27_47# _25_ 2.34e-20
C684 _52_/a_93_21# _18_ 1.97e-19
C685 _24_ net6 0.00121f
C686 _25_ _22_ 5.39e-19
C687 _31_/a_35_297# _20_ 1.69e-19
C688 _00_ net7 8.12e-21
C689 _24_ b[1] 6.01e-20
C690 VGND _50_/a_343_93# -4.3e-19
C691 p[7] p[5] 1.29e-19
C692 _29_/a_29_53# _02_ 6.76e-21
C693 net14 net15 1.07f
C694 VPWR _08_ -0.0171f
C695 _30_/a_109_53# b[1] 2.69e-20
C696 p[13] input1/a_75_212# 4.16e-19
C697 VGND input5/a_558_47# -0.00123f
C698 p[1] input5/a_558_47# 1.61e-21
C699 b[1] _38_/a_303_47# 8.14e-20
C700 VPWR _02_ 0.332f
C701 VPWR _53_/a_29_53# 0.00821f
C702 p[2] VPWR 0.121f
C703 p[8] _37_/a_27_47# 0.0017f
C704 _35_/a_556_47# _21_ 2.69e-19
C705 VGND _15_ 0.149f
C706 _17_ net2 0.181f
C707 _14_ net19 0.00714f
C708 _15_ _43_/a_193_413# 4.86e-19
C709 net12 b[3] 2.47e-19
C710 _12_ _39_/a_129_47# 0.00175f
C711 _36_/a_197_47# _06_ 6.18e-19
C712 _37_/a_197_47# net3 0.0028f
C713 _39_/a_377_297# _06_ 8.76e-20
C714 VPWR _33_/a_296_53# -1.15e-19
C715 _10_ net11 0.0109f
C716 p[14] p[12] 0.00101f
C717 _24_ _03_ 9.46e-20
C718 _42_/a_209_311# _17_ 1.22e-19
C719 net5 net17 4.21e-21
C720 VPWR _43_/a_27_47# 0.0186f
C721 net1 b[1] 0.00429f
C722 _04_ net7 0.0602f
C723 _30_/a_109_53# _03_ 0.0189f
C724 _30_/a_392_297# net10 3.4e-19
C725 net5 net15 0.0226f
C726 input4/a_75_212# p[12] 0.026f
C727 _12_ p[8] 2.09e-20
C728 _14_ input5/a_381_47# 5.68e-20
C729 _50_/a_343_93# _06_ 0.0376f
C730 net6 _21_ 2.92e-20
C731 _01_ _55_/a_300_47# 0.00113f
C732 net12 net4 2.57e-20
C733 b[1] _21_ 0.00179f
C734 _06_ input5/a_558_47# 3.55e-19
C735 b[1] net8 0.00199f
C736 _55_/a_300_47# _22_ 2.08e-19
C737 VGND _47_/a_299_297# -3.63e-19
C738 _44_/a_250_297# b[3] 0.0112f
C739 _47_/a_81_21# net3 6.66e-19
C740 _52_/a_93_21# net6 2.33e-19
C741 _45_/a_193_297# _05_ 4.84e-22
C742 input2/a_27_47# net14 0.0102f
C743 _50_/a_27_47# p[12] 1.93e-19
C744 _10_ net3 3.89e-19
C745 net5 net10 0.0316f
C746 net11 net14 9.95e-19
C747 _06_ _15_ 0.22f
C748 _15_ _27_/a_205_297# 5.5e-20
C749 VGND _18_ 0.0166f
C750 _43_/a_193_413# _18_ 0.0413f
C751 _03_ net1 0.298f
C752 _14_ output19/a_27_47# 1.43e-19
C753 _16_ _37_/a_27_47# 2.07e-19
C754 _30_/a_465_297# net12 8.01e-20
C755 _03_ _27_/a_277_297# 2.1e-20
C756 _24_ _02_ 0.0232f
C757 _31_/a_285_297# b[1] 8.82e-20
C758 _24_ _53_/a_29_53# 0.0835f
C759 _10_ p[3] 1.37e-20
C760 _03_ _21_ 0.0818f
C761 _30_/a_109_53# _02_ 5.03e-22
C762 VGND p[9] 0.0807f
C763 net2 p[14] 1.38e-19
C764 VPWR _55_/a_80_21# 0.0289f
C765 p[7] p[6] 0.768f
C766 p[9] _43_/a_193_413# 1.09e-19
C767 _03_ net8 0.0287f
C768 net13 _04_ 0.569f
C769 net14 net3 0.684f
C770 _52_/a_93_21# _03_ 0.00985f
C771 _42_/a_209_311# p[14] 3.45e-22
C772 net5 net11 0.0129f
C773 _06_ _47_/a_299_297# 0.0174f
C774 p[0] p[10] 0.015f
C775 _35_/a_226_47# b[1] 1.46e-22
C776 VGND _35_/a_556_47# 1.95e-19
C777 net15 _44_/a_93_21# 0.00573f
C778 net5 b[2] 7.33e-20
C779 VPWR _34_/a_47_47# 0.0372f
C780 input8/a_27_47# p[3] 0.0023f
C781 _06_ _18_ 0.54f
C782 _39_/a_377_297# _11_ 2.57e-20
C783 net9 net2 3.64e-20
C784 _31_/a_285_297# _03_ 0.00677f
C785 _31_/a_35_297# _04_ 1.89e-20
C786 net1 _02_ 0.00251f
C787 p[2] net1 0.0269f
C788 net18 b[3] 7.1e-19
C789 VPWR _36_/a_303_47# -4.83e-19
C790 _41_/a_59_75# p[12] 0.0562f
C791 _08_ _21_ 0.00139f
C792 VGND _26_/a_29_53# 0.0381f
C793 _52_/a_250_297# _12_ 0.0139f
C794 net12 _05_ 0.0414f
C795 _28_/a_109_297# _15_ 0.00346f
C796 _42_/a_109_93# _04_ 5.77e-22
C797 net2 _27_/a_109_297# 7.24e-20
C798 _50_/a_343_93# _11_ 0.0384f
C799 VGND net6 0.472f
C800 net6 _43_/a_193_413# 2.41e-20
C801 _06_ p[9] 0.00205f
C802 _53_/a_29_53# _21_ 0.00959f
C803 _02_ _21_ 0.397f
C804 _01_ b[3] 1.98e-19
C805 input7/a_27_47# net7 0.00318f
C806 net5 net3 0.0365f
C807 VGND b[1] 1.54f
C808 _35_/a_226_47# _03_ 0.028f
C809 net8 _02_ 0.334f
C810 p[2] net8 0.00871f
C811 b[1] p[1] 0.0426f
C812 input15/a_27_47# net15 0.00325f
C813 VPWR _50_/a_429_93# -3.61e-19
C814 b[3] _22_ 1.28e-19
C815 VGND _54_/a_75_212# 0.053f
C816 _52_/a_93_21# _02_ 0.0962f
C817 net16 _12_ 0.131f
C818 _52_/a_93_21# _53_/a_29_53# 0.00116f
C819 VPWR input5/a_664_47# 0.00488f
C820 _10_ net19 0.00224f
C821 _10_ _39_/a_47_47# 0.00824f
C822 _11_ _15_ 0.113f
C823 net2 p[10] 0.0638f
C824 _40_/a_109_297# _17_ 9.67e-19
C825 _42_/a_209_311# p[10] 2.37e-20
C826 _31_/a_285_297# _02_ 5.86e-20
C827 p[2] _31_/a_285_297# 0.00155f
C828 _36_/a_27_47# net4 0.0103f
C829 p[4] net10 0.00279f
C830 _22_ net4 0.0866f
C831 b[3] input5/a_62_47# 0.00532f
C832 _06_ _26_/a_29_53# 0.0135f
C833 VGND _03_ 0.121f
C834 _45_/a_27_47# _23_ 1.74e-19
C835 _24_ _34_/a_47_47# 6.84e-21
C836 _35_/a_226_47# _08_ 0.00117f
C837 output16/a_27_47# p[12] 0.00102f
C838 _06_ net6 0.308f
C839 _45_/a_193_297# _22_ 0.0234f
C840 _06_ b[1] 0.00237f
C841 net19 net14 0.148f
C842 _25_ net10 2.66e-19
C843 _29_/a_29_53# input9/a_75_212# 9.7e-21
C844 _23_ _07_ 1.27e-19
C845 _35_/a_226_47# _02_ 2.21e-19
C846 _11_ _47_/a_299_297# 0.00738f
C847 net1 _55_/a_80_21# 1.8e-19
C848 _06_ _54_/a_75_212# 0.00727f
C849 _50_/a_343_93# p[8] 1.03e-20
C850 _11_ _18_ 0.484f
C851 VPWR input9/a_75_212# 0.0641f
C852 _48_/a_27_47# b[1] 5.84e-19
C853 net3 _44_/a_93_21# 0.0102f
C854 _10_ output19/a_27_47# 3.23e-20
C855 p[4] net11 0.0556f
C856 _50_/a_27_47# _13_ 0.00169f
C857 _45_/a_27_47# _07_ 1.02e-20
C858 _37_/a_27_47# _14_ 0.00137f
C859 net14 input5/a_381_47# 0.00479f
C860 VGND _08_ 0.162f
C861 net8 _55_/a_80_21# 1.84e-21
C862 p[8] _15_ 0.00832f
C863 p[4] input13/a_27_47# 7.37e-20
C864 _27_/a_27_297# _49_/a_75_199# 0.011f
C865 _06_ _03_ 0.00635f
C866 VPWR _17_ 0.306f
C867 net9 _09_ 2.62e-19
C868 _03_ _27_/a_205_297# 1.46e-20
C869 _11_ p[9] 1.01e-19
C870 VGND _02_ 1.63f
C871 VGND _53_/a_29_53# -0.0168f
C872 p[2] VGND 0.136f
C873 _02_ _43_/a_193_413# 9.4e-21
C874 net5 _36_/a_109_47# 0.00144f
C875 _55_/a_300_47# net15 1.09e-19
C876 _50_/a_27_47# _09_ 1.3e-19
C877 _25_ net11 0.0262f
C878 net5 net19 0.00124f
C879 p[2] p[1] 0.121f
C880 net5 _39_/a_47_47# 0.0389f
C881 _25_ b[2] 0.0015f
C882 _34_/a_47_47# _21_ 8.93e-19
C883 _19_ net2 0.101f
C884 _50_/a_515_93# p[12] 6.6e-20
C885 _12_ _14_ 1.98e-20
C886 net14 output19/a_27_47# 0.00142f
C887 p[11] b[3] 0.157f
C888 VGND _33_/a_296_53# -1.43e-19
C889 input15/a_27_47# net3 8.74e-20
C890 _01_ net12 1.67e-21
C891 _01_ _05_ 5.03e-19
C892 VGND _43_/a_27_47# -0.0153f
C893 _36_/a_27_47# net12 0.0185f
C894 _36_/a_27_47# _05_ 3.67e-21
C895 net12 _22_ 5.73e-20
C896 _05_ _22_ 3.33e-21
C897 _10_ _47_/a_384_47# 3.53e-19
C898 net5 input5/a_381_47# 0.0546f
C899 p[13] input5/a_558_47# 0.0019f
C900 net1 input5/a_664_47# 2.41e-19
C901 p[8] _47_/a_299_297# 1.03e-19
C902 _11_ _26_/a_29_53# 1.09e-19
C903 _06_ _08_ 0.0343f
C904 net9 _32_/a_303_47# 0.00218f
C905 p[8] _18_ 1.68e-19
C906 _11_ net6 0.0257f
C907 input6/a_27_47# net15 0.00115f
C908 _06_ _53_/a_29_53# 0.0709f
C909 _06_ _02_ 0.85f
C910 _53_/a_111_297# _09_ 3.4e-19
C911 VPWR _26_/a_111_297# -5.92e-20
C912 _21_ input5/a_664_47# 9.42e-22
C913 _27_/a_27_297# input5/a_558_47# 1.57e-19
C914 _11_ b[1] 0.00239f
C915 _16_ _15_ 0.0607f
C916 net8 input5/a_664_47# 0.0116f
C917 _48_/a_27_47# _08_ 2.58e-19
C918 _11_ _54_/a_75_212# 3.22e-20
C919 _42_/a_109_93# input3/a_27_47# 0.00249f
C920 _27_/a_27_297# _15_ 9.85e-20
C921 _37_/a_303_47# net15 0.00118f
C922 p[9] p[8] 0.0807f
C923 _06_ _33_/a_296_53# 1.11e-20
C924 _48_/a_27_47# _53_/a_29_53# 3.14e-21
C925 _48_/a_27_47# _02_ 0.00435f
C926 _06_ _43_/a_27_47# 0.0329f
C927 VPWR p[14] 0.0425f
C928 net19 _44_/a_93_21# 0.0074f
C929 VGND _55_/a_80_21# 0.00281f
C930 _55_/a_80_21# _43_/a_193_413# 2.54e-19
C931 _49_/a_208_47# _09_ 5.43e-21
C932 VPWR input4/a_75_212# 0.06f
C933 _29_/a_29_53# net9 0.0205f
C934 net17 b[3] 0.00284f
C935 input9/a_75_212# net1 0.002f
C936 _44_/a_250_297# input5/a_62_47# 2.45e-20
C937 _29_/a_29_53# _50_/a_27_47# 1.44e-20
C938 _23_ net13 4.11e-19
C939 _39_/a_129_47# net6 6.91e-19
C940 b[3] net15 0.00608f
C941 VPWR net9 0.5f
C942 VGND _34_/a_47_47# 0.0901f
C943 _16_ _18_ 0.144f
C944 input9/a_75_212# _21_ 1.17e-21
C945 VPWR _50_/a_27_47# -0.00335f
C946 _00_ _26_/a_183_297# 4.53e-19
C947 net5 _47_/a_384_47# 0.00129f
C948 output16/a_27_47# _13_ 4.58e-19
C949 input15/a_27_47# net19 0.00236f
C950 p[8] net6 0.0062f
C951 VGND _36_/a_303_47# 8.14e-19
C952 VPWR _27_/a_109_297# -2.45e-19
C953 net10 b[3] 9.16e-20
C954 net15 net4 8.68e-19
C955 _19_ _09_ 4.8e-21
C956 _14_ _49_/a_75_199# 6.79e-20
C957 output19/a_27_47# _44_/a_93_21# 7.25e-20
C958 _06_ _55_/a_80_21# 5.15e-19
C959 _52_/a_250_297# _18_ 1.77e-19
C960 _17_ net8 4.52e-20
C961 _36_/a_109_47# _25_ 3.76e-21
C962 _07_ net13 0.00686f
C963 net18 _22_ 1.68e-19
C964 net2 _20_ 8.83e-19
C965 VGND _50_/a_429_93# 4.71e-19
C966 VPWR p[10] 0.218f
C967 _11_ _02_ 0.0621f
C968 _11_ _53_/a_29_53# 2.33e-20
C969 output17/a_27_47# b[1] 0.00756f
C970 VGND input5/a_664_47# 0.0134f
C971 _52_/a_584_47# _22_ 6.24e-19
C972 p[1] input5/a_664_47# 1.21e-20
C973 _01_ _22_ 0.15f
C974 _42_/a_209_311# _20_ 1.66e-20
C975 net10 net4 8.28e-22
C976 _06_ _34_/a_47_47# 0.0391f
C977 input6/a_27_47# net3 2.52e-19
C978 _12_ _47_/a_81_21# 0.00158f
C979 _36_/a_27_47# _22_ 2.82e-20
C980 net16 _18_ 8.17e-21
C981 _29_/a_183_297# _09_ 4.51e-20
C982 p[4] m1_7039_1799# 7.19e-19
C983 _10_ _12_ 0.19f
C984 _35_/a_76_199# _20_ 3.21e-20
C985 _00_ p[12] 9.97e-23
C986 _35_/a_489_413# net12 3.97e-20
C987 input2/a_27_47# b[3] 3.24e-19
C988 _11_ _43_/a_27_47# 4.27e-19
C989 net11 b[3] 0.00388f
C990 _12_ _39_/a_285_47# 0.0221f
C991 _36_/a_303_47# _06_ 5.3e-19
C992 _29_/a_29_53# _30_/a_215_297# 1.72e-19
C993 b[2] b[3] 0.0815f
C994 _37_/a_27_47# net14 0.0584f
C995 _37_/a_303_47# net3 0.00133f
C996 input5/a_841_47# net7 0.00193f
C997 VPWR _41_/a_59_75# 0.0179f
C998 VPWR _33_/a_368_53# -4.26e-19
C999 _48_/a_27_47# _34_/a_47_47# 4.45e-21
C1000 _38_/a_27_47# p[12] 5.26e-19
C1001 p[13] b[1] 0.00115f
C1002 input13/a_27_47# b[3] 1.21e-19
C1003 VPWR input10/a_27_47# 0.00986f
C1004 _16_ net6 1.62e-20
C1005 _30_/a_109_53# net9 0.0193f
C1006 _50_/a_343_93# _14_ 9.76e-19
C1007 _30_/a_297_297# _03_ 0.00117f
C1008 _30_/a_465_297# net10 0.00106f
C1009 VPWR _30_/a_215_297# -0.00472f
C1010 _03_ output17/a_27_47# 1.95e-19
C1011 _45_/a_109_297# _00_ 4.86e-20
C1012 VPWR _49_/a_208_47# -5.93e-19
C1013 input14/a_27_47# input3/a_27_47# 5.08e-20
C1014 _50_/a_429_93# _06_ 0.00169f
C1015 _33_/a_109_93# b[3] 1.86e-20
C1016 _27_/a_27_297# b[1] 7.43e-22
C1017 _40_/a_191_297# net15 8.41e-19
C1018 _06_ input5/a_664_47# 3.21e-19
C1019 _28_/a_109_297# _55_/a_80_21# 2.05e-20
C1020 net12 net17 2.11e-21
C1021 VGND input9/a_75_212# 0.0654f
C1022 net17 _05_ 0.0111f
C1023 _15_ _14_ 0.148f
C1024 b[3] net3 0.00853f
C1025 net13 net7 1.72e-19
C1026 _52_/a_250_297# net6 0.00133f
C1027 p[4] p[7] 0.127f
C1028 _49_/a_201_297# _09_ 1.74e-20
C1029 _50_/a_223_47# p[12] 2.36e-20
C1030 net5 _37_/a_27_47# 1.13e-20
C1031 net9 net1 0.47f
C1032 p[5] b[1] 0.256f
C1033 VGND _17_ 0.312f
C1034 p[3] b[3] 0.104f
C1035 net2 _00_ 0.00732f
C1036 _17_ _43_/a_193_413# 0.0503f
C1037 _31_/a_35_297# net7 0.0384f
C1038 _03_ _29_/a_111_297# 7.48e-19
C1039 net3 net4 9.28e-21
C1040 _24_ _53_/a_111_297# 9.08e-21
C1041 VPWR _19_ 0.0335f
C1042 net16 net6 8.27e-20
C1043 _20_ _13_ 7.38e-21
C1044 VPWR output16/a_27_47# 0.122f
C1045 net9 _21_ 0.0282f
C1046 _27_/a_27_297# _03_ 2.68e-19
C1047 p[8] _43_/a_27_47# 8.91e-20
C1048 VPWR _55_/a_217_297# -0.00133f
C1049 net16 b[1] 0.0107f
C1050 net10 net12 0.539f
C1051 net10 _05_ 0.457f
C1052 net9 net8 0.0605f
C1053 _50_/a_27_47# _21_ 3.38e-21
C1054 net5 _12_ 0.983f
C1055 _55_/a_472_297# _15_ 0.00626f
C1056 net16 _54_/a_75_212# 1.69e-21
C1057 _44_/a_250_297# net15 8.86e-20
C1058 _20_ _09_ 7.11e-19
C1059 input6/a_27_47# net19 0.00586f
C1060 _14_ _18_ 0.243f
C1061 net1 p[10] 0.00236f
C1062 VPWR _34_/a_377_297# -0.00192f
C1063 p[11] _22_ 3.13e-20
C1064 VPWR _29_/a_183_297# -8.13e-19
C1065 _04_ net2 0.158f
C1066 _31_/a_285_47# _03_ 8.54e-19
C1067 p[13] _02_ 5.96e-20
C1068 _07_ _34_/a_285_47# 0.00975f
C1069 _17_ _06_ 0.0341f
C1070 _16_ _02_ 0.00564f
C1071 VGND _26_/a_111_297# -2.75e-19
C1072 p[9] _14_ 2.62e-21
C1073 input2/a_27_47# _05_ 1.83e-19
C1074 p[10] net8 0.00987f
C1075 net12 net11 0.358f
C1076 net11 _05_ 2.76e-19
C1077 _42_/a_209_311# _04_ 9.84e-22
C1078 p[12] _41_/a_145_75# 0.00411f
C1079 _37_/a_27_47# _44_/a_93_21# 3.19e-19
C1080 _27_/a_27_297# _02_ 0.00179f
C1081 net6 _43_/a_297_47# 8.23e-22
C1082 _53_/a_111_297# _21_ 4.38e-19
C1083 input13/a_27_47# net12 0.0163f
C1084 p[11] input5/a_62_47# 0.00153f
C1085 input13/a_27_47# _05_ 3.93e-19
C1086 _31_/a_35_297# net13 1.86e-20
C1087 _35_/a_226_47# net9 1.22e-20
C1088 _35_/a_76_199# _04_ 0.0269f
C1089 _40_/a_109_297# _20_ 2.35e-20
C1090 _16_ _43_/a_27_47# 2.47e-19
C1091 _32_/a_303_47# _20_ 1.54e-19
C1092 _30_/a_215_297# net1 0.00375f
C1093 VPWR _50_/a_515_93# -5.03e-19
C1094 VGND p[14] 0.365f
C1095 b[3] net19 0.0439f
C1096 _40_/a_191_297# net3 1.89e-19
C1097 _52_/a_250_297# _02_ 0.0128f
C1098 net15 _43_/a_469_47# 7.41e-19
C1099 _10_ _36_/a_197_47# 1.54e-19
C1100 input8/a_27_47# _49_/a_75_199# 1.99e-20
C1101 _10_ _39_/a_377_297# 7.42e-19
C1102 input6/a_27_47# output19/a_27_47# 0.107f
C1103 VPWR _32_/a_27_47# 0.0395f
C1104 _33_/a_109_93# net12 0.0435f
C1105 _37_/a_197_47# _15_ 3.02e-19
C1106 _33_/a_109_93# _05_ 0.0206f
C1107 b[1] output18/a_27_47# 0.0028f
C1108 p[2] p[5] 3.27e-20
C1109 VGND input4/a_75_212# 0.0529f
C1110 _49_/a_75_199# net14 3.67e-19
C1111 VPWR _49_/a_201_297# 0.0185f
C1112 _30_/a_215_297# _21_ 1.48e-19
C1113 p[6] b[1] 0.0464f
C1114 _54_/a_75_212# output18/a_27_47# 2.28e-19
C1115 _14_ _26_/a_29_53# 3.67e-19
C1116 _30_/a_215_297# net8 8.14e-21
C1117 _00_ _13_ 3.77e-20
C1118 _50_/a_343_93# _47_/a_81_21# 0.00282f
C1119 _01_ net17 0.0988f
C1120 input15/a_27_47# _37_/a_27_47# 3.27e-19
C1121 net8 _49_/a_208_47# 1.4e-19
C1122 b[1] _48_/a_181_47# 4.99e-20
C1123 b[3] input5/a_381_47# 7.71e-19
C1124 p[0] input7/a_27_47# 5.13e-20
C1125 _10_ _50_/a_343_93# 0.0284f
C1126 _39_/a_47_47# net4 0.0202f
C1127 net19 net4 2.65e-20
C1128 _14_ net6 2.11e-19
C1129 _06_ _26_/a_111_297# 9e-19
C1130 net16 _02_ 8.94e-19
C1131 VGND net9 0.379f
C1132 net16 _53_/a_29_53# 2.04e-20
C1133 _01_ net15 0.0314f
C1134 _38_/a_27_47# _13_ 4.58e-19
C1135 VGND _50_/a_27_47# -0.00433f
C1136 net12 p[3] 0.00447f
C1137 _00_ _09_ 9.35e-21
C1138 p[3] _05_ 5.67e-20
C1139 _39_/a_47_47# _45_/a_193_297# 1.4e-20
C1140 _29_/a_29_53# _20_ 0.0111f
C1141 m1_7039_1799# b[3] 0.00448f
C1142 _15_ _47_/a_81_21# 0.00332f
C1143 net18 net10 3.35e-20
C1144 _19_ net1 2.86e-19
C1145 _22_ net15 2.74e-19
C1146 VGND _27_/a_109_297# -6.15e-19
C1147 _10_ _15_ 0.479f
C1148 _06_ p[14] 1.04e-19
C1149 _38_/a_27_47# _09_ 0.00195f
C1150 _44_/a_250_297# net3 0.0088f
C1151 b[3] output19/a_27_47# 0.00809f
C1152 VPWR _20_ 0.342f
C1153 _16_ _55_/a_80_21# 0.0143f
C1154 _06_ input4/a_75_212# 0.00205f
C1155 _50_/a_343_93# net14 1.07e-20
C1156 _04_ _13_ 1.17e-21
C1157 _36_/a_27_47# net10 0.0366f
C1158 _19_ net8 0.0322f
C1159 _11_ _17_ 0.197f
C1160 VGND p[10] 0.276f
C1161 _50_/a_223_47# _13_ 8.2e-20
C1162 net14 input5/a_558_47# 0.0325f
C1163 _17_ _37_/a_109_47# 8.86e-21
C1164 p[1] p[10] 8.79e-19
C1165 _25_ _12_ 1.23e-20
C1166 input7/a_27_47# net2 3.24e-19
C1167 _06_ net9 0.0505f
C1168 _04_ _09_ 0.0904f
C1169 VGND _53_/a_111_297# -2.89e-19
C1170 net5 _36_/a_197_47# 0.00254f
C1171 _15_ net14 0.225f
C1172 _06_ _50_/a_27_47# 0.00972f
C1173 net18 net11 0.00221f
C1174 net5 _39_/a_377_297# 0.00234f
C1175 _30_/a_109_53# _32_/a_27_47# 1.51e-19
C1176 _12_ _52_/a_346_47# 3.8e-19
C1177 net18 b[2] 0.0131f
C1178 _10_ _47_/a_299_297# 0.0134f
C1179 p[7] b[3] 0.0665f
C1180 _34_/a_377_297# _21_ 2.37e-19
C1181 _47_/a_81_21# _18_ 7.96e-20
C1182 _31_/a_285_297# _19_ 1.34e-19
C1183 VGND _41_/a_59_75# 0.0138f
C1184 _10_ _18_ 0.133f
C1185 VGND _33_/a_368_53# 2.38e-19
C1186 _53_/a_29_53# output18/a_27_47# 9.46e-19
C1187 _02_ output18/a_27_47# 4.13e-19
C1188 _01_ net11 3.82e-20
C1189 net13 _34_/a_285_47# 4.11e-20
C1190 VGND input10/a_27_47# 0.00285f
C1191 net5 _50_/a_343_93# 0.00124f
C1192 p[6] _02_ 3.73e-21
C1193 p[2] p[6] 0.03f
C1194 _36_/a_27_47# net11 0.0717f
C1195 VGND _30_/a_215_297# 0.016f
C1196 net11 _22_ 6.82e-21
C1197 _52_/a_256_47# _02_ 0.00344f
C1198 _34_/a_47_47# p[5] 7.86e-20
C1199 VGND _49_/a_208_47# -0.00164f
C1200 b[2] _22_ 0.00428f
C1201 net5 input5/a_558_47# 0.0597f
C1202 p[13] input5/a_664_47# 7.04e-19
C1203 _02_ _48_/a_181_47# 3.9e-19
C1204 _17_ _39_/a_129_47# 1.38e-20
C1205 _32_/a_27_47# net1 0.0211f
C1206 _10_ p[9] 0.00225f
C1207 _14_ _02_ 0.0316f
C1208 _48_/a_109_47# b[1] 4.46e-20
C1209 net1 _49_/a_201_297# 0.00304f
C1210 net5 _15_ 0.0352f
C1211 net2 input3/a_27_47# 0.0222f
C1212 _01_ _49_/a_544_297# 0.00109f
C1213 _06_ _53_/a_111_297# 3.82e-19
C1214 _53_/a_183_297# _09_ 4.18e-19
C1215 _30_/a_109_53# _20_ 8.12e-19
C1216 _27_/a_27_297# input5/a_664_47# 0.0116f
C1217 _17_ p[8] 0.00329f
C1218 net14 _18_ 0.0147f
C1219 _01_ net3 1.16e-19
C1220 _32_/a_27_47# _21_ 8.95e-19
C1221 _33_/a_109_93# _22_ 1.34e-22
C1222 input1/a_75_212# b[3] 1.21e-19
C1223 _42_/a_209_311# input3/a_27_47# 1.56e-19
C1224 VPWR _00_ 0.416f
C1225 _14_ _43_/a_27_47# 0.00938f
C1226 _32_/a_27_47# net8 0.0275f
C1227 _28_/a_109_297# net9 3.7e-19
C1228 _22_ net3 9.39e-20
C1229 _44_/a_584_47# net2 0.0053f
C1230 _44_/a_250_297# net19 0.00592f
C1231 _41_/a_59_75# _06_ 0.0429f
C1232 _06_ _33_/a_368_53# 1.7e-19
C1233 net8 _49_/a_201_297# 7.3e-19
C1234 VPWR _38_/a_27_47# -0.0142f
C1235 VGND _19_ 0.379f
C1236 VGND output16/a_27_47# 0.0728f
C1237 _19_ _43_/a_193_413# 4.85e-21
C1238 _37_/a_27_47# input6/a_27_47# 9.35e-19
C1239 p[9] net14 1.05e-19
C1240 _06_ _30_/a_215_297# 2.03e-20
C1241 _19_ p[1] 2.82e-20
C1242 _10_ _26_/a_29_53# 0.0265f
C1243 VGND _55_/a_217_297# -0.00342f
C1244 _45_/a_27_47# p[12] 6.12e-19
C1245 _55_/a_472_297# _02_ 1.25e-19
C1246 net1 _20_ 0.363f
C1247 net6 _47_/a_81_21# 2.14e-19
C1248 net5 _47_/a_299_297# 0.00198f
C1249 _29_/a_29_53# _04_ 0.0408f
C1250 _10_ net6 0.0965f
C1251 _11_ net9 5.39e-19
C1252 net3 input5/a_62_47# 0.00164f
C1253 _29_/a_29_53# _50_/a_223_47# 1.45e-20
C1254 _10_ b[1] 2.17e-19
C1255 _11_ _50_/a_27_47# 0.0592f
C1256 net5 _18_ 0.0426f
C1257 _39_/a_285_47# net6 1.53e-19
C1258 _44_/a_93_21# input5/a_558_47# 2.71e-19
C1259 VPWR _04_ 0.456f
C1260 _20_ _21_ 0.191f
C1261 VGND _34_/a_377_297# -9.51e-19
C1262 net8 _20_ 5.07e-19
C1263 VPWR _50_/a_223_47# -0.00601f
C1264 VGND _29_/a_183_297# 4.41e-19
C1265 _17_ _16_ 0.242f
C1266 _15_ _44_/a_93_21# 0.0168f
C1267 _26_/a_29_53# net14 1.33e-20
C1268 _35_/a_226_47# _49_/a_201_297# 1.66e-20
C1269 _14_ _55_/a_80_21# 0.0175f
C1270 _44_/a_250_297# output19/a_27_47# 6.42e-20
C1271 net12 p[7] 0.0351f
C1272 _35_/a_489_413# net10 0.00225f
C1273 _01_ _49_/a_315_47# 1.82e-19
C1274 input8/a_27_47# b[1] 2.46e-19
C1275 _34_/a_47_47# p[6] 0.00104f
C1276 net6 net14 2.82e-21
C1277 _27_/a_27_297# _17_ 6.78e-22
C1278 p[8] p[14] 0.0495f
C1279 _10_ _03_ 0.00244f
C1280 _06_ _55_/a_217_297# 3.46e-19
C1281 _36_/a_197_47# _25_ 2.37e-21
C1282 net17 net15 5.19e-19
C1283 VGND _50_/a_515_93# -4.75e-19
C1284 _30_/a_109_53# _00_ 3.67e-20
C1285 p[8] input4/a_75_212# 7.5e-20
C1286 _01_ net19 4.9e-19
C1287 VGND _32_/a_27_47# 0.0233f
C1288 _06_ _34_/a_377_297# 0.00427f
C1289 input15/a_27_47# _15_ 2.15e-20
C1290 VGND _49_/a_201_297# -0.00403f
C1291 net10 net17 8.67e-21
C1292 _41_/a_59_75# _11_ 8.7e-19
C1293 net5 _26_/a_29_53# 0.0237f
C1294 _22_ net19 2.17e-19
C1295 _35_/a_226_47# _20_ 5.19e-20
C1296 _50_/a_27_47# p[8] 3.39e-21
C1297 p[11] net3 0.00294f
C1298 _44_/a_93_21# _18_ 0.00485f
C1299 _45_/a_27_47# _35_/a_76_199# 2.04e-21
C1300 _03_ net14 1.5e-19
C1301 net5 net6 0.727f
C1302 net1 _00_ 9.43e-19
C1303 p[0] net7 1.36e-19
C1304 _38_/a_109_47# p[12] 8.9e-20
C1305 _10_ _08_ 1.51e-19
C1306 VPWR _41_/a_145_75# -2.46e-19
C1307 _12_ net4 0.105f
C1308 _02_ _47_/a_81_21# 1.59e-20
C1309 _30_/a_297_297# net9 7.83e-19
C1310 _30_/a_109_53# _04_ 9.19e-21
C1311 _30_/a_392_297# _03_ 6.33e-19
C1312 _35_/a_76_199# _07_ 0.00226f
C1313 _10_ _53_/a_29_53# 0.00779f
C1314 _10_ _02_ 0.0537f
C1315 _50_/a_515_93# _06_ 0.00244f
C1316 _00_ _21_ 9.26e-20
C1317 _39_/a_285_47# _02_ 0.0019f
C1318 _45_/a_193_297# _12_ 0.0103f
C1319 _40_/a_297_297# net15 4.08e-19
C1320 net8 _00_ 3.23e-19
C1321 VGND _20_ 0.471f
C1322 net17 input2/a_27_47# 0.0398f
C1323 _20_ _43_/a_193_413# 0.00161f
C1324 net11 net17 3.19e-20
C1325 _06_ _32_/a_27_47# 0.00663f
C1326 _38_/a_27_47# _21_ 3.87e-19
C1327 _10_ _43_/a_27_47# 0.0279f
C1328 input15/a_27_47# _18_ 8.27e-21
C1329 input2/a_27_47# net15 1.61e-19
C1330 net5 _03_ 1.04e-19
C1331 p[13] net9 1.72e-19
C1332 VPWR input7/a_27_47# 0.0768f
C1333 _04_ net1 0.018f
C1334 _43_/a_369_47# _18_ 1.49e-19
C1335 input8/a_27_47# _02_ 5.08e-20
C1336 input8/a_27_47# p[2] 0.0168f
C1337 _23_ _13_ 2.08e-20
C1338 _12_ _45_/a_465_47# 0.00211f
C1339 _02_ net14 0.00952f
C1340 output17/a_27_47# p[10] 0.124f
C1341 _17_ _43_/a_297_47# 5.72e-20
C1342 net2 net7 0.00234f
C1343 _31_/a_117_297# net7 0.00472f
C1344 _04_ _27_/a_277_297# 0.00113f
C1345 net9 _29_/a_111_297# 8.06e-21
C1346 p[13] _27_/a_109_297# 3.4e-20
C1347 _41_/a_59_75# p[8] 0.00214f
C1348 p[9] input15/a_27_47# 0.0195f
C1349 _23_ _09_ 0.207f
C1350 _04_ _21_ 0.39f
C1351 net10 input2/a_27_47# 1.17e-20
C1352 net10 net11 0.592f
C1353 net17 net3 3.72e-19
C1354 _04_ net8 0.02f
C1355 _50_/a_223_47# _21_ 2.91e-21
C1356 _45_/a_27_47# _13_ 0.0703f
C1357 net6 _44_/a_93_21# 1.08e-20
C1358 _43_/a_27_47# net14 4.87e-20
C1359 _55_/a_300_47# _15_ 1.42e-20
C1360 input13/a_27_47# net10 8.86e-20
C1361 net15 net3 0.394f
C1362 _52_/a_93_21# _04_ 2.35e-19
C1363 _06_ _20_ 0.133f
C1364 _27_/a_27_297# _27_/a_109_297# -3.68e-20
C1365 _35_/a_76_199# net7 1.79e-20
C1366 p[13] p[10] 0.21f
C1367 _07_ _13_ 3.22e-23
C1368 _45_/a_27_47# _09_ 0.00823f
C1369 VPWR _34_/a_129_47# -9.47e-19
C1370 p[11] net19 0.00635f
C1371 _30_/a_215_297# _30_/a_297_297# -8.88e-34
C1372 _17_ _14_ 0.489f
C1373 VPWR input3/a_27_47# 0.0687f
C1374 _33_/a_109_93# net10 0.0336f
C1375 net5 _02_ 0.233f
C1376 _10_ _55_/a_80_21# 5.49e-19
C1377 _12_ net12 7.94e-21
C1378 _12_ _05_ 2.52e-19
C1379 _07_ _09_ 0.0416f
C1380 _27_/a_27_297# p[10] 0.00116f
C1381 net16 _50_/a_27_47# 2.35e-20
C1382 input15/a_27_47# net6 0.146f
C1383 net11 b[2] 1.46e-19
C1384 _44_/a_584_47# VPWR -2.28e-19
C1385 VGND _00_ 0.139f
C1386 p[4] b[1] 0.0579f
C1387 net6 _43_/a_369_47# 3.62e-21
C1388 _00_ _43_/a_193_413# 0.00721f
C1389 _35_/a_226_47# _04_ 0.00551f
C1390 input6/a_27_47# _15_ 5.75e-19
C1391 net10 p[3] 9.6e-19
C1392 _11_ _32_/a_27_47# 1.65e-20
C1393 VPWR _50_/a_615_93# -5.34e-19
C1394 VGND _38_/a_27_47# 0.00766f
C1395 _40_/a_297_297# net3 2.54e-19
C1396 _55_/a_80_21# net14 4.7e-19
C1397 _10_ _36_/a_303_47# 4.09e-19
C1398 _25_ b[1] 0.00709f
C1399 _33_/a_109_93# net11 5.14e-19
C1400 VPWR _32_/a_109_47# 0.00124f
C1401 _33_/a_209_311# net12 0.0769f
C1402 _33_/a_209_311# _05_ 0.0311f
C1403 _31_/a_35_297# net2 0.0635f
C1404 _19_ output17/a_27_47# 7.69e-19
C1405 _25_ _54_/a_75_212# 0.0247f
C1406 _35_/a_76_199# net13 0.0337f
C1407 _28_/a_109_297# _20_ 0.00221f
C1408 input13/a_27_47# _33_/a_109_93# 0.00348f
C1409 b[0] _13_ 0.00305f
C1410 b[3] input5/a_558_47# 4.94e-19
C1411 net1 input7/a_27_47# 0.0383f
C1412 _10_ _50_/a_429_93# 0.00167f
C1413 _39_/a_377_297# net4 8.88e-19
C1414 _42_/a_109_93# net2 0.00507f
C1415 VGND _04_ 0.139f
C1416 _04_ _43_/a_193_413# 5.67e-21
C1417 p[5] input10/a_27_47# 0.0174f
C1418 _04_ p[1] 1.74e-21
C1419 net17 net19 8.84e-23
C1420 VGND _50_/a_223_47# 0.0159f
C1421 VPWR _23_ -0.00374f
C1422 net11 p[3] 3.1e-21
C1423 _06_ _00_ 0.1f
C1424 _09_ net7 0.00258f
C1425 p[14] _14_ 1.66e-20
C1426 _15_ b[3] 0.00381f
C1427 p[13] _19_ 8.22e-19
C1428 _11_ _20_ 0.268f
C1429 net19 net15 0.0501f
C1430 _39_/a_47_47# net15 9.44e-22
C1431 _25_ _03_ 0.00422f
C1432 _50_/a_343_93# net4 0.00124f
C1433 net5 _55_/a_80_21# 2.78e-19
C1434 input13/a_27_47# p[3] 0.00101f
C1435 input7/a_27_47# net8 2.03e-21
C1436 _06_ _38_/a_27_47# 0.0172f
C1437 _16_ _55_/a_217_297# 0.0017f
C1438 net17 input5/a_381_47# 1.37e-20
C1439 _29_/a_29_53# _07_ 1.19e-20
C1440 _45_/a_27_47# VPWR -0.00418f
C1441 _27_/a_27_297# _19_ 0.082f
C1442 _50_/a_429_93# net14 6.04e-21
C1443 _15_ net4 0.00427f
C1444 p[9] input6/a_27_47# 0.076f
C1445 _39_/a_47_47# net10 4.72e-22
C1446 _17_ _37_/a_197_47# 9.19e-21
C1447 net15 input5/a_381_47# 7.15e-19
C1448 net14 input5/a_664_47# 0.0179f
C1449 net18 _12_ 8.24e-19
C1450 VPWR _07_ 0.0728f
C1451 p[2] p[4] 5.33e-19
C1452 _06_ _04_ 0.0136f
C1453 _04_ _27_/a_205_297# 6.42e-19
C1454 VGND _53_/a_183_297# -4.34e-19
C1455 net5 _36_/a_303_47# 0.00256f
C1456 _06_ _50_/a_223_47# 0.0481f
C1457 net13 _13_ 4e-21
C1458 _10_ input9/a_75_212# 5.49e-21
C1459 _39_/a_129_47# _20_ 1.71e-20
C1460 _36_/a_27_47# _12_ 0.00178f
C1461 _12_ _22_ 0.196f
C1462 _25_ _53_/a_29_53# 0.00146f
C1463 _25_ _02_ 0.0156f
C1464 net15 output19/a_27_47# 6.88e-19
C1465 net13 _09_ 0.0379f
C1466 net16 output16/a_27_47# 0.0101f
C1467 _17_ _47_/a_81_21# 0.0456f
C1468 VGND _41_/a_145_75# 3.75e-19
C1469 _36_/a_197_47# net12 4.67e-20
C1470 _47_/a_299_297# net4 3.28e-19
C1471 input2/a_27_47# net19 2.9e-23
C1472 _10_ _17_ 0.0233f
C1473 _23_ _24_ 0.012f
C1474 p[8] _20_ 1.91e-20
C1475 _52_/a_346_47# _02_ 0.00526f
C1476 net5 input5/a_664_47# 0.0536f
C1477 p[9] b[3] 0.0985f
C1478 _17_ _39_/a_285_47# 7.36e-21
C1479 input6/a_27_47# net6 0.00208f
C1480 p[13] _32_/a_27_47# 6.49e-20
C1481 input8/a_27_47# input9/a_75_212# 3.09e-20
C1482 net4 _18_ 0.023f
C1483 p[6] input10/a_27_47# 0.00448f
C1484 _29_/a_29_53# net7 6.01e-19
C1485 _11_ _00_ 0.238f
C1486 _06_ _53_/a_183_297# 0.00146f
C1487 _45_/a_27_47# _24_ 4.57e-19
C1488 VGND input7/a_27_47# 0.0574f
C1489 VPWR b[0] 0.226f
C1490 _12_ _45_/a_205_47# 7.46e-19
C1491 input7/a_27_47# p[1] 0.0169f
C1492 _32_/a_109_47# net8 0.0011f
C1493 _11_ _38_/a_27_47# 0.071f
C1494 VPWR net7 0.784f
C1495 _17_ net14 0.104f
C1496 net19 net3 0.611f
C1497 _39_/a_47_47# net3 1.66e-20
C1498 _24_ _07_ 5.67e-19
C1499 input14/a_27_47# net2 0.0176f
C1500 VPWR _38_/a_109_47# -4.66e-19
C1501 net10 p[7] 5.59e-19
C1502 _10_ _26_/a_111_297# 7.13e-20
C1503 b[3] net6 7.68e-19
C1504 _55_/a_300_47# _02_ 0.00371f
C1505 _23_ _21_ 0.0217f
C1506 b[1] b[3] 1.94f
C1507 _16_ _20_ 0.00271f
C1508 net3 input5/a_381_47# 0.0299f
C1509 output16/a_27_47# output18/a_27_47# 7.85e-19
C1510 _54_/a_75_212# b[3] 0.0013f
C1511 input5/a_841_47# VPWR 0.0775f
C1512 _11_ _50_/a_223_47# 0.0329f
C1513 _39_/a_129_47# _00_ 1.63e-20
C1514 _26_/a_29_53# net4 0.00412f
C1515 _52_/a_93_21# _23_ 0.0166f
C1516 _44_/a_93_21# input5/a_664_47# 1.88e-20
C1517 _10_ p[14] 1.53e-19
C1518 VGND _34_/a_129_47# -8.76e-20
C1519 _27_/a_27_297# _20_ 3.14e-20
C1520 _07_ net1 6.08e-22
C1521 _44_/a_250_297# _15_ 0.00517f
C1522 net5 _17_ 0.00408f
C1523 VGND input3/a_27_47# 0.0414f
C1524 net6 net4 0.713f
C1525 _45_/a_27_47# _21_ 1.18e-20
C1526 _29_/a_29_53# net13 0.00104f
C1527 b[1] net4 9.59e-20
C1528 _10_ input4/a_75_212# 0.00372f
C1529 _19_ _14_ 2.71e-21
C1530 p[8] _00_ 8.85e-20
C1531 _25_ _34_/a_47_47# 1.08e-19
C1532 _01_ _49_/a_75_199# 0.009f
C1533 _14_ _55_/a_217_297# 0.0116f
C1534 output19/a_27_47# net3 0.00348f
C1535 net11 p[7] 3.28e-20
C1536 _35_/a_226_297# net10 2.48e-19
C1537 net12 _18_ 2.25e-21
C1538 _07_ _21_ 0.133f
C1539 _03_ b[3] 3.79e-21
C1540 _45_/a_193_297# net6 9.84e-20
C1541 _52_/a_93_21# _45_/a_27_47# 1.18e-19
C1542 net9 _47_/a_81_21# 3.49e-19
C1543 VPWR net13 0.599f
C1544 _34_/a_377_297# p[6] 5.88e-19
C1545 VGND _44_/a_584_47# -0.00145f
C1546 _22_ _49_/a_75_199# 9.85e-21
C1547 input13/a_27_47# p[7] 0.0157f
C1548 _10_ net9 0.0438f
C1549 _36_/a_303_47# _25_ 2.03e-21
C1550 VPWR input11/a_27_47# 0.0375f
C1551 _10_ _50_/a_27_47# 0.0154f
C1552 VGND _50_/a_615_93# -5.19e-19
C1553 p[14] net14 6.11e-20
C1554 _23_ _35_/a_226_47# 4.21e-19
C1555 _44_/a_346_47# net2 1.64e-19
C1556 _31_/a_35_297# VPWR 0.0333f
C1557 VGND _32_/a_109_47# 1.05e-19
C1558 _45_/a_465_47# net6 6.06e-20
C1559 _06_ _34_/a_129_47# 5.3e-19
C1560 input8/a_27_47# net9 3.71e-20
C1561 VPWR _42_/a_109_93# -0.00118f
C1562 _45_/a_193_297# _03_ 2.57e-20
C1563 _08_ b[3] 2.22e-20
C1564 _45_/a_27_47# _35_/a_226_47# 5.71e-21
C1565 net9 net14 7.12e-20
C1566 _37_/a_27_47# net15 0.0541f
C1567 _01_ _50_/a_343_93# 0.0131f
C1568 net1 net7 0.0712f
C1569 _38_/a_197_47# p[12] 1.05e-19
C1570 _17_ _44_/a_93_21# 0.0646f
C1571 _01_ input5/a_558_47# 3.97e-20
C1572 b[3] _02_ 2.33e-19
C1573 p[2] b[3] 0.047f
C1574 _16_ _00_ 0.00613f
C1575 p[7] p[3] 0.0664f
C1576 VGND _23_ 0.16f
C1577 _50_/a_343_93# _22_ 0.0597f
C1578 _40_/a_191_297# net6 1.16e-20
C1579 _30_/a_465_297# _03_ 7.72e-19
C1580 _30_/a_392_297# net9 9.92e-19
C1581 _35_/a_226_47# _07_ 8.96e-19
C1582 _04_ output17/a_27_47# 0.027f
C1583 _27_/a_109_297# net14 1.32e-19
C1584 net12 _26_/a_29_53# 6.55e-19
C1585 _10_ _53_/a_111_297# 2.06e-19
C1586 net19 input5/a_381_47# 0.00173f
C1587 _50_/a_615_93# _06_ 0.00264f
C1588 _01_ _15_ 0.007f
C1589 _21_ net7 3e-19
C1590 _33_/a_209_311# _35_/a_489_413# 2.77e-20
C1591 net12 net6 0.00643f
C1592 net5 input4/a_75_212# 0.0104f
C1593 net8 net7 0.295f
C1594 _41_/a_59_75# _47_/a_81_21# 1.5e-19
C1595 _12_ net15 8.14e-21
C1596 _14_ _49_/a_201_297# 4.76e-21
C1597 net12 b[1] 0.00225f
C1598 b[1] _05_ 5.56e-20
C1599 _10_ _41_/a_59_75# 0.0172f
C1600 _15_ _22_ 0.0236f
C1601 VGND _45_/a_27_47# -0.029f
C1602 net13 _30_/a_109_53# 1.05e-19
C1603 _02_ net4 0.00376f
C1604 _53_/a_29_53# net4 3.26e-19
C1605 input5/a_841_47# net1 1.33e-19
C1606 p[10] net14 3.33e-19
C1607 _45_/a_109_297# p[12] 1.52e-21
C1608 net5 net9 0.0368f
C1609 p[13] _04_ 0.00155f
C1610 _10_ _30_/a_215_297# 5.66e-20
C1611 _43_/a_469_47# _18_ 1.59e-19
C1612 net19 output19/a_27_47# 0.0279f
C1613 _17_ input15/a_27_47# 6.14e-19
C1614 net5 _50_/a_27_47# 0.0169f
C1615 VGND _07_ 0.195f
C1616 _45_/a_193_297# _02_ 0.00988f
C1617 _12_ net10 7.82e-20
C1618 _17_ _43_/a_369_47# 5.87e-19
C1619 input5/a_841_47# _21_ 1.59e-21
C1620 _31_/a_285_297# net7 0.00227f
C1621 _04_ _29_/a_111_297# 9.25e-19
C1622 _31_/a_35_297# _30_/a_109_53# 2.89e-20
C1623 _33_/a_209_311# net17 7.03e-21
C1624 input5/a_841_47# net8 0.025f
C1625 _23_ _06_ 0.218f
C1626 _27_/a_27_297# _04_ 0.0526f
C1627 VPWR input12/a_27_47# 0.0646f
C1628 _03_ net12 0.0268f
C1629 net13 net1 3.51e-19
C1630 _03_ _05_ 0.135f
C1631 _20_ _14_ 0.144f
C1632 _01_ _18_ 6.1e-20
C1633 net16 _38_/a_27_47# 0.114f
C1634 _52_/a_250_297# _04_ 3.98e-21
C1635 _35_/a_226_47# net7 2.93e-20
C1636 _36_/a_27_47# _18_ 5.46e-20
C1637 net5 p[10] 5.12e-21
C1638 p[14] _44_/a_93_21# 2.82e-20
C1639 _22_ _18_ 0.0211f
C1640 _45_/a_27_47# _06_ 0.0021f
C1641 net13 _21_ 0.13f
C1642 b[3] _55_/a_80_21# 3.94e-19
C1643 VPWR _34_/a_285_47# -0.00233f
C1644 _31_/a_35_297# net1 0.0111f
C1645 net13 net8 7.51e-20
C1646 _33_/a_209_311# net10 0.0426f
C1647 _10_ _55_/a_217_297# 1.43e-19
C1648 _12_ net11 0.00799f
C1649 _12_ b[2] 3.89e-20
C1650 _06_ _07_ 0.185f
C1651 _52_/a_93_21# net13 7.21e-19
C1652 _37_/a_27_47# net3 0.0887f
C1653 net12 _08_ 0.0269f
C1654 _08_ _05_ 0.00897f
C1655 net16 _50_/a_223_47# 4.77e-21
C1656 _55_/a_472_297# _20_ 0.00212f
C1657 VGND b[0] 0.217f
C1658 net5 _41_/a_59_75# 2.41e-19
C1659 _31_/a_35_297# net8 0.0408f
C1660 _55_/a_80_21# net4 1.06e-19
C1661 VGND net7 0.419f
C1662 net6 _43_/a_469_47# 4.85e-21
C1663 _00_ _43_/a_297_47# 1.26e-19
C1664 _48_/a_27_47# _07_ 0.0524f
C1665 _43_/a_193_413# net7 3.49e-19
C1666 p[1] net7 0.00706f
C1667 _31_/a_285_297# net13 3.85e-20
C1668 VPWR input14/a_27_47# 0.0735f
C1669 net12 _02_ 2.28e-19
C1670 input15/a_27_47# p[14] 6.15e-19
C1671 net18 _26_/a_29_53# 2.57e-21
C1672 _05_ _02_ 0.00163f
C1673 net5 _30_/a_215_297# 8.27e-21
C1674 p[2] _05_ 3.69e-19
C1675 _33_/a_109_93# _12_ 9.75e-20
C1676 _10_ _29_/a_183_297# 6.24e-20
C1677 _19_ net14 0.0512f
C1678 VGND _38_/a_109_47# 2.3e-19
C1679 net17 _49_/a_75_199# 0.00127f
C1680 _12_ net3 3.09e-20
C1681 p[11] _15_ 2.63e-19
C1682 _55_/a_217_297# net14 2.1e-19
C1683 input15/a_27_47# input4/a_75_212# 1.1e-21
C1684 net18 b[1] 0.00569f
C1685 _52_/a_584_47# _26_/a_29_53# 7.45e-20
C1686 _33_/a_209_311# net11 2.49e-19
C1687 VPWR _32_/a_197_47# 0.00146f
C1688 _33_/a_296_53# net12 1.23e-20
C1689 _33_/a_296_53# _05_ 4.53e-19
C1690 _49_/a_75_199# net15 5.13e-20
C1691 net18 _54_/a_75_212# 0.0143f
C1692 _36_/a_27_47# _26_/a_29_53# 1.6e-19
C1693 _35_/a_226_47# net13 0.00709f
C1694 _38_/a_27_47# output18/a_27_47# 8.6e-19
C1695 input13/a_27_47# _33_/a_209_311# 5.85e-20
C1696 _22_ _26_/a_29_53# 0.09f
C1697 input5/a_841_47# VGND 0.0942f
C1698 p[8] input3/a_27_47# 6.2e-19
C1699 _36_/a_27_47# net6 5.1e-19
C1700 _23_ _11_ 2e-20
C1701 _10_ _50_/a_515_93# 0.00129f
C1702 b[3] input5/a_664_47# 4.72e-19
C1703 _42_/a_209_311# net2 5.1e-19
C1704 _22_ net6 0.163f
C1705 _14_ _00_ 0.133f
C1706 _32_/a_27_47# _47_/a_81_21# 5.06e-21
C1707 b[1] _22_ 1.02e-19
C1708 VPWR _44_/a_256_47# -7.56e-19
C1709 _10_ _32_/a_27_47# 0.00217f
C1710 _06_ net7 0.00447f
C1711 net5 _19_ 6.41e-21
C1712 _44_/a_584_47# p[8] 1.27e-19
C1713 net5 output16/a_27_47# 4.14e-19
C1714 net18 _03_ 2.07e-21
C1715 _27_/a_27_297# input7/a_27_47# 0.00119f
C1716 output17/a_27_47# input3/a_27_47# 3.15e-19
C1717 _50_/a_429_93# net4 4.16e-19
C1718 net5 _55_/a_217_297# 8.84e-20
C1719 net1 input12/a_27_47# 7.44e-20
C1720 _13_ p[12] 0.00395f
C1721 _45_/a_27_47# _11_ 0.0703f
C1722 VGND net13 0.145f
C1723 _50_/a_615_93# p[8] 5.93e-20
C1724 _17_ input6/a_27_47# 7.13e-22
C1725 _01_ _03_ 2.85e-19
C1726 net17 input5/a_558_47# 2.88e-21
C1727 _09_ p[12] 0.00189f
C1728 _50_/a_515_93# net14 1.39e-20
C1729 VGND input11/a_27_47# 0.0274f
C1730 input12/a_27_47# _21_ 2.32e-19
C1731 _44_/a_346_47# VPWR -8.74e-19
C1732 _03_ _22_ 2.55e-20
C1733 _04_ _14_ 2.04e-21
C1734 net6 _45_/a_205_47# 2.59e-20
C1735 _37_/a_27_47# net19 0.0105f
C1736 _17_ _37_/a_303_47# 1.23e-20
C1737 input5/a_841_47# _06_ 1.66e-19
C1738 net15 input5/a_558_47# 0.00672f
C1739 input8/a_27_47# _49_/a_201_297# 2.46e-21
C1740 p[13] input3/a_27_47# 0.00499f
C1741 VGND _31_/a_35_297# -0.00829f
C1742 p[9] p[11] 0.0303f
C1743 _20_ _47_/a_81_21# 0.0457f
C1744 net11 _49_/a_75_199# 4.49e-19
C1745 input9/a_75_212# b[3] 1.21e-19
C1746 _49_/a_201_297# net14 1.52e-19
C1747 _10_ _20_ 0.179f
C1748 _15_ net15 0.156f
C1749 VGND _42_/a_109_93# -0.0045f
C1750 _34_/a_285_47# _21_ 6.94e-20
C1751 _41_/a_59_75# input15/a_27_47# 3.96e-20
C1752 _34_/a_47_47# net12 0.0385f
C1753 _34_/a_47_47# _05_ 1.26e-20
C1754 _39_/a_47_47# _12_ 0.0317f
C1755 net18 _53_/a_29_53# 0.0118f
C1756 net18 _02_ 8.53e-20
C1757 p[4] input10/a_27_47# 0.0217f
C1758 _17_ b[3] 0.00637f
C1759 _06_ net13 0.0766f
C1760 _36_/a_303_47# net12 1.37e-19
C1761 _52_/a_584_47# _02_ 0.00389f
C1762 _01_ _02_ 0.106f
C1763 p[2] _01_ 0.00164f
C1764 net5 _32_/a_27_47# 0.0961f
C1765 VPWR _26_/a_183_297# -3.03e-19
C1766 _49_/a_75_199# net3 2.01e-19
C1767 _25_ input10/a_27_47# 2.03e-20
C1768 _32_/a_197_47# net1 0.00142f
C1769 _36_/a_27_47# _02_ 9.37e-20
C1770 _20_ net14 8.01e-20
C1771 _22_ _02_ 0.552f
C1772 _53_/a_29_53# _22_ 0.00749f
C1773 net15 _47_/a_299_297# 1.44e-20
C1774 _17_ net4 7.52e-21
C1775 input6/a_27_47# p[14] 0.0155f
C1776 _01_ _43_/a_27_47# 9.77e-20
C1777 b[1] p[11] 1.84e-20
C1778 _35_/a_76_199# _13_ 3.01e-21
C1779 input2/a_27_47# input5/a_558_47# 2.04e-20
C1780 net15 _18_ 0.0382f
C1781 _42_/a_109_93# _06_ 5.53e-20
C1782 _32_/a_197_47# net8 3.39e-20
C1783 _22_ _43_/a_27_47# 0.091f
C1784 input2/a_27_47# _15_ 3.18e-20
C1785 _35_/a_76_199# _09_ 0.047f
C1786 VPWR _38_/a_197_47# -5.24e-19
C1787 p[9] net15 0.00306f
C1788 VGND input12/a_27_47# 0.0405f
C1789 net10 _18_ 1.47e-21
C1790 net5 _20_ 0.0651f
C1791 _00_ _47_/a_81_21# 0.0258f
C1792 VPWR p[12] 0.0895f
C1793 _40_/a_109_297# net2 0.0011f
C1794 _10_ _00_ 0.301f
C1795 net3 input5/a_558_47# 0.0137f
C1796 b[0] _39_/a_129_47# 2.6e-20
C1797 p[14] b[3] 0.0673f
C1798 VPWR p[0] 0.0906f
C1799 _39_/a_285_47# _00_ 1.47e-21
C1800 _52_/a_250_297# _23_ 3.17e-19
C1801 _10_ _38_/a_27_47# 0.0133f
C1802 VGND _34_/a_285_47# -0.00301f
C1803 _15_ net3 0.224f
C1804 VPWR _45_/a_109_297# -0.011f
C1805 _01_ _55_/a_80_21# 0.0121f
C1806 input9/a_75_212# _05_ 1.24e-21
C1807 _17_ _40_/a_191_297# 4.35e-19
C1808 _26_/a_29_53# net15 9.06e-21
C1809 _22_ _55_/a_80_21# 0.00926f
C1810 net17 b[1] 0.00731f
C1811 _35_/a_489_413# _03_ 0.0205f
C1812 _35_/a_556_47# net10 5.59e-19
C1813 _47_/a_384_47# _12_ 9.51e-20
C1814 net9 b[3] 2.37e-20
C1815 net6 net15 0.0664f
C1816 _00_ net14 4.11e-20
C1817 _34_/a_129_47# p[6] 2.01e-20
C1818 _06_ input12/a_27_47# 5.3e-22
C1819 _10_ _04_ 9.24e-20
C1820 VGND input14/a_27_47# 0.0389f
C1821 net4 input4/a_75_212# 0.0189f
C1822 _10_ _50_/a_223_47# 0.0295f
C1823 b[3] _27_/a_109_297# 5.52e-20
C1824 _13_ _09_ 0.0927f
C1825 output17/a_27_47# net7 0.00185f
C1826 net10 _26_/a_29_53# 3.48e-22
C1827 _34_/a_47_47# _22_ 3.9e-21
C1828 VPWR net2 0.918f
C1829 _47_/a_299_297# net3 2.55e-19
C1830 _31_/a_117_297# VPWR 8.41e-19
C1831 _45_/a_27_47# net16 8.68e-19
C1832 VGND _32_/a_197_47# 8.12e-20
C1833 _33_/a_209_311# p[7] 3.7e-19
C1834 _35_/a_226_297# _12_ 3.35e-20
C1835 net9 net4 1.99e-22
C1836 net10 net6 1.35e-20
C1837 _06_ _34_/a_285_47# 0.00598f
C1838 _50_/a_27_47# net4 0.0239f
C1839 net10 b[1] 0.00244f
C1840 _03_ net17 5.1e-19
C1841 net3 _18_ 7.34e-20
C1842 _29_/a_29_53# _35_/a_76_199# 9.88e-19
C1843 input8/a_27_47# _04_ 2.36e-22
C1844 VPWR _42_/a_209_311# -0.00753f
C1845 _35_/a_489_413# _08_ 5.56e-19
C1846 p[10] b[3] 0.12f
C1847 net10 _54_/a_75_212# 7.43e-19
C1848 _44_/a_250_297# _17_ 0.0336f
C1849 _03_ net15 4.26e-20
C1850 _04_ net14 0.0863f
C1851 net5 _00_ 0.00954f
C1852 p[13] net7 1.91e-19
C1853 _48_/a_27_47# _34_/a_285_47# 6.66e-20
C1854 VPWR _35_/a_76_199# -0.00947f
C1855 _38_/a_303_47# p[12] 9.56e-20
C1856 _50_/a_223_47# net14 5.89e-21
C1857 _35_/a_489_413# _02_ 3.86e-19
C1858 VGND _44_/a_256_47# -0.00184f
C1859 _16_ net7 7.5e-20
C1860 _40_/a_297_297# net6 7.47e-22
C1861 _30_/a_465_297# net9 0.00138f
C1862 p[9] net3 1.63e-19
C1863 net5 _38_/a_27_47# 1.76e-19
C1864 net11 _26_/a_29_53# 1.08e-20
C1865 _10_ _53_/a_183_297# 2.86e-19
C1866 net19 input5/a_558_47# 2.24e-20
C1867 _27_/a_27_297# net7 1.22e-19
C1868 net10 _03_ 0.321f
C1869 net11 net6 1.08e-19
C1870 b[3] input10/a_27_47# 1.21e-19
C1871 b[1] input2/a_27_47# 4.12e-19
C1872 net11 b[1] 0.0128f
C1873 _15_ net19 0.166f
C1874 b[2] b[1] 0.126f
C1875 input5/a_841_47# p[13] 1.2e-19
C1876 _30_/a_215_297# b[3] 2.74e-20
C1877 net13 _30_/a_297_297# 3.27e-20
C1878 _53_/a_111_297# net4 2.09e-19
C1879 net11 _54_/a_75_212# 0.00956f
C1880 input13/a_27_47# b[1] 2.46e-19
C1881 p[0] net1 0.00473f
C1882 _10_ _41_/a_145_75# 5.18e-19
C1883 _23_ _52_/a_256_47# 6.66e-19
C1884 VGND _44_/a_346_47# -0.00198f
C1885 net5 _04_ 0.00476f
C1886 input5/a_841_47# _16_ 8.62e-19
C1887 net17 _02_ 0.0608f
C1888 net5 _50_/a_223_47# 0.00202f
C1889 _41_/a_59_75# net4 1.76e-19
C1890 _26_/a_29_53# net3 2.83e-21
C1891 _02_ net15 0.0806f
C1892 _17_ _43_/a_469_47# 0.00177f
C1893 _31_/a_285_47# net7 0.00132f
C1894 net16 b[0] 0.0322f
C1895 _33_/a_109_93# b[1] 2.53e-20
C1896 net6 net3 0.00152f
C1897 _03_ input2/a_27_47# 2.71e-19
C1898 b[1] net3 1.6e-20
C1899 _03_ net11 0.0952f
C1900 net9 net12 0.0596f
C1901 net10 _08_ 0.194f
C1902 net9 _05_ 0.124f
C1903 _00_ _44_/a_93_21# 4.54e-20
C1904 _07_ p[6] 1.38e-19
C1905 _50_/a_27_47# net12 7.99e-21
C1906 _42_/a_109_93# output17/a_27_47# 8.6e-21
C1907 net16 _38_/a_109_47# 4.17e-19
C1908 VPWR _13_ 0.0804f
C1909 _29_/a_29_53# _09_ 0.00488f
C1910 net10 _53_/a_29_53# 7.88e-22
C1911 net10 _02_ 6.74e-19
C1912 _07_ _48_/a_181_47# 5.93e-19
C1913 _19_ b[3] 0.00431f
C1914 _01_ _17_ 1.46e-20
C1915 _39_/a_47_47# _18_ 1.23e-19
C1916 net19 _18_ 4.89e-20
C1917 b[3] _55_/a_217_297# 3.41e-19
C1918 p[3] b[1] 0.0494f
C1919 VGND _26_/a_183_297# 2.42e-19
C1920 net1 net2 1.64e-19
C1921 VPWR _09_ 0.297f
C1922 _17_ _22_ 0.00334f
C1923 _33_/a_109_93# _03_ 2.78e-19
C1924 _33_/a_296_53# net10 8.22e-20
C1925 _03_ _49_/a_544_297# 0.00568f
C1926 input8/a_27_47# input7/a_27_47# 3.2e-20
C1927 _03_ net3 4.27e-20
C1928 p[9] net19 0.0727f
C1929 p[10] _05_ 6e-20
C1930 _11_ input14/a_27_47# 1.42e-19
C1931 net13 p[5] 1.05e-19
C1932 net11 _08_ 8.83e-19
C1933 input7/a_27_47# net14 3.48e-19
C1934 output16/a_27_47# net4 0.00706f
C1935 _04_ _44_/a_93_21# 4.47e-21
C1936 net2 net8 0.0525f
C1937 _31_/a_117_297# net8 5.91e-19
C1938 _55_/a_217_297# net4 1.13e-19
C1939 net11 _53_/a_29_53# 8.31e-19
C1940 net11 _02_ 0.0327f
C1941 input11/a_27_47# p[5] 0.0491f
C1942 _53_/a_29_53# b[2] 6.22e-19
C1943 b[2] _02_ 2.81e-19
C1944 _27_/a_27_297# _42_/a_109_93# 1.35e-20
C1945 _33_/a_209_311# _12_ 2.88e-20
C1946 _03_ p[3] 0.00359f
C1947 VGND _38_/a_197_47# 2.29e-19
C1948 _42_/a_209_311# net8 7.7e-21
C1949 _35_/a_226_47# _45_/a_109_297# 1.59e-21
C1950 p[2] input13/a_27_47# 3.58e-19
C1951 _55_/a_80_21# net15 0.00759f
C1952 _35_/a_76_199# _21_ 0.0175f
C1953 VPWR _40_/a_109_297# -4.23e-19
C1954 VPWR _32_/a_303_47# 6.03e-19
C1955 _33_/a_368_53# net12 2.63e-19
C1956 _33_/a_368_53# _05_ 9.2e-19
C1957 _47_/a_384_47# _15_ 0.00112f
C1958 _06_ _26_/a_183_297# 3.16e-19
C1959 VGND p[12] 0.649f
C1960 net12 input10/a_27_47# 0.00115f
C1961 _25_ _38_/a_27_47# 5.76e-19
C1962 _10_ _44_/a_584_47# 1.14e-20
C1963 _30_/a_215_297# net12 0.00676f
C1964 _22_ _26_/a_111_297# 0.00137f
C1965 _24_ _13_ 2.47e-19
C1966 _30_/a_215_297# _05_ 0.0453f
C1967 _52_/a_93_21# _35_/a_76_199# 6.83e-21
C1968 _33_/a_109_93# _02_ 1.54e-21
C1969 VGND p[0] 0.135f
C1970 p[0] p[1] 0.062f
C1971 _10_ _50_/a_615_93# 8.82e-19
C1972 _14_ net7 0.00251f
C1973 net19 net6 0.00352f
C1974 _39_/a_47_47# net6 0.0249f
C1975 _02_ net3 9.52e-20
C1976 input3/a_27_47# net14 3.47e-19
C1977 p[9] output19/a_27_47# 0.0847f
C1978 _24_ _09_ 0.0202f
C1979 VGND _45_/a_109_297# -0.00179f
C1980 _03_ _49_/a_315_47# 9.22e-19
C1981 p[8] input14/a_27_47# 0.0169f
C1982 _06_ _38_/a_197_47# 4.32e-19
C1983 p[2] p[3] 0.124f
C1984 _44_/a_584_47# net14 7.2e-19
C1985 _07_ _48_/a_109_47# 3.01e-19
C1986 _29_/a_29_53# VPWR 0.0299f
C1987 _34_/a_47_47# net10 0.0507f
C1988 _01_ net9 0.157f
C1989 _06_ p[12] 0.0567f
C1990 _50_/a_615_93# net14 1.69e-20
C1991 _35_/a_76_199# _35_/a_226_47# -2.84e-32
C1992 _36_/a_27_47# net9 0.00493f
C1993 _10_ _23_ 0.00192f
C1994 _39_/a_47_47# _03_ 1.47e-19
C1995 net9 _22_ 0.0023f
C1996 net15 input5/a_664_47# 0.0216f
C1997 _23_ _39_/a_285_47# 1.9e-20
C1998 _36_/a_27_47# _50_/a_27_47# 6.08e-19
C1999 net1 _09_ 5.26e-20
C2000 VGND net2 0.831f
C2001 VGND _31_/a_117_297# -0.00177f
C2002 net2 _43_/a_193_413# 1.52e-19
C2003 _50_/a_27_47# _22_ 0.0276f
C2004 b[3] _20_ 1.58e-19
C2005 p[1] net2 5.99e-20
C2006 _13_ _21_ 1.69e-19
C2007 net6 output19/a_27_47# 0.00112f
C2008 _06_ _45_/a_109_297# 0.0023f
C2009 VGND _42_/a_209_311# -0.008f
C2010 input12/a_27_47# p[5] 0.00362f
C2011 p[6] input11/a_27_47# 4.64e-20
C2012 p[8] _44_/a_256_47# 6.54e-20
C2013 _10_ _45_/a_27_47# 0.0143f
C2014 _52_/a_93_21# _13_ 1.31e-19
C2015 _21_ _09_ 0.263f
C2016 _34_/a_377_297# net12 0.00251f
C2017 _34_/a_47_47# net11 0.0309f
C2018 net9 input5/a_62_47# 3.12e-19
C2019 _49_/a_315_47# _02_ 0.00134f
C2020 p[2] _49_/a_315_47# 6.65e-20
C2021 _39_/a_377_297# _12_ 6.77e-19
C2022 _01_ p[10] 1.64e-19
C2023 VGND _35_/a_76_199# -0.0034f
C2024 p[13] input14/a_27_47# 1.37e-19
C2025 _20_ net4 3.01e-20
C2026 _10_ _07_ 2.19e-19
C2027 _52_/a_93_21# _09_ 0.0227f
C2028 _55_/a_80_21# net3 2.35e-19
C2029 _36_/a_303_47# net11 7.63e-20
C2030 _37_/a_27_47# _15_ 1.11e-19
C2031 net5 _32_/a_109_47# 5.69e-21
C2032 _50_/a_343_93# _12_ 5.63e-20
C2033 net18 input10/a_27_47# 4.16e-20
C2034 _32_/a_303_47# net1 1.45e-19
C2035 _44_/a_346_47# p[8] 7.21e-20
C2036 net19 _02_ 0.0474f
C2037 _39_/a_47_47# _02_ 0.0127f
C2038 _53_/a_111_297# _22_ 4.7e-20
C2039 _06_ net2 0.0108f
C2040 p[7] b[1] 0.0436f
C2041 _42_/a_109_93# _14_ 0.00141f
C2042 _29_/a_29_53# _30_/a_109_53# 0.0103f
C2043 _35_/a_226_47# _13_ 5.62e-21
C2044 input2/a_27_47# input5/a_664_47# 4.47e-21
C2045 _12_ _15_ 0.00833f
C2046 _41_/a_59_75# _22_ 6.24e-22
C2047 _42_/a_209_311# _06_ 1.66e-19
C2048 VPWR _24_ 0.0129f
C2049 _32_/a_27_47# net12 1.52e-19
C2050 _01_ _49_/a_208_47# 2.13e-19
C2051 _32_/a_303_47# net8 2.22e-34
C2052 _32_/a_27_47# _05_ 2.2e-20
C2053 VPWR _30_/a_109_53# 0.0012f
C2054 _17_ net15 0.195f
C2055 net5 _23_ 0.0052f
C2056 _36_/a_27_47# _30_/a_215_297# 7.13e-20
C2057 _30_/a_215_297# _22_ 2.46e-21
C2058 _35_/a_76_199# _06_ 0.00425f
C2059 net10 input9/a_75_212# 0.00699f
C2060 _35_/a_226_47# _09_ 0.0599f
C2061 VPWR _38_/a_303_47# -4.83e-19
C2062 _11_ p[12] 3.93e-19
C2063 _37_/a_27_47# _18_ 3.31e-20
C2064 _29_/a_29_53# net1 9.76e-19
C2065 b[3] _00_ 1.04e-19
C2066 VGND _13_ 0.363f
C2067 net5 _45_/a_27_47# 0.0288f
C2068 _13_ _43_/a_193_413# 5.58e-21
C2069 _10_ net7 6.22e-20
C2070 input1/a_75_212# b[1] 0.00382f
C2071 _40_/a_191_297# _20_ 2.07e-20
C2072 net3 input5/a_664_47# 0.00215f
C2073 b[0] _39_/a_285_47# 1.88e-19
C2074 VPWR net1 1.17f
C2075 _11_ _45_/a_109_297# 0.00168f
C2076 _12_ _47_/a_299_297# 0.00805f
C2077 _29_/a_29_53# _21_ 0.0775f
C2078 input12/a_27_47# p[6] 0.0188f
C2079 _10_ _38_/a_109_47# 5.44e-19
C2080 p[9] _37_/a_27_47# 0.0117f
C2081 VGND _09_ 0.396f
C2082 _01_ _19_ 0.031f
C2083 net12 _20_ 0.00437f
C2084 _05_ _20_ 6.79e-19
C2085 VPWR _27_/a_277_297# -3.63e-19
C2086 _12_ _18_ 0.0115f
C2087 _00_ net4 0.0166f
C2088 _01_ _55_/a_217_297# 0.00112f
C2089 net11 input9/a_75_212# 1.1e-20
C2090 VPWR _21_ 0.871f
C2091 input13/a_27_47# input9/a_75_212# 0.00732f
C2092 input8/a_27_47# net7 1.47e-19
C2093 VPWR net8 0.703f
C2094 net19 _55_/a_80_21# 0.00423f
C2095 _08_ p[7] 0.00201f
C2096 _39_/a_129_47# p[12] 2.2e-20
C2097 _38_/a_27_47# net4 0.0119f
C2098 _35_/a_226_297# _03_ 0.00101f
C2099 _04_ b[3] 0.00415f
C2100 _45_/a_193_297# _00_ 4.38e-20
C2101 _34_/a_285_47# p[6] 2.23e-19
C2102 net14 net7 2.23e-19
C2103 p[11] p[10] 0.00297f
C2104 _52_/a_93_21# VPWR -0.00838f
C2105 p[2] p[7] 0.0856f
C2106 _11_ net2 0.234f
C2107 _06_ _13_ 0.00188f
C2108 p[14] net15 0.00132f
C2109 p[8] p[12] 0.804f
C2110 _19_ input5/a_62_47# 0.00159f
C2111 _31_/a_285_297# VPWR 0.0174f
C2112 VGND _40_/a_109_297# -0.00181f
C2113 VGND _32_/a_303_47# -4.83e-19
C2114 _37_/a_27_47# net6 4.3e-20
C2115 _06_ _09_ 0.0965f
C2116 _10_ net13 0.00151f
C2117 _50_/a_223_47# net4 0.0107f
C2118 net9 net17 1.26e-20
C2119 _29_/a_29_53# _35_/a_226_47# 2.64e-19
C2120 _35_/a_76_199# _11_ 6.99e-22
C2121 VPWR _42_/a_296_53# -6.37e-20
C2122 net5 b[0] 3.39e-19
C2123 _17_ net3 0.0698f
C2124 p[3] input9/a_75_212# 0.0162f
C2125 net9 net15 8.49e-20
C2126 net5 net7 0.195f
C2127 _12_ _26_/a_29_53# 0.00243f
C2128 VPWR _35_/a_226_47# 0.00159f
C2129 _48_/a_27_47# _09_ 0.00541f
C2130 _30_/a_109_53# net1 0.0297f
C2131 output17/a_27_47# p[0] 0.00805f
C2132 _01_ _32_/a_27_47# 0.0266f
C2133 _12_ net6 0.0891f
C2134 _01_ _49_/a_201_297# 0.0105f
C2135 _12_ b[1] 0.00685f
C2136 net19 input5/a_664_47# 1.38e-21
C2137 _36_/a_27_47# _32_/a_27_47# 0.011f
C2138 _24_ _21_ 0.0388f
C2139 _32_/a_27_47# _22_ 1.76e-19
C2140 net13 net14 2.21e-21
C2141 net10 net9 0.111f
C2142 _30_/a_109_53# _21_ 3.31e-20
C2143 _23_ _25_ 0.00465f
C2144 VGND _29_/a_29_53# 0.0544f
C2145 _05_ _00_ 5.03e-22
C2146 _22_ _49_/a_201_297# 2.45e-20
C2147 net17 p[10] 0.181f
C2148 _30_/a_109_53# net8 1.76e-20
C2149 _40_/a_109_297# _06_ 0.00175f
C2150 _50_/a_27_47# net10 3.78e-21
C2151 _52_/a_93_21# _24_ 0.0211f
C2152 input5/a_841_47# net5 0.0221f
C2153 p[8] net2 0.00972f
C2154 net13 _30_/a_392_297# 6.64e-20
C2155 p[13] p[0] 4.11e-19
C2156 input8/a_27_47# _31_/a_35_297# 0.00955f
C2157 p[10] net15 0.0101f
C2158 VGND VPWR -0.433f
C2159 VPWR _43_/a_193_413# 0.0063f
C2160 VPWR p[1] 0.0804f
C2161 _14_ _44_/a_256_47# 0.00124f
C2162 _50_/a_343_93# _15_ 0.0098f
C2163 _12_ _03_ 2.76e-20
C2164 net1 _21_ 0.0252f
C2165 _01_ _20_ 0.161f
C2166 output17/a_27_47# net2 0.0285f
C2167 _15_ input5/a_558_47# 0.00166f
C2168 _42_/a_109_93# net14 0.00351f
C2169 _52_/a_250_297# p[12] 1.84e-20
C2170 net1 net8 0.381f
C2171 _44_/a_250_297# _00_ 6.39e-20
C2172 _11_ _13_ 0.164f
C2173 input7/a_27_47# b[3] 1.21e-19
C2174 net5 net13 0.127f
C2175 _36_/a_27_47# _20_ 0.00148f
C2176 net9 net11 0.136f
C2177 _04_ net12 0.267f
C2178 _34_/a_47_47# p[7] 2.88e-19
C2179 _04_ _05_ 0.0352f
C2180 _20_ _22_ 0.183f
C2181 _30_/a_215_297# net17 4.69e-20
C2182 _41_/a_59_75# net15 1.16e-20
C2183 p[14] net3 0.00446f
C2184 _50_/a_27_47# net11 6.05e-21
C2185 net8 _27_/a_277_297# 7.99e-20
C2186 net16 _38_/a_197_47# 5.89e-19
C2187 input13/a_27_47# net9 2.42e-19
C2188 _29_/a_29_53# _06_ 0.00111f
C2189 _11_ _09_ 0.0665f
C2190 _44_/a_346_47# _14_ 3.76e-19
C2191 net8 _21_ 0.00656f
C2192 net16 p[12] 2.15e-19
C2193 p[13] net2 0.0257f
C2194 net5 _31_/a_35_297# 2.04e-21
C2195 _31_/a_285_297# net1 5.85e-19
C2196 VPWR _06_ 1.4f
C2197 _52_/a_93_21# _21_ 9.4e-19
C2198 VPWR _27_/a_205_297# 1.05e-19
C2199 _39_/a_47_47# _17_ 1.47e-20
C2200 _17_ net19 0.0269f
C2201 _33_/a_209_311# _03_ 8.38e-19
C2202 _33_/a_368_53# net10 0.00171f
C2203 _33_/a_109_93# net9 0.00211f
C2204 _16_ net2 0.00654f
C2205 net10 input10/a_27_47# 0.00321f
C2206 net5 _42_/a_109_93# 0.00109f
C2207 _44_/a_250_297# _04_ 5.57e-21
C2208 net9 net3 5.09e-20
C2209 _50_/a_343_93# _18_ 0.0276f
C2210 input2/a_27_47# p[10] 0.0108f
C2211 _30_/a_215_297# net10 0.0512f
C2212 _12_ _02_ 0.265f
C2213 _12_ _53_/a_29_53# 3.46e-20
C2214 _27_/a_27_297# net2 0.0131f
C2215 _48_/a_27_47# VPWR 0.0158f
C2216 net16 _45_/a_109_297# 5.1e-20
C2217 _42_/a_209_311# _16_ 0.00129f
C2218 VGND _24_ -0.00863f
C2219 _31_/a_285_297# net8 0.0215f
C2220 _15_ _47_/a_299_297# 0.0103f
C2221 input3/a_27_47# b[3] 0.0133f
C2222 _35_/a_226_47# net1 1.3e-20
C2223 _19_ net17 0.0211f
C2224 _27_/a_109_297# net3 5.45e-19
C2225 VGND _30_/a_109_53# -0.00695f
C2226 _27_/a_27_297# _42_/a_209_311# 4.7e-20
C2227 _40_/a_109_297# _11_ 0.00522f
C2228 net9 p[3] 0.0376f
C2229 _15_ _18_ 0.042f
C2230 _19_ net15 0.00628f
C2231 _12_ _43_/a_27_47# 2.33e-21
C2232 VGND _38_/a_303_47# 1.78e-19
C2233 _14_ _26_/a_183_297# 6.98e-22
C2234 _55_/a_217_297# net15 7.79e-19
C2235 _35_/a_226_47# _21_ 9.87e-19
C2236 _44_/a_584_47# b[3] 0.00109f
C2237 _33_/a_209_311# _08_ 0.0122f
C2238 net11 input10/a_27_47# 0.112f
C2239 p[10] net3 8.47e-19
C2240 net18 _38_/a_27_47# 0.00997f
C2241 _30_/a_215_297# input2/a_27_47# 3.51e-20
C2242 _01_ _00_ 0.00124f
C2243 _30_/a_215_297# net11 1.04e-19
C2244 p[9] _15_ 2.06e-19
C2245 _52_/a_93_21# _35_/a_226_47# 4.89e-20
C2246 _52_/a_250_297# _35_/a_76_199# 3.4e-21
C2247 _17_ output19/a_27_47# 0.00122f
C2248 VGND net1 0.513f
C2249 _36_/a_197_47# net6 6.94e-20
C2250 net1 p[1] 0.0291f
C2251 _39_/a_377_297# net6 0.00143f
C2252 _22_ _00_ 0.477f
C2253 _28_/a_109_297# VPWR -1.71e-19
C2254 _24_ _06_ 0.113f
C2255 VGND _27_/a_277_297# -4.65e-19
C2256 p[7] input9/a_75_212# 0.00102f
C2257 _50_/a_343_93# _26_/a_29_53# 2.61e-19
C2258 _03_ _49_/a_75_199# 0.0849f
C2259 p[14] net19 0.101f
C2260 _22_ _38_/a_27_47# 2.86e-19
C2261 _06_ _30_/a_109_53# 1.96e-19
C2262 VGND _21_ 0.295f
C2263 _42_/a_109_93# _44_/a_93_21# 1.25e-19
C2264 VGND net8 0.405f
C2265 _30_/a_215_297# _33_/a_109_93# 0.00104f
C2266 net8 _43_/a_193_413# 1.62e-20
C2267 _50_/a_343_93# net6 0.00214f
C2268 p[4] net13 2.34e-20
C2269 p[1] net8 0.00115f
C2270 _34_/a_377_297# net10 1.62e-19
C2271 _39_/a_47_47# input4/a_75_212# 3.1e-19
C2272 VPWR _11_ 0.352f
C2273 _52_/a_93_21# VGND -0.0175f
C2274 VPWR _37_/a_109_47# -4.38e-19
C2275 input14/a_27_47# net14 0.0232f
C2276 _52_/a_584_47# _04_ 2.5e-19
C2277 _01_ _04_ 0.119f
C2278 _15_ _26_/a_29_53# 0.00192f
C2279 p[4] input11/a_27_47# 0.0644f
C2280 _40_/a_109_297# p[8] 5.45e-19
C2281 _19_ input2/a_27_47# 5.26e-20
C2282 _36_/a_27_47# _04_ 0.00169f
C2283 net11 _19_ 6.27e-21
C2284 _25_ net13 0.00297f
C2285 _15_ net6 0.17f
C2286 _04_ _22_ 1.76e-20
C2287 _47_/a_384_47# _17_ 1.1e-20
C2288 _36_/a_27_47# _50_/a_223_47# 1.27e-20
C2289 _06_ net1 0.0115f
C2290 VGND _31_/a_285_297# -0.00136f
C2291 _50_/a_223_47# _22_ 0.031f
C2292 _30_/a_215_297# p[3] 2.31e-19
C2293 _49_/a_201_297# net15 1.41e-19
C2294 _29_/a_111_297# _09_ 5.79e-20
C2295 _52_/a_250_297# _13_ 5.43e-19
C2296 _06_ _21_ 0.143f
C2297 _49_/a_75_199# _02_ 0.0354f
C2298 p[2] _49_/a_75_199# 1.06e-19
C2299 p[14] output19/a_27_47# 0.0937f
C2300 net9 input5/a_381_47# 3.4e-19
C2301 _04_ input5/a_62_47# 0.00345f
C2302 _07_ b[3] 3.54e-20
C2303 _10_ _44_/a_346_47# 9.13e-21
C2304 _06_ net8 0.00282f
C2305 VGND _35_/a_226_47# -0.0111f
C2306 net10 _32_/a_27_47# 2.76e-20
C2307 net11 _29_/a_183_297# 3.64e-19
C2308 _44_/a_256_47# net14 0.00379f
C2309 _23_ _45_/a_193_297# 4.13e-19
C2310 _19_ net3 0.0122f
C2311 VPWR _39_/a_129_47# -9.47e-19
C2312 _55_/a_217_297# net3 5.78e-20
C2313 _52_/a_93_21# _06_ 0.0584f
C2314 _52_/a_250_297# _09_ 1.97e-20
C2315 p[10] net19 1.26e-21
C2316 _03_ _15_ 7.39e-20
C2317 net17 _20_ 4e-20
C2318 _45_/a_27_47# net4 0.024f
C2319 net6 _47_/a_299_297# 3.63e-19
C2320 _26_/a_29_53# _18_ 5.26e-20
C2321 _48_/a_27_47# _21_ 0.0121f
C2322 net2 _14_ 0.0104f
C2323 net16 _13_ 0.0198f
C2324 net5 _32_/a_197_47# 5.61e-21
C2325 net6 _18_ 0.166f
C2326 _20_ net15 0.0021f
C2327 VPWR p[8] 0.285f
C2328 _53_/a_183_297# _22_ 3.71e-20
C2329 _33_/a_209_311# _34_/a_47_47# 0.017f
C2330 _31_/a_285_297# _06_ 1.01e-20
C2331 _24_ _11_ 7.29e-20
C2332 _42_/a_209_311# _14_ 0.00142f
C2333 net16 _09_ 0.00707f
C2334 _44_/a_346_47# net14 0.00464f
C2335 _44_/a_250_297# input3/a_27_47# 2.07e-19
C2336 _29_/a_183_297# net3 7.38e-21
C2337 VGND _43_/a_193_413# -0.0147f
C2338 VGND p[1] 0.134f
C2339 _41_/a_59_75# net19 3.1e-20
C2340 _50_/a_343_93# _02_ 6.94e-19
C2341 p[9] net6 0.14f
C2342 _10_ _26_/a_183_297# 5.74e-19
C2343 VPWR _30_/a_297_297# -4.57e-19
C2344 net10 _20_ 3.23e-19
C2345 net11 _49_/a_201_297# 1.42e-19
C2346 VPWR output17/a_27_47# 0.0263f
C2347 _35_/a_226_47# _06_ 0.00487f
C2348 p[4] input12/a_27_47# 9.28e-19
C2349 net9 p[7] 8.26e-19
C2350 _03_ _18_ 7.25e-23
C2351 b[3] net7 0.00175f
C2352 _15_ _02_ 0.101f
C2353 _49_/a_315_47# _19_ 1.33e-19
C2354 _23_ net12 2.28e-21
C2355 _17_ _37_/a_27_47# 0.00277f
C2356 _40_/a_297_297# _20_ 9.18e-21
C2357 p[13] VPWR 0.209f
C2358 _10_ _38_/a_197_47# 6.29e-19
C2359 net6 _26_/a_29_53# 0.0032f
C2360 _15_ _43_/a_27_47# 8.96e-20
C2361 VPWR _16_ 0.126f
C2362 _11_ _21_ 9.98e-20
C2363 VGND _06_ 1.09f
C2364 VGND _27_/a_205_297# -3.36e-19
C2365 b[0] net4 0.00301f
C2366 _06_ _43_/a_193_413# 0.0138f
C2367 net11 _20_ 0.00128f
C2368 _11_ net8 1.81e-20
C2369 VPWR _29_/a_111_297# -5.85e-19
C2370 _45_/a_27_47# _05_ 9.34e-23
C2371 _10_ p[12] 0.109f
C2372 _27_/a_27_297# VPWR 0.0329f
C2373 input5/a_841_47# b[3] 2.04e-19
C2374 _17_ _12_ 0.0109f
C2375 _39_/a_285_47# p[12] 3.75e-19
C2376 _38_/a_109_47# net4 7.32e-19
C2377 _48_/a_27_47# VGND 0.0548f
C2378 _07_ net12 0.18f
C2379 _00_ net15 0.00147f
C2380 _07_ _05_ 1.21e-19
C2381 _54_/a_75_212# b[1] 7.35e-19
C2382 _52_/a_250_297# VPWR 0.019f
C2383 _14_ _13_ 1.47e-20
C2384 _44_/a_256_47# _44_/a_93_21# -6.6e-20
C2385 _02_ _18_ 2.96e-20
C2386 _37_/a_197_47# net2 4.74e-20
C2387 VPWR p[5] 0.14f
C2388 _10_ _45_/a_109_297# 0.00202f
C2389 _20_ net3 4.07e-19
C2390 _03_ _26_/a_29_53# 7.93e-21
C2391 input3/a_27_47# _22_ 5.13e-20
C2392 net13 b[3] 1.08e-19
C2393 _31_/a_285_47# VPWR -2.91e-19
C2394 _03_ net6 2.9e-20
C2395 _43_/a_27_47# _18_ 0.0201f
C2396 p[7] input10/a_27_47# 4.26e-20
C2397 VPWR net16 0.518f
C2398 _04_ net17 0.0218f
C2399 _03_ b[1] 0.00143f
C2400 input11/a_27_47# b[3] 1.21e-19
C2401 _15_ _55_/a_80_21# 0.107f
C2402 VPWR _42_/a_368_53# -3.03e-19
C2403 _44_/a_346_47# _44_/a_93_21# -5.12e-20
C2404 _35_/a_556_47# _08_ 7.71e-19
C2405 _37_/a_27_47# p[14] 1.37e-19
C2406 _03_ _54_/a_75_212# 5.45e-21
C2407 _04_ net15 0.0569f
C2408 input1/a_75_212# p[10] 0.00372f
C2409 _31_/a_35_297# b[3] 9.28e-20
C2410 net2 _47_/a_81_21# 4.95e-19
C2411 VGND _28_/a_109_297# -9.87e-19
C2412 _48_/a_27_47# _06_ 0.0251f
C2413 net13 net4 2.48e-19
C2414 input3/a_27_47# input5/a_62_47# 0.00179f
C2415 _30_/a_297_297# net1 7.34e-20
C2416 _10_ net2 2.65e-19
C2417 output17/a_27_47# net1 8.12e-19
C2418 _01_ _32_/a_109_47# 0.00129f
C2419 _42_/a_109_93# b[3] 6.56e-19
C2420 _40_/a_109_297# _14_ -1.78e-33
C2421 net10 _04_ 0.121f
C2422 net5 p[12] 0.00365f
C2423 _23_ net18 -4.05e-24
C2424 net12 net7 1.57e-19
C2425 _05_ net7 0.0129f
C2426 VGND _11_ 0.0908f
C2427 _02_ _26_/a_29_53# 0.0466f
C2428 _11_ _43_/a_193_413# 5.45e-19
C2429 _30_/a_297_297# net8 2.42e-21
C2430 VGND _37_/a_109_47# -7.9e-19
C2431 _08_ b[1] 1.17e-19
C2432 output17/a_27_47# net8 0.0043f
C2433 _10_ _35_/a_76_199# 7.19e-20
C2434 _52_/a_250_297# _24_ 3.03e-19
C2435 net13 _30_/a_465_297# 6.36e-20
C2436 p[13] net1 2.13e-19
C2437 _12_ input4/a_75_212# 2.09e-20
C2438 net6 _02_ 0.00427f
C2439 net11 _38_/a_27_47# 1.68e-20
C2440 _53_/a_29_53# net6 2.11e-20
C2441 VPWR _43_/a_297_47# -2.11e-19
C2442 _53_/a_29_53# b[1] 3.63e-19
C2443 b[1] _02_ 0.00178f
C2444 p[2] b[1] 0.0428f
C2445 net2 net14 0.151f
C2446 _55_/a_80_21# _18_ 1.44e-20
C2447 p[13] _27_/a_277_297# 4.24e-20
C2448 _23_ _36_/a_27_47# 0.00118f
C2449 net5 _45_/a_109_297# 0.0184f
C2450 _54_/a_75_212# _02_ 6.6e-20
C2451 _23_ _22_ 0.0187f
C2452 _50_/a_429_93# _15_ 6.82e-19
C2453 _12_ net9 4.39e-22
C2454 _27_/a_27_297# net1 6.05e-21
C2455 net6 _43_/a_27_47# 9.07e-20
C2456 _42_/a_209_311# net14 0.0238f
C2457 VPWR output18/a_27_47# 0.0689f
C2458 net16 _24_ 6.93e-19
C2459 _15_ input5/a_664_47# 9.15e-22
C2460 p[13] net8 0.0034f
C2461 _50_/a_27_47# _12_ 0.00354f
C2462 _00_ net3 2.12e-19
C2463 VPWR p[6] 0.079f
C2464 _04_ input2/a_27_47# 4.5e-21
C2465 _03_ _08_ 0.0144f
C2466 _04_ net11 0.078f
C2467 _39_/a_47_47# _20_ 2.3e-20
C2468 _20_ net19 1.29e-19
C2469 _16_ net8 0.00624f
C2470 VPWR _52_/a_256_47# -9.47e-19
C2471 VPWR _48_/a_181_47# -3.35e-19
C2472 net16 _38_/a_303_47# 6.47e-19
C2473 _45_/a_27_47# _22_ 0.0131f
C2474 VGND _39_/a_129_47# -0.00126f
C2475 _11_ _06_ 0.493f
C2476 _03_ _02_ 0.00474f
C2477 _27_/a_27_297# net8 0.0108f
C2478 p[11] input3/a_27_47# 0.014f
C2479 VPWR _14_ 0.186f
C2480 input12/a_27_47# b[3] 1.21e-19
C2481 net5 net2 0.0616f
C2482 _07_ _22_ 1.19e-20
C2483 net13 net12 0.363f
C2484 net13 _05_ 0.192f
C2485 _33_/a_209_311# net9 4.33e-20
C2486 _33_/a_109_93# _04_ 0.0299f
C2487 VGND p[8] 0.35f
C2488 p[8] _43_/a_193_413# 3.24e-19
C2489 net17 input7/a_27_47# 4.99e-20
C2490 _04_ _49_/a_544_297# 0.00204f
C2491 net5 _42_/a_209_311# 3.27e-21
C2492 _04_ net3 0.112f
C2493 _10_ _13_ 0.0621f
C2494 _52_/a_93_21# _52_/a_250_297# -6.97e-22
C2495 input7/a_27_47# net15 1.88e-19
C2496 _39_/a_285_47# _13_ 0.00451f
C2497 _18_ input5/a_664_47# 1.09e-20
C2498 net5 _35_/a_76_199# 3.38e-19
C2499 _50_/a_343_93# _17_ 0.0015f
C2500 _31_/a_35_297# _05_ 0.00649f
C2501 _31_/a_285_47# net8 0.00129f
C2502 net16 _21_ 1.89e-19
C2503 VGND _30_/a_297_297# -4.43e-19
C2504 _10_ _09_ 0.0222f
C2505 _17_ input5/a_558_47# 2.13e-21
C2506 _08_ _02_ 2.26e-20
C2507 VGND output17/a_27_47# 0.00231f
C2508 VPWR _55_/a_472_297# 0.00488f
C2509 _41_/a_59_75# _12_ 0.00101f
C2510 _04_ p[3] 5.34e-19
C2511 _53_/a_29_53# _02_ 0.0388f
C2512 p[2] _02_ 7.08e-19
C2513 input15/a_27_47# p[12] 5.48e-19
C2514 _17_ _15_ 0.0752f
C2515 input14/a_27_47# b[3] 0.0211f
C2516 _34_/a_47_47# b[1] 4.35e-19
C2517 _01_ net7 0.233f
C2518 _28_/a_109_297# _11_ 6.29e-19
C2519 _06_ p[8] 0.00489f
C2520 _52_/a_250_297# _35_/a_226_47# 2.63e-20
C2521 p[13] VGND 0.0891f
C2522 _43_/a_27_47# _02_ 1.88e-21
C2523 _36_/a_303_47# net6 1.25e-19
C2524 _39_/a_47_47# _00_ 1.85e-20
C2525 net2 _44_/a_93_21# 0.0273f
C2526 _22_ net7 2.73e-20
C2527 VGND _16_ -0.00582f
C2528 _16_ _43_/a_193_413# 0.0261f
C2529 input3/a_27_47# net15 6.19e-20
C2530 _44_/a_250_297# _42_/a_109_93# 6.38e-19
C2531 VGND _29_/a_111_297# -1.9e-19
C2532 net9 _49_/a_75_199# 0.00382f
C2533 VGND _27_/a_27_297# -0.0157f
C2534 _04_ _49_/a_315_47# 7.71e-19
C2535 _42_/a_209_311# _44_/a_93_21# 2.21e-19
C2536 _27_/a_27_297# p[1] 2.27e-19
C2537 input7/a_27_47# input2/a_27_47# 1.62e-19
C2538 _47_/a_384_47# _20_ 1.72e-19
C2539 _30_/a_215_297# _33_/a_209_311# 1.56e-19
C2540 net1 p[6] 3.12e-20
C2541 _50_/a_429_93# net6 6.18e-19
C2542 _34_/a_129_47# net10 0.003f
C2543 _34_/a_47_47# _03_ 4.5e-20
C2544 net7 input5/a_62_47# 2.04e-19
C2545 net5 _13_ 0.0381f
C2546 _52_/a_250_297# VGND -0.00314f
C2547 VPWR _37_/a_197_47# -3.27e-19
C2548 _17_ _18_ 0.271f
C2549 _21_ output18/a_27_47# 0.00103f
C2550 VGND p[5] 0.15f
C2551 p[6] _21_ 0.00203f
C2552 _36_/a_109_47# _04_ 2.39e-19
C2553 input15/a_27_47# net2 0.00296f
C2554 net12 input12/a_27_47# 0.0297f
C2555 _04_ net19 2.07e-20
C2556 net5 _09_ 5.18e-19
C2557 p[13] _27_/a_205_297# 5.22e-20
C2558 p[10] _49_/a_75_199# 2.29e-20
C2559 _16_ _06_ 0.00162f
C2560 _45_/a_27_47# _35_/a_489_413# 3.89e-21
C2561 p[14] _15_ 5.32e-19
C2562 _17_ p[9] 1.03e-20
C2563 VGND net16 0.144f
C2564 _01_ net13 0.00228f
C2565 _10_ _29_/a_29_53# 5.17e-19
C2566 _02_ _55_/a_80_21# 0.164f
C2567 _52_/a_93_21# _52_/a_256_47# -6.6e-20
C2568 _06_ _29_/a_111_297# 6.74e-20
C2569 net8 _14_ 4.23e-19
C2570 VGND _42_/a_368_53# -4.05e-19
C2571 _50_/a_343_93# net9 6.64e-19
C2572 _36_/a_27_47# net13 0.0488f
C2573 VPWR _47_/a_81_21# 0.00889f
C2574 net13 _22_ 4.63e-20
C2575 _34_/a_129_47# net11 0.00242f
C2576 _34_/a_285_47# net12 8.07e-20
C2577 _07_ _35_/a_489_413# 0.00429f
C2578 _34_/a_47_47# _08_ 0.00123f
C2579 _50_/a_343_93# _50_/a_27_47# -7.11e-33
C2580 _34_/a_285_47# _05_ 7.85e-21
C2581 _10_ VPWR 0.577f
C2582 net9 input5/a_558_47# 4.42e-19
C2583 VPWR _39_/a_285_47# -9.53e-19
C2584 _43_/a_27_47# _55_/a_80_21# 1.56e-19
C2585 _31_/a_35_297# _01_ 4.27e-19
C2586 _34_/a_47_47# _02_ 1.09e-19
C2587 _52_/a_250_297# _06_ 0.0058f
C2588 _34_/a_47_47# _53_/a_29_53# 5.88e-22
C2589 net9 _15_ 0.00113f
C2590 _11_ p[8] 0.0039f
C2591 p[8] _37_/a_109_47# 3.95e-21
C2592 input9/a_75_212# b[1] 2.46e-19
C2593 _50_/a_27_47# _15_ 5.65e-19
C2594 net5 _32_/a_303_47# 7.18e-21
C2595 _29_/a_29_53# net14 1.61e-20
C2596 input8/a_27_47# VPWR 0.0863f
C2597 _23_ net10 0.00216f
C2598 _42_/a_109_93# _22_ 1.21e-19
C2599 _17_ net6 3.12e-19
C2600 net16 _06_ 0.0511f
C2601 VPWR net14 0.182f
C2602 _47_/a_384_47# _00_ 5.15e-20
C2603 input3/a_27_47# net3 0.0299f
C2604 p[10] input5/a_558_47# 1.09e-19
C2605 VGND _43_/a_297_47# -1.33e-19
C2606 input6/a_27_47# p[12] 2.78e-19
C2607 _18_ input4/a_75_212# 4.36e-19
C2608 _28_/a_109_297# _16_ 1.26e-19
C2609 _02_ input5/a_664_47# 0.00187f
C2610 _03_ input9/a_75_212# 9.32e-20
C2611 VGND output18/a_27_47# 0.0581f
C2612 p[9] p[14] 0.415f
C2613 _50_/a_343_93# _41_/a_59_75# 6.13e-22
C2614 VGND p[6] 0.13f
C2615 net5 _29_/a_29_53# 8.1e-20
C2616 _44_/a_250_297# input14/a_27_47# 8.25e-21
C2617 net9 _18_ 1.51e-19
C2618 VGND _52_/a_256_47# -0.00161f
C2619 _19_ _49_/a_75_199# 0.0206f
C2620 _07_ net10 0.0605f
C2621 _50_/a_27_47# _18_ 0.0665f
C2622 VGND _48_/a_181_47# 3.03e-19
C2623 _10_ _24_ 0.00484f
C2624 _23_ net11 0.0461f
C2625 _11_ _16_ 4.42e-20
C2626 _23_ b[2] 2.87e-20
C2627 _12_ _20_ 3.9e-19
C2628 VGND _14_ 0.226f
C2629 net5 VPWR 0.613f
C2630 _14_ _43_/a_193_413# 0.0297f
C2631 _41_/a_59_75# _15_ 0.0139f
C2632 net6 _26_/a_111_297# 1.12e-19
C2633 _10_ _38_/a_303_47# 7.36e-19
C2634 _06_ _43_/a_297_47# 4.81e-20
C2635 b[3] p[12] 7.54e-20
C2636 _45_/a_27_47# net11 3.64e-20
C2637 net17 net7 0.2f
C2638 p[0] b[3] 0.0791f
C2639 _25_ _09_ 1.49e-19
C2640 net1 _47_/a_81_21# 1.58e-21
C2641 _38_/a_197_47# net4 7.64e-19
C2642 net2 input6/a_27_47# 0.0047f
C2643 _35_/a_226_297# _04_ 4.51e-19
C2644 _06_ output18/a_27_47# 0.0114f
C2645 p[2] input9/a_75_212# 7.58e-20
C2646 p[14] net6 0.00237f
C2647 _10_ net1 4.34e-19
C2648 _07_ net11 0.0206f
C2649 net15 net7 2.91e-19
C2650 _06_ p[6] 0.00262f
C2651 _06_ _52_/a_256_47# 0.00207f
C2652 net4 p[12] 0.0233f
C2653 VGND _55_/a_472_297# -0.00188f
C2654 net6 input4/a_75_212# 0.0273f
C2655 _06_ _48_/a_181_47# 6.4e-19
C2656 _37_/a_303_47# net2 4.41e-19
C2657 _41_/a_59_75# _47_/a_299_297# 0.00146f
C2658 net16 _11_ 0.172f
C2659 net9 _26_/a_29_53# 0.00343f
C2660 net8 _47_/a_81_21# 2.08e-21
C2661 _17_ _02_ 0.00482f
C2662 _10_ _21_ 0.00421f
C2663 _06_ _14_ 0.0556f
C2664 net13 _35_/a_489_413# 7.36e-20
C2665 _48_/a_27_47# p[6] 2.32e-19
C2666 input3/a_27_47# net19 0.00105f
C2667 _45_/a_193_297# p[12] 1.55e-20
C2668 _10_ net8 5.86e-19
C2669 _50_/a_27_47# _26_/a_29_53# 5.56e-19
C2670 p[13] p[8] 0.00172f
C2671 _37_/a_27_47# _00_ 6.15e-20
C2672 net10 net7 1.65e-36
C2673 input8/a_27_47# net1 0.0347f
C2674 _07_ _33_/a_109_93# 3.2e-19
C2675 _19_ _15_ 1.46e-20
C2676 net9 b[1] 3.31e-20
C2677 _45_/a_109_297# net4 6.43e-20
C2678 _16_ p[8] 1.59e-19
C2679 _10_ _52_/a_93_21# 0.00534f
C2680 _50_/a_27_47# net6 0.0428f
C2681 input5/a_841_47# net15 0.00585f
C2682 _15_ _55_/a_217_297# 0.0474f
C2683 net1 net14 6.64e-20
C2684 _17_ _43_/a_27_47# 0.00131f
C2685 VPWR _44_/a_93_21# 0.005f
C2686 net5 _24_ 5.83e-20
C2687 net2 b[3] 0.318f
C2688 _31_/a_117_297# b[3] 1.21e-20
C2689 net5 _30_/a_109_53# 5.84e-22
C2690 _41_/a_59_75# p[9] 1.02e-19
C2691 _27_/a_277_297# net14 5.1e-19
C2692 p[13] output17/a_27_47# 0.00122f
C2693 _45_/a_465_47# p[12] 5.2e-20
C2694 input8/a_27_47# net8 0.0181f
C2695 _01_ _32_/a_197_47# 0.00156f
C2696 _12_ _00_ 0.00396f
C2697 net13 net17 5.21e-20
C2698 net14 _21_ 7.17e-21
C2699 _42_/a_209_311# b[3] 8.61e-19
C2700 VGND _48_/a_109_47# 9.44e-19
C2701 net8 net14 0.0516f
C2702 net13 net15 8.84e-19
C2703 b[0] b[2] 0.0783f
C2704 input2/a_27_47# net7 0.00213f
C2705 _12_ _38_/a_27_47# 0.0527f
C2706 _03_ net9 0.15f
C2707 net11 net7 1.77e-19
C2708 b[1] p[10] 0.2f
C2709 VGND _37_/a_197_47# -4.58e-19
C2710 _10_ _35_/a_226_47# 1.25e-19
C2711 VPWR input15/a_27_47# 0.0113f
C2712 _31_/a_35_297# net17 0.0514f
C2713 input3/a_27_47# output19/a_27_47# 4.77e-21
C2714 net5 net1 0.0772f
C2715 VPWR p[4] 0.118f
C2716 input8/a_27_47# _31_/a_285_297# 1.04e-19
C2717 _20_ _49_/a_75_199# 0.0233f
C2718 _03_ _27_/a_109_297# 1.97e-20
C2719 VPWR _43_/a_369_47# -3.75e-19
C2720 _50_/a_343_93# _32_/a_27_47# 6.48e-20
C2721 _53_/a_111_297# b[1] 2.85e-20
C2722 _28_/a_109_297# _14_ 5.66e-19
C2723 _42_/a_109_93# net17 3.1e-21
C2724 _23_ _36_/a_109_47# 3.44e-19
C2725 net13 net10 0.375f
C2726 _23_ _39_/a_47_47# 5.24e-21
C2727 _50_/a_515_93# _15_ 0.00147f
C2728 _41_/a_59_75# net6 0.0373f
C2729 _12_ _04_ 1.42e-19
C2730 _17_ _55_/a_80_21# 7.64e-21
C2731 p[13] _27_/a_27_297# 4.67e-19
C2732 VPWR _25_ 0.0829f
C2733 net5 _21_ 0.00784f
C2734 _49_/a_544_297# net7 2.72e-19
C2735 _42_/a_109_93# net15 4.62e-19
C2736 net5 net8 0.48f
C2737 _42_/a_296_53# net14 2.18e-19
C2738 _50_/a_223_47# _12_ 0.00327f
C2739 net3 net7 7.45e-20
C2740 b[1] input10/a_27_47# 8.3e-19
C2741 _32_/a_27_47# _15_ 1.19e-19
C2742 _27_/a_27_297# _16_ 3.74e-22
C2743 _30_/a_215_297# net6 3.3e-21
C2744 _03_ p[10] 8.74e-20
C2745 VGND _47_/a_81_21# -0.0112f
C2746 net9 _08_ 7.71e-21
C2747 _06_ _48_/a_109_47# 9.47e-19
C2748 _30_/a_215_297# b[1] 3.95e-20
C2749 _10_ VGND 1.11f
C2750 _52_/a_93_21# net5 0.0124f
C2751 _11_ _14_ 0.0415f
C2752 VPWR _52_/a_346_47# -0.00109f
C2753 input1/a_75_212# input7/a_27_47# 3.2e-20
C2754 _54_/a_75_212# input10/a_27_47# 1.17e-22
C2755 _31_/a_35_297# net10 3.95e-20
C2756 _10_ _43_/a_193_413# 0.0174f
C2757 _05_ _45_/a_109_297# 2.79e-22
C2758 VGND _39_/a_285_47# -0.0046f
C2759 _45_/a_27_47# _39_/a_47_47# 1.31e-19
C2760 net9 _02_ 0.00611f
C2761 p[2] net9 1.4e-20
C2762 _50_/a_27_47# _02_ 2.09e-19
C2763 _50_/a_343_93# _20_ 0.00826f
C2764 net13 net11 0.093f
C2765 _33_/a_209_311# _04_ 0.00133f
C2766 _40_/a_191_297# net2 0.00143f
C2767 input8/a_27_47# VGND 0.0573f
C2768 input13/a_27_47# net13 0.00139f
C2769 input8/a_27_47# p[1] 5.13e-20
C2770 net11 input11/a_27_47# 0.00318f
C2771 _30_/a_215_297# _03_ 0.0393f
C2772 input14/a_27_47# p[11] 3.98e-20
C2773 VGND net14 0.441f
C2774 net14 _43_/a_193_413# 1.11e-19
C2775 p[1] net14 0.0025f
C2776 _03_ _49_/a_208_47# 3.86e-19
C2777 _15_ _20_ 0.691f
C2778 _31_/a_35_297# input2/a_27_47# 0.00136f
C2779 net2 _05_ 4.03e-20
C2780 output16/a_27_47# net6 1.5e-19
C2781 _32_/a_27_47# _18_ 1.18e-20
C2782 _06_ _47_/a_81_21# 0.0388f
C2783 output16/a_27_47# b[1] 6.65e-20
C2784 VGND _30_/a_392_297# 7.67e-19
C2785 net13 _33_/a_109_93# 0.0254f
C2786 p[10] _02_ 1.8e-19
C2787 _10_ _06_ 1.14f
C2788 VPWR _55_/a_300_47# -4.61e-19
C2789 net13 _49_/a_544_297# 3.43e-19
C2790 _13_ net4 0.212f
C2791 _06_ _39_/a_285_47# 1.23e-20
C2792 net13 net3 3.25e-21
C2793 _22_ _26_/a_183_297# 0.00184f
C2794 _49_/a_315_47# net7 0.00706f
C2795 _53_/a_111_297# _02_ 9.57e-20
C2796 p[8] _14_ 0.00748f
C2797 _33_/a_368_53# _08_ 5.04e-19
C2798 _10_ _48_/a_27_47# 4.55e-19
C2799 _35_/a_76_199# net12 0.0132f
C2800 _35_/a_76_199# _05_ 0.00238f
C2801 _09_ net4 0.00262f
C2802 _34_/a_377_297# b[1] 6.01e-20
C2803 net13 p[3] 0.00174f
C2804 net5 VGND 1.2f
C2805 _44_/a_250_297# net2 0.0169f
C2806 net5 _43_/a_193_413# 1.39e-20
C2807 _20_ _47_/a_299_297# 0.002f
C2808 _03_ _19_ 0.0019f
C2809 _39_/a_47_47# b[0] 2.04e-19
C2810 p[2] input10/a_27_47# 1.02e-20
C2811 _45_/a_193_297# _09_ 0.00961f
C2812 net10 input12/a_27_47# 0.00182f
C2813 _06_ net14 1.94e-19
C2814 net14 _27_/a_205_297# 3.63e-19
C2815 _30_/a_215_297# _02_ 3.58e-21
C2816 _20_ _18_ 0.0151f
C2817 _42_/a_109_93# net3 0.0423f
C2818 _49_/a_208_47# _02_ 0.00193f
C2819 _45_/a_465_47# _13_ 0.00134f
C2820 _04_ _49_/a_75_199# 0.0782f
C2821 VPWR input6/a_27_47# 0.00162f
C2822 _50_/a_515_93# net6 4.7e-19
C2823 _50_/a_343_93# _00_ 0.102f
C2824 _07_ p[7] 0.00227f
C2825 _45_/a_465_47# _09_ 2.77e-19
C2826 _22_ p[12] 2.13e-21
C2827 _34_/a_285_47# net10 0.0454f
C2828 _34_/a_377_297# _03_ 3.13e-20
C2829 _34_/a_47_47# net9 1.41e-20
C2830 net7 input5/a_381_47# 4.91e-19
C2831 VPWR _37_/a_303_47# -3.13e-19
C2832 _25_ _21_ 0.00164f
C2833 _03_ _29_/a_183_297# 7.36e-19
C2834 _10_ _28_/a_109_297# 4.34e-19
C2835 _15_ _00_ 0.207f
C2836 net11 input12/a_27_47# 0.00246f
C2837 _16_ _14_ 0.0584f
C2838 net5 _06_ 0.41f
C2839 _45_/a_109_297# _22_ 0.0426f
C2840 _19_ _02_ 0.213f
C2841 _11_ _47_/a_81_21# 0.0454f
C2842 _27_/a_27_297# _14_ 1.66e-21
C2843 _05_ _13_ 2.57e-20
C2844 _02_ _55_/a_217_297# 6.01e-19
C2845 _10_ _11_ 0.176f
C2846 _52_/a_93_21# _52_/a_346_47# -5.12e-20
C2847 p[6] p[5] 0.304f
C2848 VPWR b[3] 0.48f
C2849 VGND _44_/a_93_21# -0.0223f
C2850 _36_/a_109_47# net13 0.00126f
C2851 p[0] input5/a_62_47# 1.39e-19
C2852 _44_/a_93_21# _43_/a_193_413# 0.0161f
C2853 _20_ _26_/a_29_53# 0.00447f
C2854 net12 _09_ 0.0374f
C2855 net9 input5/a_664_47# 5.29e-19
C2856 _04_ input5/a_558_47# 1.25e-20
C2857 _05_ _09_ 0.0683f
C2858 net16 output18/a_27_47# 3.45e-19
C2859 _03_ _32_/a_27_47# 1.9e-19
C2860 _43_/a_27_47# _55_/a_217_297# 2.18e-19
C2861 _01_ net2 2.72e-19
C2862 _20_ net6 9.69e-20
C2863 _03_ _49_/a_201_297# 0.00842f
C2864 _04_ _15_ 3.61e-20
C2865 b[1] _20_ 3.48e-20
C2866 _00_ _47_/a_299_297# 7.59e-21
C2867 _16_ _55_/a_472_297# 3.71e-19
C2868 p[8] _37_/a_197_47# 1.03e-19
C2869 net2 _22_ 1.93e-20
C2870 VPWR net4 1.07f
C2871 _50_/a_223_47# _15_ 0.00698f
C2872 _01_ _42_/a_209_311# 1.58e-19
C2873 _00_ _18_ 0.157f
C2874 _11_ net14 5e-19
C2875 _37_/a_109_47# net14 1.71e-19
C2876 VGND input15/a_27_47# 0.0156f
C2877 _42_/a_109_93# net19 0.0448f
C2878 _42_/a_209_311# _22_ 1.72e-19
C2879 VPWR _45_/a_193_297# -0.00859f
C2880 _01_ _35_/a_76_199# 3.08e-21
C2881 input15/a_27_47# _43_/a_193_413# 1.62e-20
C2882 VGND p[4] 0.332f
C2883 _10_ _39_/a_129_47# 2.51e-19
C2884 VGND _43_/a_369_47# -8.43e-19
C2885 _35_/a_76_199# _36_/a_27_47# 3.22e-19
C2886 _43_/a_193_413# _43_/a_369_47# -1.25e-19
C2887 _35_/a_76_199# _22_ 6.58e-21
C2888 net2 input5/a_62_47# 0.0197f
C2889 _17_ p[14] 5.46e-21
C2890 VPWR _30_/a_465_297# -4.57e-19
C2891 _03_ _20_ 0.0794f
C2892 p[8] _47_/a_81_21# 3.81e-19
C2893 net9 input9/a_75_212# 0.0247f
C2894 VGND _25_ 0.199f
C2895 _10_ p[8] 9.43e-19
C2896 _32_/a_27_47# _02_ 0.00247f
C2897 _42_/a_109_93# input5/a_381_47# 0.00763f
C2898 _50_/a_223_47# _47_/a_299_297# 2.74e-20
C2899 _23_ _12_ 0.00743f
C2900 VPWR _45_/a_465_47# -5.05e-19
C2901 p[2] _49_/a_201_297# 4.58e-20
C2902 _04_ _18_ 1.94e-21
C2903 _55_/a_80_21# _55_/a_217_297# 1.42e-32
C2904 net5 _11_ 0.207f
C2905 VGND _52_/a_346_47# -0.00175f
C2906 _30_/a_109_53# b[3] 1.92e-20
C2907 _50_/a_223_47# _18_ 0.0367f
C2908 input1/a_75_212# net7 3.77e-19
C2909 _17_ net9 2.89e-23
C2910 _32_/a_27_47# _43_/a_27_47# 2.01e-20
C2911 _10_ _30_/a_297_297# 1.25e-20
C2912 _14_ _43_/a_297_47# 9.11e-19
C2913 _17_ _50_/a_27_47# 3.93e-20
C2914 _06_ input15/a_27_47# 4.73e-19
C2915 _45_/a_27_47# _12_ 0.0867f
C2916 _00_ _26_/a_29_53# 0.0466f
C2917 _42_/a_109_93# output19/a_27_47# 1.56e-20
C2918 net13 p[7] 0.00514f
C2919 _29_/a_29_53# net12 0.0132f
C2920 VPWR _40_/a_191_297# -6.82e-19
C2921 _29_/a_29_53# _05_ 3.79e-20
C2922 _06_ _43_/a_369_47# -2.02e-19
C2923 p[8] net14 0.013f
C2924 _24_ net4 8.65e-20
C2925 p[6] _48_/a_181_47# 1.44e-20
C2926 net6 _00_ 0.00178f
C2927 _07_ _12_ 2.94e-23
C2928 p[7] input11/a_27_47# 4.26e-20
C2929 net1 b[3] 7.79e-20
C2930 _06_ _25_ 0.144f
C2931 VPWR net12 0.82f
C2932 _20_ _02_ 0.1f
C2933 net18 _09_ 1.97e-21
C2934 VPWR _05_ 0.127f
C2935 _38_/a_303_47# net4 5.95e-19
C2936 _44_/a_256_47# net3 0.00101f
C2937 input7/a_27_47# input5/a_558_47# 1.22e-20
C2938 b[1] _38_/a_27_47# 4.87e-19
C2939 _22_ _13_ 0.00309f
C2940 b[3] _27_/a_277_297# 2.46e-20
C2941 net5 _39_/a_129_47# 0.00344f
C2942 _10_ _16_ 0.00486f
C2943 _06_ _52_/a_346_47# 0.0031f
C2944 p[11] net2 0.0122f
C2945 _01_ _09_ 4.69e-21
C2946 _54_/a_75_212# _38_/a_27_47# 2.67e-19
C2947 VGND _55_/a_300_47# -0.00109f
C2948 b[3] _21_ 2.41e-21
C2949 _20_ _43_/a_27_47# 0.0124f
C2950 net8 b[3] 0.00179f
C2951 _04_ _26_/a_29_53# 2.3e-21
C2952 _19_ input5/a_664_47# 2.19e-21
C2953 _22_ _09_ 0.0279f
C2954 net13 _35_/a_226_297# 6.88e-19
C2955 _30_/a_215_297# input9/a_75_212# 6.24e-21
C2956 _50_/a_223_47# _26_/a_29_53# 0.00124f
C2957 net5 p[8] 5.53e-19
C2958 _11_ _44_/a_93_21# 4.78e-20
C2959 net15 p[12] 2.99e-19
C2960 _04_ net6 2.61e-20
C2961 _03_ _00_ 2.31e-20
C2962 _44_/a_346_47# net3 8.04e-19
C2963 VPWR _44_/a_250_297# 0.0231f
C2964 _07_ _33_/a_209_311# 0.00859f
C2965 _04_ b[1] 6.5e-19
C2966 _50_/a_223_47# net6 0.0194f
C2967 _10_ _52_/a_250_297# 0.00368f
C2968 p[13] net14 5.21e-19
C2969 _41_/a_59_75# _17_ 0.00149f
C2970 _21_ net4 0.00535f
C2971 _16_ net14 0.00266f
C2972 _13_ _45_/a_205_47# 7.51e-20
C2973 net5 output17/a_27_47# 5.01e-20
C2974 input14/a_27_47# net19 1.44e-19
C2975 _55_/a_472_297# _14_ 0.00192f
C2976 b[0] _12_ 2.61e-20
C2977 _52_/a_93_21# net4 7.93e-20
C2978 _01_ _32_/a_303_47# 8.58e-19
C2979 _27_/a_27_297# net14 0.0118f
C2980 _42_/a_296_53# b[3] 2.07e-20
C2981 VGND input6/a_27_47# -0.00259f
C2982 _10_ net16 0.0338f
C2983 input5/a_841_47# _37_/a_27_47# 4.64e-20
C2984 _06_ _55_/a_300_47# 2.5e-20
C2985 input3/a_27_47# _15_ 7.53e-19
C2986 _11_ input15/a_27_47# 4.4e-19
C2987 net16 _39_/a_285_47# 1.29e-19
C2988 _52_/a_93_21# _45_/a_193_297# 6.01e-19
C2989 _12_ _38_/a_109_47# 0.00179f
C2990 _03_ _04_ 0.586f
C2991 _30_/a_109_53# net12 4.25e-20
C2992 _20_ _55_/a_80_21# 0.0291f
C2993 _30_/a_109_53# _05_ 0.033f
C2994 VGND _37_/a_303_47# -1.63e-19
C2995 _50_/a_223_47# _03_ 1.41e-21
C2996 p[13] net5 0.008f
C2997 net17 net2 0.261f
C2998 _31_/a_117_297# net17 0.00149f
C2999 _00_ _02_ 0.0269f
C3000 VPWR _43_/a_469_47# -2.75e-19
C3001 p[7] input12/a_27_47# 1.95e-19
C3002 _48_/a_109_47# p[6] 7.26e-22
C3003 _53_/a_183_297# b[1] 4.4e-20
C3004 net5 _16_ 1.99e-20
C3005 _11_ _25_ 7.05e-19
C3006 net2 net15 0.324f
C3007 _42_/a_209_311# net17 1.04e-21
C3008 _17_ _19_ 8.82e-21
C3009 _53_/a_29_53# _38_/a_27_47# 1.29e-19
C3010 _38_/a_27_47# _02_ 0.00103f
C3011 p[8] _44_/a_93_21# 5.51e-19
C3012 _50_/a_615_93# _15_ 0.00183f
C3013 net5 _27_/a_27_297# 3.48e-19
C3014 VPWR net18 0.104f
C3015 _29_/a_29_53# _01_ 8.33e-20
C3016 _00_ _43_/a_27_47# 0.0431f
C3017 _07_ _49_/a_75_199# 4.05e-21
C3018 _42_/a_209_311# net15 0.0157f
C3019 _42_/a_368_53# net14 7.39e-19
C3020 input14/a_27_47# output19/a_27_47# 0.0101f
C3021 net12 net1 1.17e-19
C3022 VGND b[3] 0.222f
C3023 net1 _05_ 0.151f
C3024 _29_/a_29_53# _36_/a_27_47# 6.92e-20
C3025 p[1] b[3] 0.045f
C3026 _06_ input6/a_27_47# 2.85e-19
C3027 _41_/a_59_75# p[14] 5.13e-20
C3028 _29_/a_29_53# _22_ 2.24e-21
C3029 _04_ _08_ 5.99e-19
C3030 _34_/a_285_47# p[7] 9.55e-20
C3031 _35_/a_226_47# _45_/a_193_297# 8.15e-21
C3032 _52_/a_250_297# net5 0.018f
C3033 VPWR _52_/a_584_47# -9.47e-19
C3034 _10_ _43_/a_297_47# 0.00118f
C3035 _01_ VPWR 0.521f
C3036 net10 net2 2.05e-20
C3037 net11 _45_/a_109_297# 7.46e-20
C3038 net13 _12_ 0.00632f
C3039 _41_/a_59_75# input4/a_75_212# 0.00153f
C3040 VPWR _36_/a_27_47# -0.00832f
C3041 _04_ _02_ 0.0541f
C3042 p[2] _04_ 1.83e-20
C3043 net12 _21_ 0.23f
C3044 VPWR _22_ 1.4f
C3045 _44_/a_346_47# net19 0.00124f
C3046 _05_ _21_ 0.0104f
C3047 net12 net8 0.00458f
C3048 _50_/a_223_47# _02_ 2.51e-20
C3049 _42_/a_109_93# _37_/a_27_47# 2.55e-20
C3050 net8 _05_ 0.0146f
C3051 VGND net4 0.564f
C3052 input15/a_27_47# p[8] 0.00758f
C3053 net5 net16 0.00476f
C3054 _35_/a_76_199# net10 0.0226f
C3055 _52_/a_93_21# _05_ 1.12e-20
C3056 p[8] _43_/a_369_47# 8.49e-20
C3057 _40_/a_297_297# net2 0.00101f
C3058 b[1] input7/a_27_47# 8.24e-19
C3059 _10_ _52_/a_256_47# 1.65e-19
C3060 _41_/a_59_75# _50_/a_27_47# 9.59e-22
C3061 VGND _45_/a_193_297# -0.00241f
C3062 _14_ _47_/a_81_21# 6.24e-20
C3063 _30_/a_215_297# net9 0.0458f
C3064 net14 _43_/a_297_47# 1.09e-21
C3065 VPWR input5/a_62_47# 0.0601f
C3066 _10_ _14_ 0.0571f
C3067 _35_/a_489_413# _09_ 0.0296f
C3068 net2 input2/a_27_47# 0.024f
C3069 _06_ b[3] 3.15e-19
C3070 _16_ _44_/a_93_21# 0.00354f
C3071 b[3] _27_/a_205_297# 3.05e-20
C3072 _31_/a_285_297# _05_ 6.12e-19
C3073 _00_ _55_/a_80_21# 5.5e-19
C3074 p[3] p[0] 0.0462f
C3075 net13 _33_/a_209_311# 0.0227f
C3076 VGND _30_/a_465_297# 0.00105f
C3077 VPWR _45_/a_205_47# -1.62e-19
C3078 _42_/a_209_311# input2/a_27_47# 1e-22
C3079 _49_/a_75_199# net7 0.09f
C3080 _24_ net18 5.57e-21
C3081 VGND _45_/a_465_47# -8.14e-19
C3082 _53_/a_183_297# _02_ 4.14e-19
C3083 _35_/a_76_199# net11 4e-19
C3084 _35_/a_226_47# net12 8.29e-19
C3085 _35_/a_226_47# _05_ 0.0134f
C3086 _06_ net4 0.281f
C3087 _34_/a_129_47# b[1] 1.01e-19
C3088 _14_ net14 0.184f
C3089 m1_7039_1799# 0 0.143f
C3090 _04_ 0 0.338f
C3091 net9 0 0.306f
C3092 _03_ 0 0.36f
C3093 net10 0 0.412f
C3094 _30_/a_109_53# 0 0.159f
C3095 _30_/a_215_297# 0 0.142f
C3096 _05_ 0 0.152f
C3097 net8 0 0.384f
C3098 _31_/a_285_297# 0 0.00137f
C3099 _31_/a_35_297# 0 0.255f
C3100 _06_ 0 0.804f
C3101 _32_/a_27_47# 0 0.175f
C3102 _11_ 0 0.261f
C3103 _50_/a_343_93# 0 0.172f
C3104 _50_/a_223_47# 0 0.141f
C3105 _50_/a_27_47# 0 0.259f
C3106 _07_ 0 0.285f
C3107 net13 0 0.382f
C3108 _33_/a_209_311# 0 0.143f
C3109 _33_/a_109_93# 0 0.158f
C3110 _08_ 0 0.128f
C3111 net11 0 0.717f
C3112 net12 0 0.517f
C3113 _34_/a_285_47# 0 0.0174f
C3114 _34_/a_47_47# 0 0.199f
C3115 _23_ 0 0.106f
C3116 p[9] 0 0.434f
C3117 input15/a_27_47# 0 0.208f
C3118 _35_/a_489_413# 0 0.0254f
C3119 _35_/a_226_47# 0 0.162f
C3120 _35_/a_76_199# 0 0.141f
C3121 _24_ 0 0.135f
C3122 _12_ 0 0.372f
C3123 _52_/a_250_297# 0 0.0278f
C3124 _52_/a_93_21# 0 0.151f
C3125 _10_ 0 0.629f
C3126 _36_/a_27_47# 0 0.175f
C3127 p[8] 0 0.725f
C3128 input14/a_27_47# 0 0.208f
C3129 _53_/a_29_53# 0 0.18f
C3130 _37_/a_27_47# 0 0.175f
C3131 p[7] 0 0.603f
C3132 input13/a_27_47# 0 0.208f
C3133 net18 0 0.201f
C3134 _25_ 0 0.184f
C3135 _54_/a_75_212# 0 0.21f
C3136 _38_/a_27_47# 0 0.175f
C3137 net19 0 0.171f
C3138 _22_ 0 0.215f
C3139 _14_ 0 0.219f
C3140 _15_ 0 0.333f
C3141 _55_/a_217_297# 0 0.00117f
C3142 _55_/a_80_21# 0 0.21f
C3143 p[6] 0 1.25f
C3144 input12/a_27_47# 0 0.208f
C3145 p[3] 0 3.15f
C3146 input9/a_75_212# 0 0.21f
C3147 _39_/a_285_47# 0 0.0174f
C3148 _39_/a_47_47# 0 0.199f
C3149 p[5] 0 0.927f
C3150 input11/a_27_47# 0 0.208f
C3151 p[2] 0 1.1f
C3152 input8/a_27_47# 0 0.208f
C3153 p[4] 0 1.77f
C3154 input10/a_27_47# 0 0.208f
C3155 net7 0 0.458f
C3156 p[1] 0 1.1f
C3157 input7/a_27_47# 0 0.208f
C3158 p[14] 0 0.547f
C3159 input6/a_27_47# 0 0.208f
C3160 net5 0 0.819f
C3161 p[13] 0 0.763f
C3162 input5/a_841_47# 0 0.0929f
C3163 input5/a_664_47# 0 0.13f
C3164 input5/a_558_47# 0 0.164f
C3165 input5/a_381_47# 0 0.11f
C3166 input5/a_62_47# 0 0.169f
C3167 p[12] 0 0.44f
C3168 input4/a_75_212# 0 0.21f
C3169 p[11] 0 0.522f
C3170 input3/a_27_47# 0 0.208f
C3171 net2 0 0.66f
C3172 p[10] 0 0.917f
C3173 input2/a_27_47# 0 0.208f
C3174 net1 0 0.338f
C3175 p[0] 0 1.46f
C3176 input1/a_75_212# 0 0.21f
C3177 b[3] 0 3.49f
C3178 output19/a_27_47# 0 0.543f
C3179 b[2] 0 0.429f
C3180 output18/a_27_47# 0 0.543f
C3181 b[1] 0 0.422f
C3182 net17 0 0.17f
C3183 output17/a_27_47# 0 0.543f
C3184 _41_/a_59_75# 0 0.177f
C3185 b[0] 0 0.788f
C3186 output16/a_27_47# 0 0.543f
C3187 _16_ 0 0.125f
C3188 _42_/a_209_311# 0 0.143f
C3189 _42_/a_109_93# 0 0.158f
C3190 _17_ 0 0.248f
C3191 _43_/a_193_413# 0 0.136f
C3192 _43_/a_27_47# 0 0.224f
C3193 _00_ 0 0.377f
C3194 net6 0 0.527f
C3195 net4 0 0.311f
C3196 _26_/a_29_53# 0 0.18f
C3197 _01_ 0 0.15f
C3198 net14 0 0.511f
C3199 net3 0 0.472f
C3200 net15 0 0.441f
C3201 _27_/a_27_297# 0 0.163f
C3202 _18_ 0 0.143f
C3203 _44_/a_250_297# 0 0.0278f
C3204 _44_/a_93_21# 0 0.151f
C3205 net16 0 0.218f
C3206 _09_ 0 0.14f
C3207 _13_ 0 0.13f
C3208 _45_/a_193_297# 0 0.0011f
C3209 _45_/a_109_297# 0 7.11e-19
C3210 _45_/a_27_47# 0 0.216f
C3211 _29_/a_29_53# 0 0.18f
C3212 _19_ 0 0.114f
C3213 _47_/a_299_297# 0 0.0348f
C3214 _47_/a_81_21# 0 0.147f
C3215 VPWR 0 40.6f
C3216 VGND 0 12.7f
C3217 _48_/a_27_47# 0 0.177f
C3218 _21_ 0 0.288f
C3219 _20_ 0 0.238f
C3220 _02_ 0 0.446f
C3221 _49_/a_201_297# 0 0.00345f
C3222 _49_/a_75_199# 0 0.205f
.ends

.subckt analog_therm
Xx1 x1/Vin x1/Vp x1/V1 x1/V2 x1/V3 x1/V4 x1/V5 x1/V6 x1/V7 x1/V8 x1/V10 x1/V11 x1/V12
+ x1/V13 x1/V14 x1/V15 x1/x28/m1_1594_n962# x1/x29/m1_1074_6# x1/Vp x1/x22/m1_451_n1105#
+ x1/x30/Vin x1/x29/m1_915_n714# x1/x28/m1_710_n388# x1/x28/m1_2498_n384# x1/x21/m1_400_n1066#
+ x1/x27/m1_724_n958# x1/x26/m1_532_n361# x1/x30/Vin x1/x31/m1_931_n929# x1/x25/m1_717_301#
+ x1/th10_0/m1_718_n418# x1/x30/Vin x1/x16/m1_1199_9# x1/x17/m1_522_n210# x1/x26/m1_773_n853#
+ x1/x17/li_1010_10# x1/x30/Vin x1/x16/m1_4146_502# VSUBS x1/x19/m1_836_n724# x1/x20/m1_528_n874#
+ x1/x23/m1_891_n977# x1/x23/m1_1725_85# x1/x30/Vin x1/x27/m1_546_n454# x1/Vp x1/x25/m1_509_303#
+ x1/Vp x1/Vp x1/Vp x1/Vp x1/x17/m1_782_n682# x1/V9 x1/x30/Vin x1/x30/Vin x1/x18/m1_960_n972#
+ x1/x18/m1_397_n357# VSUBS x1/x29/m1_1076_814# Analog
Xx2 x2/b[0] x2/b[2] x1/V12 x1/V13 x1/V14 x1/V15 x1/V3 x1/V6 x1/V9 x2/input3/a_27_47#
+ x2/_35_/a_226_47# x2/input4/a_75_212# x2/_50_/a_27_47# x2/_45_/a_465_47# x2/net7
+ x2/input13/a_27_47# x2/_45_/a_205_47# x2/_30_/a_215_297# x2/output19/a_27_47# x2/net19
+ x2/_45_/a_27_47# x2/input10/a_27_47# x2/_18_ x2/_10_ x2/_31_/a_285_47# x2/_31_/a_35_297#
+ x2/_50_/a_429_93# x2/_07_ x2/input7/a_27_47# x2/_04_ x2/output16/a_27_47# x2/input9/a_75_212#
+ x2/_30_/a_109_53# x2/_39_/a_129_47# x2/b[1] x2/_27_/a_27_297# x2/input1/a_75_212#
+ x2/_41_/a_59_75# x2/input5/a_62_47# x2/net3 x2/input14/a_27_47# x2/b[3] x2/_31_/a_285_297#
+ x2/_11_ x2/net2 x2/_47_/a_81_21# x2/_49_/a_208_47# x1/V1 x2/_09_ x2/net14 x2/_13_
+ x2/_34_/a_47_47# x2/_19_ x2/input11/a_27_47# x2/net12 x2/_34_/a_285_47# x2/_49_/a_75_199#
+ x2/net4 x2/_47_/a_384_47# x2/net8 x2/net6 x2/_17_ x2/input8/a_27_47# x2/_33_/a_209_311#
+ x2/_41_/a_145_75# x2/output17/a_27_47# x1/V8 x2/_01_ x2/_37_/a_27_47# x2/_38_/a_109_47#
+ x2/_47_/a_299_297# x2/_44_/a_93_21# x2/_44_/a_250_297# x1/V10 x2/net13 x2/_02_ x2/input15/a_27_47#
+ x2/_39_/a_47_47# x2/_43_/a_27_47# x1/V2 x2/_50_/a_223_47# x2/_50_/a_515_93# x2/input2/a_27_47#
+ x2/_38_/a_197_47# x2/_15_ x2/_50_/a_615_93# x2/_14_ x2/input12/a_27_47# x1/V4 x2/_20_
+ x2/net1 x2/_38_/a_27_47# x1/Vp x2/_34_/a_129_47# x2/net11 x2/_03_ x2/_06_ x2/_49_/a_315_47#
+ x2/net16 x2/net10 x2/output18/a_27_47# x2/_08_ x2/_16_ x2/_34_/a_377_297# x2/_12_
+ x2/net9 x2/_00_ x2/_05_ x1/V5 x2/input6/a_27_47# x2/_39_/a_285_47# x2/net17 x2/_31_/a_117_297#
+ VSUBS x2/_50_/a_343_93# x2/net5 x1/V11 x2/_39_/a_377_297# x2/net15 VSUBS x1/V7 therm
C0 x1/Vp x2/_31_/a_285_47# 2.02e-19
C1 x2/net16 x1/V13 2.61e-19
C2 x2/input10/a_27_47# x1/Vp 4.48e-20
C3 x1/Vp x2/_07_ 5.15e-19
C4 x1/x23/m1_891_n977# x1/Vp -2.74e-20
C5 x1/x28/m1_2498_n384# x1/V12 3.29e-19
C6 x2/net14 VSUBS 7.36e-21
C7 x1/Vp x1/x29/m1_1076_814# 0.00259f
C8 x1/x27/m1_724_n958# VSUBS 5.85e-20
C9 x1/x25/m1_717_301# VSUBS -0.0087f
C10 x2/output19/a_27_47# x1/V15 0.00109f
C11 x2/net15 x1/V15 1.08e-19
C12 x1/x23/m1_891_n977# x1/x27/m1_546_n454# -0.00212f
C13 x1/V3 x1/x17/li_1010_10# 0.0803f
C14 x1/x20/m1_528_n874# x1/Vp 1.25e-19
C15 x1/th10_0/m1_718_n418# VSUBS 0.00114f
C16 x2/b[1] x1/x17/li_1010_10# 5.1e-20
C17 x2/_01_ VSUBS 1.42e-32
C18 x1/x27/m1_546_n454# x1/x29/m1_1076_814# -2.28e-19
C19 x1/V11 x1/x25/m1_717_301# 0.0286f
C20 x1/Vp x2/_50_/a_343_93# 1.47e-20
C21 x1/Vp x2/b[3] 0.966f
C22 x2/b[1] x1/V1 -0.0017f
C23 x1/Vp x1/x26/m1_773_n853# 0.0055f
C24 x1/x22/m1_451_n1105# x2/b[3] 0.00378f
C25 x2/_30_/a_109_53# x1/x16/m1_4146_502# 1.22e-19
C26 x1/V4 x1/x31/m1_931_n929# -0.0169f
C27 x1/x28/m1_2498_n384# VSUBS 6.56e-19
C28 x2/output18/a_27_47# x1/x30/Vin 9.47e-21
C29 x2/_39_/a_47_47# x1/Vp 0.00244f
C30 x2/_19_ x1/Vp 4.43e-19
C31 x1/x29/m1_915_n714# VSUBS 0.0156f
C32 x1/x16/m1_1199_9# x1/V4 0.00202f
C33 x2/b[1] x2/_34_/a_47_47# -3.19e-20
C34 x1/x20/m1_528_n874# x1/V7 0.00258f
C35 x2/_38_/a_109_47# x1/Vp 1.11e-19
C36 x1/V15 x1/x30/Vin 0.00517f
C37 x2/input15/a_27_47# VSUBS 1.28e-19
C38 x1/Vp x2/net13 1.18e-19
C39 x2/b[1] x1/V3 -9.6e-20
C40 x1/Vp x2/net12 0.00206f
C41 x2/_47_/a_299_297# x1/Vp 0.00107f
C42 x2/_38_/a_197_47# x1/Vp 9.52e-20
C43 x1/x29/m1_1074_6# x1/V15 2.45e-19
C44 VSUBS x2/net2 0.00474f
C45 x2/b[2] x2/b[1] -7.17e-19
C46 x2/_31_/a_35_297# x1/Vp 0.00138f
C47 x1/V9 x1/x30/Vin 0.00435f
C48 x2/input1/a_75_212# x1/x28/m1_710_n388# 9.92e-21
C49 x2/net6 x2/net2 5.55e-35
C50 x1/x21/m1_400_n1066# x1/x30/Vin -5.68e-32
C51 x1/x19/m1_836_n724# x1/V7 0.0116f
C52 x1/x16/m1_4146_502# x1/V4 0.214f
C53 x1/x29/m1_1074_6# x1/V9 2.24e-21
C54 x1/x28/m1_710_n388# x1/V1 7.62e-20
C55 x1/V14 x2/b[3] 0.073f
C56 x2/b[1] x2/_34_/a_377_297# -2.08e-20
C57 x2/output19/a_27_47# x1/Vp 2.83e-19
C58 x2/net15 x1/Vp 5.92e-20
C59 x2/net16 x1/Vp 1.23e-19
C60 x2/_37_/a_27_47# x1/V15 4.31e-21
C61 x1/V13 VSUBS 0.0287f
C62 x1/x17/m1_522_n210# x1/V2 3.71e-19
C63 x2/input4/a_75_212# x1/V15 4.55e-20
C64 x2/input12/a_27_47# x1/x17/li_1010_10# 3.04e-20
C65 x2/_30_/a_109_53# x2/b[3] -3.47e-36
C66 x2/b[1] x1/x28/m1_710_n388# 6.49e-20
C67 x2/input7/a_27_47# x1/Vp 0.00549f
C68 x1/x16/m1_4146_502# x2/b[3] 2.81e-19
C69 x1/V10 x1/x29/m1_1076_814# 5.18e-19
C70 x1/x21/m1_400_n1066# x1/V8 1.6e-20
C71 x2/input11/a_27_47# x1/Vp 4.48e-20
C72 x1/V15 VSUBS 0.109f
C73 x2/_04_ x1/Vp 1.98e-19
C74 x1/x25/m1_717_301# x1/V1 0.00428f
C75 x1/Vp x1/x30/Vin 1.85f
C76 x1/x22/m1_451_n1105# x1/x30/Vin -3.71e-20
C77 x2/net6 x1/V15 2.29e-20
C78 x1/V10 x2/b[3] -1.42e-20
C79 x2/net5 x1/x28/m1_710_n388# 6.72e-22
C80 x2/_31_/a_117_297# x1/Vp 5.01e-19
C81 x1/V9 VSUBS 0.0728f
C82 x1/Vp x1/V2 0.37f
C83 x1/x17/m1_782_n682# x1/V7 1.95e-20
C84 x2/_37_/a_27_47# x2/net3 2.84e-32
C85 x2/b[0] x1/x30/Vin 0.0688f
C86 x2/_14_ x1/V15 1.2e-20
C87 x2/b[3] x1/V4 -0.00234f
C88 x2/net1 x1/V3 -1.73e-20
C89 x1/x27/m1_724_n958# x2/b[1] 8.7e-21
C90 x2/_45_/a_465_47# x1/Vp 6.63e-20
C91 x1/V7 x1/x30/Vin 0.069f
C92 x1/Vp x2/net10 0.00102f
C93 x2/_09_ x1/Vp 7.15e-20
C94 x1/Vp x1/V8 0.132f
C95 x2/input4/a_75_212# x1/Vp 0.00341f
C96 x1/V12 x1/Vp 0.0523f
C97 x2/net3 VSUBS 2.04e-20
C98 x1/x30/Vin x1/x31/m1_931_n929# 0.00651f
C99 x1/x22/m1_451_n1105# x1/V8 0.00976f
C100 x2/_41_/a_59_75# VSUBS 9.12e-20
C101 x2/_15_ x1/Vp 0.00491f
C102 x2/_06_ x2/net10 2.84e-32
C103 x1/x16/m1_1199_9# x1/x30/Vin -0.0164f
C104 x2/_34_/a_285_47# x1/Vp 5.81e-19
C105 x2/_17_ x2/net2 -2.84e-32
C106 x1/x20/m1_528_n874# x2/b[3] 0.00287f
C107 x2/_10_ x1/V15 5.92e-20
C108 x2/_16_ VSUBS 3.55e-33
C109 x2/output16/a_27_47# x1/V13 6.08e-20
C110 x2/_49_/a_315_47# x1/Vp 7.63e-21
C111 x1/x25/m1_509_303# x1/Vp 0.0375f
C112 x2/_47_/a_384_47# x1/Vp 6.21e-20
C113 x2/input9/a_75_212# x1/V3 -2.54e-21
C114 x2/output17/a_27_47# VSUBS 2e-20
C115 x1/x16/m1_1199_9# x1/V2 1.55e-19
C116 x2/net11 x1/x30/Vin 4.48e-19
C117 x1/Vp VSUBS 1.99f
C118 x1/V10 x2/net15 6.08e-21
C119 x1/Vp x2/net8 0.00652f
C120 x1/V15 x2/input6/a_27_47# 2.43e-19
C121 x1/V7 x1/V8 0.253f
C122 x1/x22/m1_451_n1105# VSUBS 3.63e-21
C123 x1/Vp x1/V6 0.155f
C124 x1/V11 x1/Vp 0.177f
C125 x1/x26/m1_532_n361# x1/Vp 0.0363f
C126 x1/x27/m1_546_n454# VSUBS 0.00694f
C127 x2/net1 x1/x28/m1_710_n388# 1.2e-20
C128 x2/net6 x1/Vp 0.00481f
C129 x2/_31_/a_285_297# x1/Vp 4.79e-19
C130 x2/_06_ VSUBS 1.11e-19
C131 x2/_39_/a_377_297# x1/Vp 3.97e-19
C132 x1/th10_0/m1_718_n418# x1/x28/m1_710_n388# 3.92e-19
C133 x1/Vp x2/_49_/a_208_47# 2.29e-20
C134 x2/net7 x1/Vp 0.0069f
C135 x2/b[0] VSUBS 0.0511f
C136 x1/x21/m1_400_n1066# x1/V5 6.29e-19
C137 x1/x16/m1_4146_502# x1/x30/Vin -0.0056f
C138 x2/_30_/a_109_53# x1/V2 1.65e-20
C139 x1/V12 x1/V14 0.00499f
C140 x1/V7 VSUBS 0.36f
C141 x2/_08_ x1/Vp 6.6e-19
C142 x1/V7 x1/V6 -0.0155f
C143 x1/V15 x2/_17_ 4.4e-22
C144 x1/V10 x1/x30/Vin 0.00287f
C145 x1/x16/m1_4146_502# x1/V2 0.126f
C146 x1/Vp x2/_33_/a_209_311# 1.21e-21
C147 x1/x25/m1_509_303# x1/x31/m1_931_n929# -0.0022f
C148 x1/x17/m1_782_n682# x1/V4 0.0101f
C149 x1/Vp x2/_13_ 0.00257f
C150 x2/net15 x1/x29/m1_1076_814# 4.68e-20
C151 x1/x18/m1_397_n357# x1/Vp 2.29e-19
C152 x1/x31/m1_931_n929# VSUBS 0.114f
C153 x1/Vp x2/input8/a_27_47# 0.00419f
C154 x1/x16/m1_1199_9# VSUBS 0.0629f
C155 x1/V14 VSUBS 0.021f
C156 x1/x30/Vin x1/V4 0.632f
C157 x2/net19 x1/V15 2.1e-19
C158 x1/x16/m1_4146_502# x2/net10 4.87e-21
C159 x1/V11 x1/x16/m1_1199_9# 1.51e-19
C160 x2/_10_ x1/Vp 0.00418f
C161 x1/x28/m1_1594_n962# x1/Vp 8.18e-20
C162 x1/V11 x1/V14 0.0919f
C163 x1/x28/m1_710_n388# x2/net2 1.86e-20
C164 x2/input13/a_27_47# x1/Vp 3.64e-19
C165 x2/input10/a_27_47# x1/x30/Vin 0.00121f
C166 x2/_35_/a_226_47# x1/Vp 5.68e-32
C167 x1/Vp x1/V5 0.229f
C168 x1/V2 x1/V4 0.0745f
C169 x2/_12_ x1/V13 7.61e-22
C170 x1/x22/m1_451_n1105# x1/V5 0.0218f
C171 x2/net11 x1/V6 -0.00685f
C172 x1/Vp x2/input6/a_27_47# 2.52e-20
C173 x1/x17/m1_782_n682# x2/b[3] 2.4e-20
C174 x2/_37_/a_27_47# x1/V10 2.05e-20
C175 x1/V10 x1/V12 0.0056f
C176 x2/_43_/a_27_47# VSUBS 2.84e-32
C177 x2/net5 x1/V15 7.26e-21
C178 x1/x16/m1_4146_502# VSUBS 0.0251f
C179 x1/V3 x1/x17/m1_522_n210# 0.00261f
C180 x1/x30/Vin x2/b[3] 0.366f
C181 x2/output16/a_27_47# x1/x27/m1_546_n454# 1.15e-19
C182 x1/x30/Vin x1/x26/m1_773_n853# 0.0251f
C183 x2/_12_ x1/V15 5.5e-21
C184 x2/_47_/a_81_21# VSUBS 2.06e-20
C185 x1/V5 x1/V7 0.00522f
C186 x2/input1/a_75_212# x1/Vp 0.00577f
C187 x1/Vp x2/_03_ 3.58e-20
C188 x1/V10 VSUBS 0.0168f
C189 x1/Vp x1/V1 0.577f
C190 x2/b[3] x1/V2 -0.00101f
C191 x1/Vp x2/_17_ 6.82e-19
C192 x1/x19/m1_836_n724# x1/x30/Vin -2.9e-20
C193 x2/net6 x1/V10 -5.68e-32
C194 x2/_37_/a_27_47# x1/x29/m1_1076_814# 8.05e-20
C195 x1/x20/m1_528_n874# x1/V8 -6.58e-19
C196 x1/V4 VSUBS 0.856f
C197 x2/net13 x1/x30/Vin 6.02e-19
C198 x2/_00_ VSUBS 1.42e-31
C199 x1/x30/Vin x2/net12 6.06e-19
C200 x1/x28/m1_2498_n384# x2/net2 2.31e-19
C201 x1/Vp x2/_34_/a_47_47# 0.00222f
C202 x1/x17/li_1010_10# x1/V7 9.05e-20
C203 x1/V8 x2/b[3] 1.78e-33
C204 x1/x16/m1_4146_502# x1/x18/m1_397_n357# -3.84e-19
C205 x1/V12 x2/b[3] 6.93e-19
C206 x1/V3 x1/Vp 0.776f
C207 x2/b[1] x1/Vp 0.116f
C208 x2/_20_ x1/Vp 4.47e-19
C209 x1/x22/m1_451_n1105# x1/V3 0.00381f
C210 x1/x18/m1_960_n972# x1/Vp 0.001f
C211 x2/b[2] x1/Vp 0.0143f
C212 x1/x29/m1_1076_814# VSUBS 0.0247f
C213 x1/x20/m1_528_n874# VSUBS 4.22e-19
C214 x2/b[1] x2/_06_ -4.61e-19
C215 x1/V1 x1/x31/m1_931_n929# 5.68e-32
C216 x1/x19/m1_836_n724# x1/V8 -0.00357f
C217 x1/x25/m1_509_303# x2/b[3] 5.1e-21
C218 x2/net6 x1/x29/m1_1076_814# 6.33e-20
C219 x1/x20/m1_528_n874# x1/V6 0.00476f
C220 x2/net14 x1/V15 2.63e-20
C221 x2/_50_/a_429_93# x1/Vp 5.73e-20
C222 x1/x16/m1_1199_9# x1/V1 0.0151f
C223 x2/_50_/a_343_93# VSUBS -7.11e-33
C224 x2/b[3] VSUBS 0.153f
C225 x1/V14 x1/V1 -1.81e-19
C226 x2/net5 x1/Vp 0.00362f
C227 x2/output19/a_27_47# x1/x29/m1_1074_6# 1.14e-20
C228 x2/_34_/a_377_297# x1/Vp 1.63e-19
C229 x1/x18/m1_397_n357# x1/V4 9.29e-19
C230 x2/b[3] x1/V6 -0.00218f
C231 x1/V11 x2/b[3] 0.00987f
C232 x2/_12_ x1/Vp 0.00229f
C233 x1/Vp x2/net9 1.13e-19
C234 x1/V3 x1/V7 1.13e-19
C235 x2/net6 x2/b[3] -2.22e-34
C236 x1/x29/m1_915_n714# x1/V15 9.36e-19
C237 x2/input11/a_27_47# x1/x30/Vin 0.00123f
C238 x1/V12 x2/input3/a_27_47# 2.84e-32
C239 x1/x28/m1_710_n388# x1/Vp 0.0084f
C240 x1/Vp x2/_41_/a_145_75# 3.55e-19
C241 x1/x17/m1_782_n682# x1/V2 1.63e-21
C242 x1/x16/m1_4146_502# x2/_03_ 1.59e-21
C243 x2/input7/a_27_47# x1/V2 -1.2e-20
C244 x1/x16/m1_4146_502# x1/V1 0.00499f
C245 x2/input15/a_27_47# x1/V15 1.72e-19
C246 x1/x29/m1_915_n714# x1/V9 9.46e-20
C247 x1/Vp x2/net17 0.00167f
C248 x2/_31_/a_35_297# VSUBS 9.34e-21
C249 x1/x30/Vin x1/V2 0.269f
C250 x2/b[1] x2/net11 -1.86e-19
C251 x1/V15 x2/net2 3.61e-20
C252 x1/x17/m1_782_n682# x1/V8 3.08e-20
C253 x2/input12/a_27_47# x1/Vp 4.48e-20
C254 x1/x17/li_1010_10# x1/V4 0.0308f
C255 x1/x20/m1_528_n874# x1/V5 0.0107f
C256 x2/output19/a_27_47# VSUBS 7.4e-19
C257 x2/input6/a_27_47# x1/x29/m1_1076_814# 1.12e-20
C258 x2/net15 VSUBS 5.06e-20
C259 x2/_50_/a_515_93# x1/Vp 9.87e-20
C260 x1/x30/Vin x2/net10 6.01e-19
C261 x2/net16 VSUBS 2.99e-20
C262 x1/x16/m1_4146_502# x1/V3 0.019f
C263 x2/input10/a_27_47# x1/x17/li_1010_10# 3.42e-20
C264 x1/V5 x2/b[3] -6.14e-20
C265 x2/b[1] x1/x16/m1_4146_502# 1.41e-19
C266 x2/net14 x1/Vp 6.13e-20
C267 x1/V1 x1/V4 -0.0454f
C268 x2/net1 x1/Vp 0.00672f
C269 x1/x30/Vin x1/V8 0.00885f
C270 x1/x25/m1_717_301# x1/Vp 0.0206f
C271 x1/V12 x1/x30/Vin 5.32e-20
C272 x2/net19 x1/V10 1.63e-20
C273 x1/th10_0/m1_718_n418# x1/Vp 8.17e-19
C274 x2/_01_ x1/Vp 6.26e-20
C275 x1/V13 x1/V15 4.14e-19
C276 x1/x28/m1_710_n388# x1/V14 0.0787f
C277 x1/x17/m1_782_n682# VSUBS 2.56e-20
C278 x1/x19/m1_836_n724# x1/V5 0.0407f
C279 x2/input7/a_27_47# VSUBS 2.73e-20
C280 x1/x27/m1_724_n958# x2/b[0] 0.0054f
C281 x1/x28/m1_2498_n384# x1/Vp 3.74e-19
C282 x1/x25/m1_509_303# x1/x30/Vin 0.005f
C283 x1/x23/m1_1725_85# x1/V9 0.0382f
C284 x2/input14/a_27_47# x2/net2 2.22e-34
C285 x1/V13 x1/V9 0.183f
C286 x1/V11 x2/input7/a_27_47# 2.22e-34
C287 x1/x29/m1_915_n714# x1/Vp 1.59e-19
C288 x1/x17/li_1010_10# x2/b[3] 6.8e-20
C289 x1/x30/Vin VSUBS 0.684f
C290 x1/x16/m1_4146_502# x2/net9 9.47e-21
C291 x1/V3 x1/V4 -0.00444f
C292 x2/net8 x1/x30/Vin 1.77e-20
C293 x1/x30/Vin x1/V6 0.339f
C294 x1/V11 x1/x30/Vin 6.89e-20
C295 x1/x26/m1_532_n361# x1/x30/Vin 3.98e-20
C296 x1/x18/m1_960_n972# x1/V4 6.61e-19
C297 x2/input9/a_75_212# x1/Vp 0.00113f
C298 x1/x29/m1_1074_6# VSUBS 3.62e-19
C299 x1/V1 x2/b[3] -0.00159f
C300 x2/_05_ x1/Vp 2.87e-19
C301 x1/Vp x2/_02_ 9.59e-20
C302 x2/input15/a_27_47# x1/Vp 2.4e-20
C303 x2/_44_/a_93_21# VSUBS -5.68e-32
C304 x1/V2 VSUBS 0.0461f
C305 x1/V15 x1/V9 0.353f
C306 x1/Vp x2/net2 0.00334f
C307 x2/b[1] x1/x20/m1_528_n874# 7.29e-21
C308 x2/_50_/a_615_93# x1/Vp 1.07e-19
C309 x1/V10 x1/x28/m1_710_n388# -6.8e-21
C310 x1/V3 x2/b[3] -0.00226f
C311 x1/V8 VSUBS -0.0221f
C312 x2/b[1] x2/b[3] -6.38e-19
C313 x2/_37_/a_27_47# VSUBS 1.66e-21
C314 x2/input4/a_75_212# VSUBS 7.71e-20
C315 x1/V12 VSUBS 0.0114f
C316 x1/x28/m1_2498_n384# x1/V14 0.0267f
C317 x1/x30/Vin x2/input8/a_27_47# 3.42e-19
C318 x2/input14/a_27_47# x1/V15 3.98e-20
C319 x2/_34_/a_129_47# x1/Vp 1.22e-19
C320 x1/Vp x2/_18_ 9.91e-20
C321 x1/V13 x1/Vp 0.0257f
C322 x2/net3 x1/V15 1.07e-19
C323 x2/_27_/a_27_297# x1/Vp 2.53e-19
C324 x2/_41_/a_59_75# x1/V15 5.91e-20
C325 x1/x27/m1_546_n454# x1/x23/m1_1725_85# -2.91e-19
C326 x1/x28/m1_1594_n962# x1/x30/Vin 0.0193f
C327 x1/x27/m1_546_n454# x1/V13 -5.17e-20
C328 x1/x25/m1_509_303# VSUBS -0.00786f
C329 x2/input13/a_27_47# x1/x30/Vin 0.00122f
C330 x2/_16_ x1/V15 2.48e-21
C331 x1/V5 x1/x30/Vin 0.121f
C332 x1/x25/m1_509_303# x1/V11 0.00995f
C333 x2/net8 VSUBS 9.41e-20
C334 x1/V13 x2/b[0] 4.93e-19
C335 x2/b[1] x2/net12 -3.49e-20
C336 x1/V6 VSUBS 0.00382f
C337 x1/V11 VSUBS 0.681f
C338 x2/net14 x1/V10 2.16e-19
C339 x2/net6 VSUBS 8.38e-21
C340 x1/Vp x1/V15 0.0232f
C341 x1/V10 x1/th10_0/m1_718_n418# 0.00288f
C342 x2/net7 VSUBS 3.18e-19
C343 x1/x27/m1_546_n454# x1/V15 -9.98e-19
C344 x2/output16/a_27_47# x1/x30/Vin 5.02e-19
C345 x1/V13 x2/_38_/a_27_47# 4.09e-20
C346 x1/x28/m1_710_n388# x2/b[3] 0.0129f
C347 x1/V15 x2/_06_ 6.92e-20
C348 x1/V11 x2/net7 2.22e-34
C349 x2/_14_ VSUBS -1.14e-31
C350 x1/Vp x1/V9 0.317f
C351 x1/x25/m1_717_301# x1/V4 -9.85e-19
C352 x2/input9/a_75_212# x1/x16/m1_4146_502# 6.09e-20
C353 x1/x29/m1_915_n714# x1/V10 4.86e-19
C354 x2/_19_ x1/x28/m1_710_n388# 2.44e-20
C355 x1/x27/m1_546_n454# x1/V9 0.208f
C356 x1/V1 x1/x30/Vin 0.166f
C357 x1/V5 x1/V8 0.0686f
C358 x1/x17/li_1010_10# x1/V2 0.00198f
C359 x1/x18/m1_397_n357# VSUBS 0.00233f
C360 x2/input8/a_27_47# VSUBS 6.94e-20
C361 x1/x17/m1_782_n682# x1/V3 0.0115f
C362 x2/b[1] x1/x17/m1_782_n682# 1.85e-20
C363 x2/net3 x1/Vp 5.92e-20
C364 x1/Vp x2/_39_/a_285_47# 6.21e-19
C365 x2/_10_ VSUBS 8.77e-20
C366 x1/V11 x1/Vin 3.64e-19
C367 x1/V10 x2/net2 5.29e-19
C368 x2/_41_/a_59_75# x1/Vp 0.00259f
C369 x1/Vp x2/_49_/a_75_199# 2.53e-19
C370 x2/input13/a_27_47# VSUBS 3.74e-21
C371 x1/x21/m1_400_n1066# x1/V7 0.00413f
C372 x1/V5 VSUBS 0.29f
C373 x1/x17/li_1010_10# x1/V8 2.35e-19
C374 x1/V3 x1/x30/Vin 0.423f
C375 x2/b[1] x1/x30/Vin 0.143f
C376 x1/Vp x2/net4 0.00699f
C377 x1/V5 x1/V6 4.11e-19
C378 x2/input6/a_27_47# VSUBS 1.75e-19
C379 x1/x18/m1_960_n972# x1/x30/Vin 1.28e-21
C380 x2/b[2] x1/x30/Vin 0.0471f
C381 x2/output17/a_27_47# x1/Vp 0.00644f
C382 x2/net6 x2/input6/a_27_47# 4.26e-32
C383 x1/V3 x1/V2 0.0548f
C384 x1/x28/m1_2498_n384# x2/b[3] 0.0373f
C385 x2/b[1] x1/V2 -2.18e-20
C386 x2/output16/a_27_47# VSUBS 3.5e-20
C387 x2/_30_/a_215_297# x1/Vp 1.17e-20
C388 x1/x27/m1_546_n454# x1/Vp 0.00106f
C389 x2/input15/a_27_47# x1/x29/m1_1076_814# 2.66e-20
C390 x1/x17/li_1010_10# VSUBS 0.00635f
C391 x1/Vp x2/_06_ 0.00399f
C392 x1/x25/m1_509_303# x1/V1 0.00256f
C393 x2/input1/a_75_212# VSUBS 5.9e-20
C394 x1/x29/m1_1076_814# x2/net2 5.25e-20
C395 x2/b[0] x1/Vp 0.0311f
C396 x2/b[1] x2/net10 -1.03e-20
C397 x2/_45_/a_27_47# x1/Vp 8.43e-19
C398 x1/V1 VSUBS 0.474f
C399 x1/Vp x2/_50_/a_27_47# 2.02e-19
C400 x1/V11 x2/input1/a_75_212# -1.33e-33
C401 x2/_47_/a_81_21# x1/V15 1.32e-21
C402 x1/V3 x1/V8 3.88e-19
C403 x2/_17_ VSUBS 1.83e-20
C404 x1/x27/m1_546_n454# x2/b[0] 0.00421f
C405 x1/V11 x1/V1 0.00263f
C406 x1/Vp x1/V7 0.0345f
C407 x1/V10 x1/V15 0.0116f
C408 x1/x22/m1_451_n1105# x1/V7 0.00397f
C409 x1/x28/m1_710_n388# x1/x30/Vin 0.0013f
C410 x2/_38_/a_27_47# x1/Vp 2.55e-19
C411 x2/net19 VSUBS 4.66e-20
C412 x1/Vp x1/x31/m1_931_n929# 0.0155f
C413 x1/V13 x1/x29/m1_1076_814# 3.47e-19
C414 x2/output17/a_27_47# x1/V14 9.62e-21
C415 x1/V10 x1/V9 0.00767f
C416 x1/x16/m1_1199_9# x1/Vp 0.0108f
C417 x1/V3 VSUBS 0.0756f
C418 x1/V14 x1/Vp 0.0723f
C419 x2/b[1] VSUBS 0.101f
C420 x1/V3 x2/net8 -1.25e-19
C421 x2/_20_ VSUBS -5.68e-32
C422 x1/x18/m1_960_n972# VSUBS 0.00319f
C423 x1/V11 x2/b[1] -5.92e-19
C424 VSUBS x2/_44_/a_250_297# -2.22e-34
C425 x2/b[2] VSUBS -1.79e-20
C426 x2/input12/a_27_47# x1/x30/Vin 0.00124f
C427 x2/net11 x1/Vp 0.0142f
C428 x2/output19/a_27_47# x1/x29/m1_915_n714# 2.24e-20
C429 x1/x18/m1_397_n357# x1/V1 2.1e-19
C430 x2/_39_/a_129_47# x1/Vp 6.96e-20
C431 x1/V15 x1/x29/m1_1076_814# 1.1e-19
C432 x2/_45_/a_205_47# x1/Vp 1.27e-20
C433 x2/_11_ x1/Vp 8.15e-19
C434 x1/x17/m1_522_n210# x1/V4 0.0102f
C435 x2/_30_/a_109_53# x1/Vp 1.26e-19
C436 x1/x28/m1_710_n388# x2/input5/a_62_47# 2.7e-20
C437 x1/V10 x2/input14/a_27_47# 3.18e-19
C438 x2/net5 VSUBS 6.84e-20
C439 x1/x17/li_1010_10# x1/V5 3.68e-20
C440 x1/x25/m1_717_301# x1/x30/Vin 0.0149f
C441 x2/net11 x2/_06_ 7.11e-33
C442 x1/V12 x1/x28/m1_710_n388# 8.88e-34
C443 x1/V10 x2/net3 0.00147f
C444 x2/_12_ VSUBS 2.35e-20
C445 x1/x23/m1_891_n977# x1/V9 0.028f
C446 x1/V15 x2/b[3] 3.63e-19
C447 x2/input2/a_27_47# x1/Vp 0.00193f
C448 x1/V9 x1/x29/m1_1076_814# 0.0223f
C449 x1/x16/m1_4146_502# x1/Vp 1.62e-19
C450 x2/_08_ x2/b[1] -2.59e-20
C451 x1/Vp x2/_50_/a_223_47# 9.53e-20
C452 x2/_47_/a_81_21# x1/Vp 6.37e-19
C453 x2/_30_/a_215_297# x1/x16/m1_4146_502# 9.48e-22
C454 x1/V3 x2/input8/a_27_47# -7.11e-21
C455 x1/x16/m1_1199_9# x1/V14 -0.00147f
C456 x1/V10 x1/Vp 0.0237f
C457 x1/x28/m1_710_n388# VSUBS 0.00968f
C458 x1/V11 x1/x28/m1_710_n388# 0.0173f
C459 x2/input13/a_27_47# x1/V3 1.73e-36
C460 x2/net3 x1/x29/m1_1076_814# 8.2e-21
C461 x1/V3 x1/V5 -5.19e-19
C462 x1/Vp x1/V4 0.477f
C463 x2/b[1] x1/V5 -6.14e-20
C464 x2/_04_ 0 0.338f
C465 x2/net9 0 0.306f
C466 x2/_03_ 0 0.36f
C467 x2/net10 0 0.412f
C468 x2/_30_/a_109_53# 0 0.159f
C469 x2/_30_/a_215_297# 0 0.142f
C470 x2/_05_ 0 0.152f
C471 x2/net8 0 0.384f
C472 x2/_31_/a_285_297# 0 0.00137f
C473 x2/_31_/a_35_297# 0 0.255f
C474 x2/_06_ 0 0.804f
C475 x2/_32_/a_27_47# 0 0.175f
C476 x2/_11_ 0 0.261f
C477 x2/_50_/a_343_93# 0 0.172f
C478 x2/_50_/a_223_47# 0 0.141f
C479 x2/_50_/a_27_47# 0 0.259f
C480 x2/_07_ 0 0.285f
C481 x2/net13 0 0.382f
C482 x2/_33_/a_209_311# 0 0.143f
C483 x2/_33_/a_109_93# 0 0.158f
C484 x2/_08_ 0 0.128f
C485 x2/net11 0 0.717f
C486 x2/net12 0 0.517f
C487 x2/_34_/a_285_47# 0 0.0174f
C488 x2/_34_/a_47_47# 0 0.199f
C489 x2/_23_ 0 0.106f
C490 x2/input15/a_27_47# 0 0.208f
C491 x2/_35_/a_489_413# 0 0.0254f
C492 x2/_35_/a_226_47# 0 0.162f
C493 x2/_35_/a_76_199# 0 0.141f
C494 x2/_24_ 0 0.135f
C495 x2/_12_ 0 0.372f
C496 x2/_52_/a_250_297# 0 0.0278f
C497 x2/_52_/a_93_21# 0 0.151f
C498 x2/_10_ 0 0.629f
C499 x2/_36_/a_27_47# 0 0.175f
C500 x2/input14/a_27_47# 0 0.208f
C501 x2/_53_/a_29_53# 0 0.18f
C502 x2/_37_/a_27_47# 0 0.175f
C503 x2/input13/a_27_47# 0 0.208f
C504 x2/net18 0 0.201f
C505 x2/_25_ 0 0.184f
C506 x2/_54_/a_75_212# 0 0.21f
C507 x2/_38_/a_27_47# 0 0.175f
C508 x2/net19 0 0.171f
C509 x2/_22_ 0 0.215f
C510 x2/_14_ 0 0.219f
C511 x2/_15_ 0 0.333f
C512 x2/_55_/a_217_297# 0 0.00117f
C513 x2/_55_/a_80_21# 0 0.21f
C514 x2/input12/a_27_47# 0 0.208f
C515 x2/input9/a_75_212# 0 0.21f
C516 x2/_39_/a_285_47# 0 0.0174f
C517 x2/_39_/a_47_47# 0 0.199f
C518 x2/input11/a_27_47# 0 0.208f
C519 x2/input8/a_27_47# 0 0.208f
C520 x2/input10/a_27_47# 0 0.208f
C521 x2/net7 0 0.458f
C522 x2/input7/a_27_47# 0 0.208f
C523 x2/input6/a_27_47# 0 0.208f
C524 x2/net5 0 0.819f
C525 x2/input5/a_841_47# 0 0.0929f
C526 x2/input5/a_664_47# 0 0.13f
C527 x2/input5/a_558_47# 0 0.164f
C528 x2/input5/a_381_47# 0 0.11f
C529 x2/input5/a_62_47# 0 0.169f
C530 x2/input4/a_75_212# 0 0.21f
C531 x2/input3/a_27_47# 0 0.208f
C532 x2/net2 0 0.66f
C533 x2/input2/a_27_47# 0 0.208f
C534 x2/net1 0 0.338f
C535 x2/input1/a_75_212# 0 0.21f
C536 x2/b[3] 0 3.49f
C537 x2/output19/a_27_47# 0 0.543f
C538 x2/b[2] 0 0.429f
C539 x2/output18/a_27_47# 0 0.543f
C540 x2/b[1] 0 0.422f
C541 x2/net17 0 0.17f
C542 x2/output17/a_27_47# 0 0.543f
C543 x2/_41_/a_59_75# 0 0.177f
C544 x2/b[0] 0 0.788f
C545 x2/output16/a_27_47# 0 0.543f
C546 x2/_16_ 0 0.125f
C547 x2/_42_/a_209_311# 0 0.143f
C548 x2/_42_/a_109_93# 0 0.158f
C549 x2/_17_ 0 0.248f
C550 x2/_43_/a_193_413# 0 0.136f
C551 x2/_43_/a_27_47# 0 0.224f
C552 x2/_00_ 0 0.377f
C553 x2/net6 0 0.527f
C554 x2/net4 0 0.311f
C555 x2/_26_/a_29_53# 0 0.18f
C556 x2/_01_ 0 0.15f
C557 x2/net14 0 0.511f
C558 x2/net3 0 0.472f
C559 x2/net15 0 0.441f
C560 x2/_27_/a_27_297# 0 0.163f
C561 x2/_18_ 0 0.143f
C562 x2/_44_/a_250_297# 0 0.0278f
C563 x2/_44_/a_93_21# 0 0.151f
C564 x2/net16 0 0.218f
C565 x2/_09_ 0 0.14f
C566 x2/_13_ 0 0.13f
C567 x2/_45_/a_193_297# 0 0.0011f
C568 x2/_45_/a_109_297# 0 7.11e-19
C569 x2/_45_/a_27_47# 0 0.216f
C570 x2/_29_/a_29_53# 0 0.18f
C571 x2/_19_ 0 0.114f
C572 x2/_47_/a_299_297# 0 0.0348f
C573 x2/_47_/a_81_21# 0 0.147f
C574 x1/Vp 0 0.131p
C575 VSUBS 0 25.4f
C576 x2/_48_/a_27_47# 0 0.177f
C577 x2/_21_ 0 0.288f
C578 x2/_20_ 0 0.238f
C579 x2/_02_ 0 0.446f
C580 x2/_49_/a_201_297# 0 0.00345f
C581 x2/_49_/a_75_199# 0 0.205f
C582 x1/Vin 0 0.181f
C583 x1/V5 0 1.61f
C584 x1/x19/m1_836_n724# 0 1.02f
C585 x1/V4 0 2.79f
C586 x1/x18/m1_960_n972# 0 0.53f
C587 x1/x18/m1_397_n357# 0 0.189f
C588 x1/x29/m1_4024_602# 0 0.411f
C589 x1/V15 0 2.36f
C590 x1/x29/m1_1076_814# 0 5.99f
C591 x1/x29/m1_1074_6# 0 0.643f
C592 x1/x29/m1_915_n714# 0 0.787f
C593 x1/V3 0 1.16f
C594 x1/x17/m1_782_n682# 0 1.41f
C595 x1/x17/m1_522_n210# 0 0.24f
C596 x1/x17/li_1010_10# 0 2.8f
C597 x1/V14 0 1.48f
C598 x1/x28/m1_710_n388# 0 3.52f
C599 x1/x28/m1_2498_n384# 0 0.297f
C600 x1/x28/m1_1594_n962# 0 0.292f
C601 x1/x16/m1_4146_502# 0 7.92f
C602 x1/V2 0 1.24f
C603 x1/x16/m1_1199_9# 0 0.377f
C604 x1/V13 0 1.05f
C605 x1/x27/m1_546_n454# 0 1.54f
C606 x1/x27/m1_724_n958# 0 0.188f
C607 x1/x25/m1_509_303# 0 0.622f
C608 x1/V11 0 1.33f
C609 x1/x25/m1_717_301# 0 0.231f
C610 x1/x26/m1_532_n361# 0 0.839f
C611 x1/V12 0 1.43f
C612 x1/x26/m1_773_n853# 0 0.183f
C613 x1/x23/m1_891_n977# 0 1.14f
C614 x1/V9 0 0.591f
C615 x1/x23/m1_1725_85# 0 0.13f
C616 x1/x22/m1_451_n1105# 0 0.667f
C617 x1/V8 0 0.816f
C618 x1/x21/m1_400_n1066# 0 0.735f
C619 x1/V7 0 1.18f
C620 x1/V1 0 1.35f
C621 x1/x31/m1_931_n929# 0 2.11f
C622 x1/x20/m1_528_n874# 0 0.726f
C623 x1/V6 0 1.4f
C624 x1/x30/Vin 0 39.3f
C625 x1/th10_0/m1_718_n418# 0 0.567f
C626 x1/V10 0 0.761f
C627 x1/th10_0/m1_878_n414# 0 0.16f
.ends

