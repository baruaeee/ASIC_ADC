magic
tech sky130A
magscale 1 2
timestamp 1706270854
<< psubdiff >>
rect 1098 -727 1132 -673
<< nsubdiff >>
rect 367 382 441 416
rect 875 282 1047 316
<< locali >>
rect 375 382 404 416
rect 911 282 1070 316
rect 743 -249 777 -71
rect 689 -283 777 -249
rect 689 -724 723 -283
rect 669 -758 723 -724
rect 1098 -691 1132 -665
<< viali >>
rect 341 382 375 416
rect 877 282 911 316
rect 1098 -725 1132 -691
<< metal1 >>
rect 335 421 381 428
rect 658 421 758 452
rect 273 416 758 421
rect 273 387 341 416
rect 273 208 307 387
rect 335 382 341 387
rect 375 387 758 416
rect 375 382 381 387
rect 335 370 381 382
rect 658 352 758 387
rect 464 274 528 326
rect 871 316 917 328
rect 871 282 877 316
rect 911 282 917 316
rect 871 270 917 282
rect 273 174 457 208
rect 536 174 687 208
rect 653 161 687 174
rect 876 170 910 270
rect 740 161 794 170
rect 991 162 997 164
rect 653 127 794 161
rect 460 108 512 114
rect 740 110 794 127
rect 966 120 997 162
rect 991 112 997 120
rect 1049 112 1055 164
rect 460 50 512 56
rect 851 77 907 111
rect 851 21 885 77
rect 851 -13 948 21
rect 410 -61 777 -15
rect 410 -76 449 -61
rect 415 -115 449 -76
rect 741 -107 777 -61
rect 502 -495 536 -116
rect 741 -119 775 -107
rect 914 -113 948 -13
rect 1038 -113 1138 -84
rect 914 -147 1138 -113
rect 346 -528 446 -502
rect 914 -515 948 -147
rect 1038 -184 1138 -147
rect 346 -580 376 -528
rect 428 -580 446 -528
rect 885 -549 948 -515
rect 914 -550 948 -549
rect 346 -602 446 -580
rect 746 -608 752 -556
rect 804 -560 810 -556
rect 804 -608 836 -560
rect 788 -610 836 -608
rect 498 -620 550 -614
rect 498 -678 550 -672
rect 912 -689 946 -610
rect 992 -614 1046 -550
rect 1086 -689 1144 -685
rect 912 -691 1144 -689
rect 738 -737 838 -694
rect 912 -723 1098 -691
rect 912 -737 946 -723
rect 1086 -725 1098 -723
rect 1132 -725 1144 -691
rect 1086 -731 1144 -725
rect 738 -771 946 -737
rect 738 -794 838 -771
<< via1 >>
rect 997 112 1049 164
rect 460 56 512 108
rect 376 -580 428 -528
rect 752 -608 804 -556
rect 498 -672 550 -620
<< metal2 >>
rect 997 164 1049 170
rect 454 99 460 108
rect 274 65 460 99
rect 274 -537 308 65
rect 454 56 460 65
rect 512 56 518 108
rect 997 106 1049 112
rect 1006 -37 1040 106
rect 967 -71 1040 -37
rect 967 -431 1001 -71
rect 761 -465 1001 -431
rect 370 -537 376 -528
rect 274 -571 376 -537
rect 370 -580 376 -571
rect 428 -580 434 -528
rect 761 -550 795 -465
rect 752 -556 804 -550
rect 752 -614 804 -608
rect 492 -672 498 -620
rect 550 -629 556 -620
rect 752 -629 795 -614
rect 550 -663 795 -629
rect 550 -672 556 -663
use sky130_fd_pr__pfet_01v8_XGS3BL  XM0
timestamp 1706239161
transform 0 -1 591 1 0 -89
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_4L9AWD  XM1
timestamp 1706239161
transform 0 -1 522 1 0 -552
box -242 -252 242 252
use sky130_fd_pr__pfet_01v8_EZD9Q7  XM2
timestamp 1706239161
transform 1 0 496 0 1 191
box -224 -261 224 261
use sky130_fd_pr__pfet_01v8_M479BZ  XM3
timestamp 1706239161
transform 0 -1 879 1 0 141
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_4BNSKG  XM4
timestamp 1706239161
transform 0 -1 916 1 0 -580
box -214 -252 214 252
<< labels >>
flabel metal1 1038 -184 1138 -84 0 FreeSans 256 0 0 0 V10
port 1 nsew
flabel metal1 738 -794 838 -694 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 346 -602 446 -502 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 658 352 758 452 0 FreeSans 256 0 0 0 Vp
port 0 nsew
<< end >>
