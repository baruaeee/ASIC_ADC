magic
tech sky130A
magscale 1 2
timestamp 1705440135
<< pwell >>
rect 440 -1078 478 -938
rect 522 -976 586 -920
rect 540 -1164 574 -1130
<< psubdiff >>
rect 279 8 631 42
rect 279 -1231 313 8
rect 279 -1265 411 -1231
<< locali >>
rect 380 -136 418 -55
rect 592 -1088 734 -1016
rect 1024 -1082 1166 -1010
<< viali >>
rect 380 -55 418 -17
<< metal1 >>
rect 342 258 542 364
rect 639 297 803 359
rect 639 258 701 297
rect 0 0 200 200
rect 342 196 738 258
rect 797 229 895 263
rect 797 225 831 229
rect 833 225 895 229
rect 342 164 542 196
rect 380 105 418 164
rect 639 151 701 196
rect 797 191 895 225
rect 805 179 895 191
rect 459 117 511 123
rect 380 67 459 105
rect 380 -11 418 67
rect 639 89 799 151
rect 459 59 511 65
rect 861 -11 895 179
rect 368 -17 430 -11
rect 368 -55 380 -17
rect 418 -55 430 -17
rect 368 -61 430 -55
rect 629 -45 895 -11
rect 1016 -20 1216 180
rect 397 -123 431 -119
rect 629 -123 663 -45
rect 397 -157 663 -123
rect 0 -400 200 -200
rect 397 -281 431 -157
rect 528 -240 590 -188
rect 397 -291 507 -281
rect 742 -286 748 -234
rect 800 -286 806 -234
rect 958 -246 1018 -190
rect 1063 -279 1101 -20
rect 397 -343 525 -291
rect 586 -295 664 -290
rect 397 -357 509 -343
rect 585 -361 669 -295
rect 750 -298 806 -286
rect 1035 -289 1101 -279
rect 1025 -290 1101 -289
rect 750 -354 954 -298
rect 586 -364 669 -361
rect 588 -370 669 -364
rect 1024 -368 1101 -290
rect 342 -449 581 -415
rect 631 -420 669 -370
rect 1026 -372 1101 -368
rect 342 -592 376 -449
rect 631 -458 1029 -420
rect 0 -800 200 -600
rect 342 -792 542 -592
rect 0 -1200 200 -1000
rect 342 -1135 376 -792
rect 631 -853 669 -458
rect 1063 -519 1101 -372
rect 874 -557 1101 -519
rect 440 -891 837 -853
rect 440 -979 478 -891
rect 522 -976 586 -920
rect 440 -1009 489 -979
rect 440 -1075 525 -1009
rect 440 -1078 489 -1075
rect 592 -1078 733 -1020
rect 451 -1083 489 -1078
rect 540 -1135 574 -1130
rect 342 -1169 587 -1135
rect 675 -1231 733 -1078
rect 799 -1127 837 -891
rect 874 -999 912 -557
rect 1010 -792 1210 -592
rect 960 -972 1020 -918
rect 874 -1019 925 -999
rect 1127 -1019 1185 -792
rect 874 -1087 959 -1019
rect 1021 -1077 1189 -1019
rect 799 -1165 1015 -1127
rect 1131 -1231 1189 -1077
rect 675 -1289 1189 -1231
<< via1 >>
rect 459 65 511 117
rect 748 -286 800 -234
<< metal2 >>
rect 453 65 459 117
rect 511 65 517 117
rect 466 -47 504 65
rect 466 -85 793 -47
rect 755 -228 793 -85
rect 748 -234 800 -228
rect 748 -292 800 -286
use sky130_fd_pr__nfet_01v8_42G4RD  XM0
timestamp 1704404416
transform 1 0 556 0 1 -1048
box -218 -252 218 252
use sky130_fd_pr__pfet_01v8_DDPLQ8  XM1
timestamp 1704404416
transform 1 0 557 0 1 -325
box -215 -261 215 261
use sky130_fd_pr__nfet_01v8_VWP3K3  XM2
timestamp 1704404416
transform 1 0 767 0 1 224
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_LZD9A4  XM3
timestamp 1704404416
transform 1 0 988 0 1 -327
box -218 -261 218 261
use sky130_fd_pr__nfet_01v8_VRD6K3  XM4
timestamp 1704404416
transform 1 0 989 0 1 -1048
box -215 -252 215 252
<< labels >>
flabel metal1 1016 -20 1216 180 0 FreeSans 256 0 0 0 V04
port 1 nsew
flabel metal1 342 -792 542 -592 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 1010 -792 1210 -592 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 342 164 542 364 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 V04
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
<< end >>
