magic
tech sky130A
magscale 1 2
timestamp 1704418840
<< pwell >>
rect 548 -740 592 -680
rect 1544 -788 1618 -730
<< psubdiff >>
rect 1039 229 1173 263
rect 1139 -534 1173 229
rect 979 -568 1403 -534
<< locali >>
rect 1010 10 1398 64
rect 636 -884 696 -736
<< metal1 >>
rect 1122 528 1322 696
rect 1514 530 1580 584
rect 1120 496 1322 528
rect 522 486 574 490
rect 522 408 602 486
rect 1120 480 1196 496
rect 918 420 1196 480
rect 522 -130 574 408
rect 918 404 1524 420
rect 954 372 1006 404
rect 858 320 1006 372
rect 1118 344 1524 404
rect 1580 346 1828 422
rect 928 100 1576 152
rect 928 -122 980 100
rect 1752 -28 1828 346
rect 522 -202 598 -130
rect 896 -174 980 -122
rect 1640 -150 1840 -28
rect 900 -198 980 -174
rect 522 -210 574 -202
rect 414 -410 614 -396
rect 660 -410 712 -248
rect 414 -462 712 -410
rect 928 -444 980 -198
rect 1542 -228 1840 -150
rect 1542 -246 1682 -228
rect 1542 -414 1618 -246
rect 414 -596 614 -462
rect 782 -496 1504 -444
rect 510 -680 562 -596
rect 510 -738 592 -680
rect 782 -682 834 -496
rect 548 -740 592 -738
rect 770 -852 822 -736
rect 912 -742 968 -678
rect 1114 -852 1314 -716
rect 1544 -788 1618 -730
rect 1566 -852 1618 -788
rect 770 -904 1618 -852
rect 1114 -916 1314 -904
use sky130_fd_pr__nfet_01v8_8X7S4D  XM0
timestamp 1704418840
transform 0 -1 754 1 0 -709
box -211 -340 211 340
use sky130_fd_pr__pfet_01v8_GZD9X3  XM1
timestamp 1704418840
transform 1 0 749 0 1 -161
box -335 -261 335 261
use sky130_fd_pr__nfet_01v8_LH5FDA  XM2
timestamp 1704418840
transform 1 0 760 0 1 446
box -346 -252 346 252
use sky130_fd_pr__pfet_01v8_XJP3BL  XM3
timestamp 1704418840
transform 1 0 1551 0 1 337
box -211 -369 211 369
use sky130_fd_pr__nfet_01v8_LH5FDA  XM4
timestamp 1704418840
transform 0 -1 1584 1 0 -570
box -346 -252 346 252
<< labels >>
flabel metal1 1122 496 1322 696 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 1640 -228 1840 -28 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 1114 -916 1314 -716 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 414 -596 614 -396 0 FreeSans 256 0 0 0 Vin
port 2 nsew
<< end >>
