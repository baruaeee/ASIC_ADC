magic
tech sky130A
magscale 1 2
timestamp 1703792416
<< error_s >>
rect 8662 1446 8720 1452
rect 8662 1412 8674 1446
rect 8662 1406 8720 1412
rect 8662 1252 8720 1258
rect 8662 1218 8674 1252
rect 8662 1212 8720 1218
rect 8824 774 8882 780
rect 8824 740 8836 774
rect 8824 734 8882 740
rect 8824 562 8882 568
rect 8824 528 8836 562
rect 8824 522 8882 528
<< metal1 >>
rect 7084 2358 7284 2558
rect 5170 728 5370 928
rect 9618 816 9818 1016
rect 7064 -678 7264 -478
use sky130_fd_pr__pfet_01v8_MQKFYN  XM1
timestamp 1703732895
transform 1 0 6930 0 1 -133
box -1396 -261 1396 261
use sky130_fd_pr__nfet_01v8_RYBV7U  XM2
timestamp 1703732895
transform 1 0 6924 0 1 1976
box -1396 -252 1396 252
use sky130_fd_pr__pfet_01v8_VZ9GCW  XM3
timestamp 1703732895
transform -1 0 9172 0 1 1973
box -696 -261 696 261
use sky130_fd_pr__nfet_01v8_L7T3GD  XM4
timestamp 1703732895
transform 1 0 8691 0 1 1332
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_MQKFYN  XM5
timestamp 1703732895
transform 1 0 6924 0 1 651
box -1396 -261 1396 261
use sky130_fd_pr__nfet_01v8_RYBV7U  XM6
timestamp 1703732895
transform 1 0 6930 0 1 1328
box -1396 -252 1396 252
use sky130_fd_pr__pfet_01v8_M479BZ  XM7
timestamp 1703732895
transform 1 0 8853 0 1 651
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_LHZPBA  XM10
timestamp 1703732895
transform 1 0 9126 0 1 -142
box -646 -252 646 252
<< labels >>
flabel metal1 5170 728 5370 928 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 7064 -678 7264 -478 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 7084 2358 7284 2558 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 9618 816 9818 1016 0 FreeSans 256 0 0 0 Vout
port 2 nsew
<< end >>
