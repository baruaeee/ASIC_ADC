magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 2031 29 2037
rect -29 1997 -17 2031
rect -29 1991 29 1997
rect -29 -1997 29 -1991
rect -29 -2031 -17 -1997
rect -29 -2037 29 -2031
<< nwell >>
rect -211 -2169 211 2169
<< pmos >>
rect -15 -1950 15 1950
<< pdiff >>
rect -73 1938 -15 1950
rect -73 -1938 -61 1938
rect -27 -1938 -15 1938
rect -73 -1950 -15 -1938
rect 15 1938 73 1950
rect 15 -1938 27 1938
rect 61 -1938 73 1938
rect 15 -1950 73 -1938
<< pdiffc >>
rect -61 -1938 -27 1938
rect 27 -1938 61 1938
<< nsubdiff >>
rect -175 2099 -79 2133
rect 79 2099 175 2133
rect -175 2037 -141 2099
rect 141 2037 175 2099
rect -175 -2099 -141 -2037
rect 141 -2099 175 -2037
rect -175 -2133 -79 -2099
rect 79 -2133 175 -2099
<< nsubdiffcont >>
rect -79 2099 79 2133
rect -175 -2037 -141 2037
rect 141 -2037 175 2037
rect -79 -2133 79 -2099
<< poly >>
rect -33 2031 33 2047
rect -33 1997 -17 2031
rect 17 1997 33 2031
rect -33 1981 33 1997
rect -15 1950 15 1981
rect -15 -1981 15 -1950
rect -33 -1997 33 -1981
rect -33 -2031 -17 -1997
rect 17 -2031 33 -1997
rect -33 -2047 33 -2031
<< polycont >>
rect -17 1997 17 2031
rect -17 -2031 17 -1997
<< locali >>
rect -175 2099 -79 2133
rect 79 2099 175 2133
rect -175 2037 -141 2099
rect 141 2037 175 2099
rect -33 1997 -17 2031
rect 17 1997 33 2031
rect -61 1938 -27 1954
rect -61 -1954 -27 -1938
rect 27 1938 61 1954
rect 27 -1954 61 -1938
rect -33 -2031 -17 -1997
rect 17 -2031 33 -1997
rect -175 -2099 -141 -2037
rect 141 -2099 175 -2037
rect -175 -2133 -79 -2099
rect 79 -2133 175 -2099
<< viali >>
rect -17 1997 17 2031
rect -61 -1938 -27 1938
rect 27 -1938 61 1938
rect -17 -2031 17 -1997
<< metal1 >>
rect -29 2031 29 2037
rect -29 1997 -17 2031
rect 17 1997 29 2031
rect -29 1991 29 1997
rect -67 1938 -21 1950
rect -67 -1938 -61 1938
rect -27 -1938 -21 1938
rect -67 -1950 -21 -1938
rect 21 1938 67 1950
rect 21 -1938 27 1938
rect 61 -1938 67 1938
rect 21 -1950 67 -1938
rect -29 -1997 29 -1991
rect -29 -2031 -17 -1997
rect 17 -2031 29 -1997
rect -29 -2037 29 -2031
<< properties >>
string FIXED_BBOX -158 -2116 158 2116
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 19.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
