magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 181 29 187
rect -29 147 -17 181
rect -29 141 29 147
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect -29 -187 29 -181
<< nwell >>
rect -216 -319 216 319
<< pmos >>
rect -20 -100 20 100
<< pdiff >>
rect -78 88 -20 100
rect -78 -88 -66 88
rect -32 -88 -20 88
rect -78 -100 -20 -88
rect 20 88 78 100
rect 20 -88 32 88
rect 66 -88 78 88
rect 20 -100 78 -88
<< pdiffc >>
rect -66 -88 -32 88
rect 32 -88 66 88
<< nsubdiff >>
rect -180 249 -84 283
rect 84 249 180 283
rect -180 187 -146 249
rect 146 187 180 249
rect -180 -249 -146 -187
rect 146 -249 180 -187
rect -180 -283 -84 -249
rect 84 -283 180 -249
<< nsubdiffcont >>
rect -84 249 84 283
rect -180 -187 -146 187
rect 146 -187 180 187
rect -84 -283 84 -249
<< poly >>
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect -20 100 20 131
rect -20 -131 20 -100
rect -33 -147 33 -131
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -197 33 -181
<< polycont >>
rect -17 147 17 181
rect -17 -181 17 -147
<< locali >>
rect -180 249 -84 283
rect 84 249 180 283
rect -180 187 -146 249
rect 146 187 180 249
rect -33 147 -17 181
rect 17 147 33 181
rect -66 88 -32 104
rect -66 -104 -32 -88
rect 32 88 66 104
rect 32 -104 66 -88
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -180 -249 -146 -187
rect 146 -249 180 -187
rect -180 -283 -84 -249
rect 84 -283 180 -249
<< viali >>
rect -17 147 17 181
rect -66 -88 -32 88
rect 32 -88 66 88
rect -17 -181 17 -147
<< metal1 >>
rect -29 181 29 187
rect -29 147 -17 181
rect 17 147 29 181
rect -29 141 29 147
rect -72 88 -26 100
rect -72 -88 -66 88
rect -32 -88 -26 88
rect -72 -100 -26 -88
rect 26 88 72 100
rect 26 -88 32 88
rect 66 -88 72 88
rect 26 -100 72 -88
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect 17 -181 29 -147
rect -29 -187 29 -181
<< properties >>
string FIXED_BBOX -163 -266 163 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
