magic
tech sky130A
magscale 1 2
timestamp 1705440829
<< nwell >>
rect 722 -1022 776 -958
<< locali >>
rect 2068 272 2156 340
rect 2216 272 2470 340
rect 2402 -152 2470 272
rect 2022 -400 2241 -302
rect 1868 -872 1992 -814
rect 2902 -1166 3000 -1018
<< viali >>
rect 2156 272 2216 340
rect 2241 -400 2301 -302
rect 1992 -873 2052 -813
<< metal1 >>
rect 1300 700 1500 772
rect 1300 640 2274 700
rect 436 280 782 340
rect 1300 338 1500 640
rect 2214 472 2274 640
rect 2214 412 2582 472
rect 2214 352 2274 412
rect 3704 392 3802 480
rect 2150 340 2274 352
rect 436 -300 496 280
rect 948 80 1008 282
rect 1960 280 2020 340
rect 2150 272 2156 340
rect 2216 272 2274 340
rect 2150 260 2274 272
rect 1156 80 1216 86
rect 710 20 1156 80
rect 2214 70 2274 260
rect 2500 80 2560 86
rect 2714 80 2774 348
rect 300 -440 500 -300
rect 710 -388 770 20
rect 1156 14 1216 20
rect 2094 10 2274 70
rect 2384 20 2500 80
rect 2560 20 2774 80
rect 3742 44 3802 392
rect 1938 -314 1998 -300
rect 1908 -374 1998 -314
rect 1910 -380 1998 -374
rect 300 -500 918 -440
rect 1938 -674 1998 -380
rect 1594 -734 1998 -674
rect 722 -1022 776 -958
rect 1594 -962 1654 -734
rect 1986 -813 2058 -801
rect 2094 -813 2154 10
rect 2235 -302 2307 -290
rect 2235 -400 2241 -302
rect 2301 -400 2307 -302
rect 2235 -412 2307 -400
rect 1986 -873 1992 -813
rect 2052 -873 2154 -813
rect 1986 -885 2058 -873
rect 1756 -1000 1816 -958
rect 2242 -1000 2302 -412
rect 1674 -1060 2302 -1000
rect 2384 -424 2444 20
rect 2500 14 2560 20
rect 2840 -16 3802 44
rect 2840 -50 2900 -16
rect 2498 -110 2900 -50
rect 2498 -312 2558 -110
rect 2498 -382 2580 -312
rect 3700 -362 3802 -302
rect 2498 -384 2558 -382
rect 2384 -484 2650 -424
rect 2384 -970 2444 -484
rect 3742 -648 3802 -362
rect 3972 -648 4172 -600
rect 3504 -708 4172 -648
rect 3504 -964 3564 -708
rect 3972 -800 4172 -708
rect 2384 -1030 2580 -970
rect 2100 -1108 2302 -1060
rect 2762 -1108 2822 -1016
rect 3736 -1022 3796 -962
rect 2100 -1168 2822 -1108
rect 2100 -1200 2300 -1168
<< via1 >>
rect 1156 20 1216 80
rect 2500 20 2560 80
<< metal2 >>
rect 1150 20 1156 80
rect 1216 20 2500 80
rect 2560 20 2566 80
use sky130_fd_pr__pfet_01v8_XJ7SDL  XM0
timestamp 1704305861
transform 0 -1 1269 1 0 -989
box -211 -669 211 669
use sky130_fd_pr__nfet_01v8_ZFMUVB  XM1
timestamp 1704305861
transform 1 0 1346 0 1 -350
box -746 -252 746 252
use sky130_fd_pr__pfet_01v8_UJPVTG  XM2
timestamp 1704305861
transform 0 -1 1369 1 0 311
box -211 -769 211 769
use sky130_fd_pr__pfet_01v8_VZ9GTR  XM3
timestamp 1704305861
transform 1 0 3146 0 1 437
box -746 -261 746 261
use sky130_fd_pr__pfet_01v8_VZ9GTR  XM4
timestamp 1704305861
transform 1 0 3144 0 1 -341
box -746 -261 746 261
use sky130_fd_pr__nfet_01v8_9GNSAM  XM5
timestamp 1704305861
transform 0 -1 3158 1 0 -989
box -211 -760 211 760
<< labels >>
flabel metal1 2100 -1200 2300 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 1300 572 1500 772 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 300 -500 500 -300 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 3972 -800 4172 -600 0 FreeSans 256 0 0 0 Vout
port 1 nsew
<< end >>
