magic
tech sky130A
magscale 1 2
timestamp 1704962958
<< error_p >>
rect -29 391 29 397
rect -29 357 -17 391
rect -29 351 29 357
rect -29 -357 29 -351
rect -29 -391 -17 -357
rect -29 -397 29 -391
<< nwell >>
rect -211 -529 211 529
<< pmos >>
rect -15 -310 15 310
<< pdiff >>
rect -73 298 -15 310
rect -73 -298 -61 298
rect -27 -298 -15 298
rect -73 -310 -15 -298
rect 15 298 73 310
rect 15 -298 27 298
rect 61 -298 73 298
rect 15 -310 73 -298
<< pdiffc >>
rect -61 -298 -27 298
rect 27 -298 61 298
<< nsubdiff >>
rect -175 459 -79 493
rect 79 459 175 493
rect -175 397 -141 459
rect 141 397 175 459
rect -175 -459 -141 -397
rect 141 -459 175 -397
rect -175 -493 -79 -459
rect 79 -493 175 -459
<< nsubdiffcont >>
rect -79 459 79 493
rect -175 -397 -141 397
rect 141 -397 175 397
rect -79 -493 79 -459
<< poly >>
rect -33 391 33 407
rect -33 357 -17 391
rect 17 357 33 391
rect -33 341 33 357
rect -15 310 15 341
rect -15 -341 15 -310
rect -33 -357 33 -341
rect -33 -391 -17 -357
rect 17 -391 33 -357
rect -33 -407 33 -391
<< polycont >>
rect -17 357 17 391
rect -17 -391 17 -357
<< locali >>
rect -175 459 -79 493
rect 79 459 175 493
rect -175 397 -141 459
rect 141 397 175 459
rect -33 357 -17 391
rect 17 357 33 391
rect -61 298 -27 314
rect -61 -314 -27 -298
rect 27 298 61 314
rect 27 -314 61 -298
rect -33 -391 -17 -357
rect 17 -391 33 -357
rect -175 -459 -141 -397
rect 141 -459 175 -397
rect -175 -493 -79 -459
rect 79 -493 175 -459
<< viali >>
rect -17 357 17 391
rect -61 -298 -27 298
rect 27 -298 61 298
rect -17 -391 17 -357
<< metal1 >>
rect -29 391 29 397
rect -29 357 -17 391
rect 17 357 29 391
rect -29 351 29 357
rect -67 298 -21 310
rect -67 -298 -61 298
rect -27 -298 -21 298
rect -67 -310 -21 -298
rect 21 298 67 310
rect 21 -298 27 298
rect 61 -298 67 298
rect 21 -310 67 -298
rect -29 -357 29 -351
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -397 29 -391
<< properties >>
string FIXED_BBOX -158 -476 158 476
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.1 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
