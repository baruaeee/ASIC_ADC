************************************************************************
* auCdl Netlist:
* 
* Library Name:  ADC
* Top Cell Name: preampF_comm_B
* View Name:     schematic
* Netlisted on:  Dec  5 17:31:30 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: ADC
* Cell Name:    preampF_comm_B
* View Name:    schematic
************************************************************************

.SUBCKT preampF_comm_B A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MNM0 VDD A Y Y nfet_01v8 W=1.02u L=150n M=1
MPM1 VSS A Y Y pfet_01v8 W=550n L=1.05u M=1
.ENDS

