magic
tech sky130A
magscale 1 2
timestamp 1702941825
<< checkpaint >>
rect 2194 2339 5136 2546
rect -21 2258 5136 2339
rect -944 -766 5136 2258
rect -21 -819 5136 -766
rect 348 -872 5136 -819
rect 1271 -925 5136 -872
rect 2194 -978 5136 -925
<< error_s >>
rect 129 1431 187 1437
rect 129 1397 141 1431
rect 129 1391 187 1397
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_M4JX2X  XM1
timestamp 0
transform 1 0 158 0 1 1058
box -211 -511 211 511
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 0
transform 1 0 1450 0 1 760
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_YPGKLK  XM3
timestamp 0
transform 1 0 804 0 1 746
box -488 -252 488 252
use sky130_fd_pr__pfet_01v8_JRKFSA  XM7
timestamp 0
transform 1 0 2096 0 1 649
box -488 -261 488 261
use sky130_fd_pr__pfet_01v8_JRKFSA  XM9
timestamp 0
transform 1 0 3019 0 1 596
box -488 -261 488 261
use sky130_fd_pr__nfet_01v8_USW3YZ  XM10
timestamp 0
transform 1 0 3665 0 1 784
box -211 -502 211 502
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
