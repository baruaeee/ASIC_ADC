magic
tech sky130A
magscale 1 2
timestamp 1704305861
<< error_p >>
rect -29 631 29 637
rect -29 597 -17 631
rect -29 591 29 597
rect -29 -597 29 -591
rect -29 -631 -17 -597
rect -29 -637 29 -631
<< nwell >>
rect -211 -769 211 769
<< pmos >>
rect -15 -550 15 550
<< pdiff >>
rect -73 538 -15 550
rect -73 -538 -61 538
rect -27 -538 -15 538
rect -73 -550 -15 -538
rect 15 538 73 550
rect 15 -538 27 538
rect 61 -538 73 538
rect 15 -550 73 -538
<< pdiffc >>
rect -61 -538 -27 538
rect 27 -538 61 538
<< nsubdiff >>
rect -175 699 -79 733
rect 79 699 175 733
rect -175 637 -141 699
rect 141 637 175 699
rect -175 -699 -141 -637
rect 141 -699 175 -637
rect -175 -733 -79 -699
rect 79 -733 175 -699
<< nsubdiffcont >>
rect -79 699 79 733
rect -175 -637 -141 637
rect 141 -637 175 637
rect -79 -733 79 -699
<< poly >>
rect -33 631 33 647
rect -33 597 -17 631
rect 17 597 33 631
rect -33 581 33 597
rect -15 550 15 581
rect -15 -581 15 -550
rect -33 -597 33 -581
rect -33 -631 -17 -597
rect 17 -631 33 -597
rect -33 -647 33 -631
<< polycont >>
rect -17 597 17 631
rect -17 -631 17 -597
<< locali >>
rect -175 699 -79 733
rect 79 699 175 733
rect -175 637 -141 699
rect 141 637 175 699
rect -33 597 -17 631
rect 17 597 33 631
rect -61 538 -27 554
rect -61 -554 -27 -538
rect 27 538 61 554
rect 27 -554 61 -538
rect -33 -631 -17 -597
rect 17 -631 33 -597
rect -175 -699 -141 -637
rect 141 -699 175 -637
rect -175 -733 -79 -699
rect 79 -733 175 -699
<< viali >>
rect -17 597 17 631
rect -61 -538 -27 538
rect 27 -538 61 538
rect -17 -631 17 -597
<< metal1 >>
rect -29 631 29 637
rect -29 597 -17 631
rect 17 597 29 631
rect -29 591 29 597
rect -67 538 -21 550
rect -67 -538 -61 538
rect -27 -538 -21 538
rect -67 -550 -21 -538
rect 21 538 67 550
rect 21 -538 27 538
rect 61 -538 67 538
rect 21 -550 67 -538
rect -29 -597 29 -591
rect -29 -631 -17 -597
rect 17 -631 29 -597
rect -29 -637 29 -631
<< properties >>
string FIXED_BBOX -158 -716 158 716
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
