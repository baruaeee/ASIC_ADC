magic
tech sky130A
timestamp 1703732895
<< pwell >>
rect -323 -126 323 126
<< nmos >>
rect -225 -21 225 21
<< ndiff >>
rect -254 15 -225 21
rect -254 -15 -248 15
rect -231 -15 -225 15
rect -254 -21 -225 -15
rect 225 15 254 21
rect 225 -15 231 15
rect 248 -15 254 15
rect 225 -21 254 -15
<< ndiffc >>
rect -248 -15 -231 15
rect 231 -15 248 15
<< psubdiff >>
rect -305 91 -257 108
rect 257 91 305 108
rect -305 60 -288 91
rect 288 60 305 91
rect -305 -91 -288 -60
rect 288 -91 305 -60
rect -305 -108 -257 -91
rect 257 -108 305 -91
<< psubdiffcont >>
rect -257 91 257 108
rect -305 -60 -288 60
rect 288 -60 305 60
rect -257 -108 257 -91
<< poly >>
rect -225 57 225 65
rect -225 40 -217 57
rect 217 40 225 57
rect -225 21 225 40
rect -225 -40 225 -21
rect -225 -57 -217 -40
rect 217 -57 225 -40
rect -225 -65 225 -57
<< polycont >>
rect -217 40 217 57
rect -217 -57 217 -40
<< locali >>
rect -305 91 -257 108
rect 257 91 305 108
rect -305 60 -288 91
rect 288 60 305 91
rect -225 40 -217 57
rect 217 40 225 57
rect -248 15 -231 23
rect -248 -23 -231 -15
rect 231 15 248 23
rect 231 -23 248 -15
rect -225 -57 -217 -40
rect 217 -57 225 -40
rect -305 -91 -288 -60
rect 288 -91 305 -60
rect -305 -108 -257 -91
rect 257 -108 305 -91
<< viali >>
rect -217 40 217 57
rect -248 -15 -231 15
rect 231 -15 248 15
rect -217 -57 217 -40
<< metal1 >>
rect -223 57 223 60
rect -223 40 -217 57
rect 217 40 223 57
rect -223 37 223 40
rect -251 15 -228 21
rect -251 -15 -248 15
rect -231 -15 -228 15
rect -251 -21 -228 -15
rect 228 15 251 21
rect 228 -15 231 15
rect 248 -15 251 15
rect 228 -21 251 -15
rect -223 -40 223 -37
rect -223 -57 -217 -40
rect 217 -57 223 -40
rect -223 -60 223 -57
<< properties >>
string FIXED_BBOX -296 -99 296 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 4.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
