magic
tech sky130A
magscale 1 2
timestamp 1706203507
<< error_p >>
rect -29 144 29 150
rect -29 110 -17 144
rect -29 104 29 110
rect -29 -110 29 -104
rect -29 -144 -17 -110
rect -29 -150 29 -144
<< nwell >>
rect -211 -282 211 282
<< pmos >>
rect -15 -63 15 63
<< pdiff >>
rect -73 51 -15 63
rect -73 -51 -61 51
rect -27 -51 -15 51
rect -73 -63 -15 -51
rect 15 51 73 63
rect 15 -51 27 51
rect 61 -51 73 51
rect 15 -63 73 -51
<< pdiffc >>
rect -61 -51 -27 51
rect 27 -51 61 51
<< nsubdiff >>
rect -175 212 -79 246
rect 79 212 175 246
rect -175 150 -141 212
rect 141 150 175 212
rect -175 -212 -141 -150
rect 141 -212 175 -150
rect -175 -246 -79 -212
rect 79 -246 175 -212
<< nsubdiffcont >>
rect -79 212 79 246
rect -175 -150 -141 150
rect 141 -150 175 150
rect -79 -246 79 -212
<< poly >>
rect -33 144 33 160
rect -33 110 -17 144
rect 17 110 33 144
rect -33 94 33 110
rect -15 63 15 94
rect -15 -94 15 -63
rect -33 -110 33 -94
rect -33 -144 -17 -110
rect 17 -144 33 -110
rect -33 -160 33 -144
<< polycont >>
rect -17 110 17 144
rect -17 -144 17 -110
<< locali >>
rect -175 212 -79 246
rect 79 212 175 246
rect -175 150 -141 212
rect 141 150 175 212
rect -33 110 -17 144
rect 17 110 33 144
rect -61 51 -27 67
rect -61 -67 -27 -51
rect 27 51 61 67
rect 27 -67 61 -51
rect -33 -144 -17 -110
rect 17 -144 33 -110
rect -175 -212 -141 -150
rect 141 -212 175 -150
rect -175 -246 -79 -212
rect 79 -246 175 -212
<< viali >>
rect -17 110 17 144
rect -61 -51 -27 51
rect 27 -51 61 51
rect -17 -144 17 -110
<< metal1 >>
rect -29 144 29 150
rect -29 110 -17 144
rect 17 110 29 144
rect -29 104 29 110
rect -67 51 -21 63
rect -67 -51 -61 51
rect -27 -51 -21 51
rect -67 -63 -21 -51
rect 21 51 67 63
rect 21 -51 27 51
rect 61 -51 67 51
rect 21 -63 67 -51
rect -29 -110 29 -104
rect -29 -144 -17 -110
rect 17 -144 29 -110
rect -29 -150 29 -144
<< properties >>
string FIXED_BBOX -158 -229 158 229
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.63 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
