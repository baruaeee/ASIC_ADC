magic
tech sky130A
magscale 1 2
timestamp 1704962958
<< error_p >>
rect -29 382 29 388
rect -29 348 -17 382
rect -29 342 29 348
rect -29 -348 29 -342
rect -29 -382 -17 -348
rect -29 -388 29 -382
<< pwell >>
rect -211 -520 211 520
<< nmos >>
rect -15 -310 15 310
<< ndiff >>
rect -73 298 -15 310
rect -73 -298 -61 298
rect -27 -298 -15 298
rect -73 -310 -15 -298
rect 15 298 73 310
rect 15 -298 27 298
rect 61 -298 73 298
rect 15 -310 73 -298
<< ndiffc >>
rect -61 -298 -27 298
rect 27 -298 61 298
<< psubdiff >>
rect -175 450 -79 484
rect 79 450 175 484
rect -175 388 -141 450
rect 141 388 175 450
rect -175 -450 -141 -388
rect 141 -450 175 -388
rect -175 -484 -79 -450
rect 79 -484 175 -450
<< psubdiffcont >>
rect -79 450 79 484
rect -175 -388 -141 388
rect 141 -388 175 388
rect -79 -484 79 -450
<< poly >>
rect -33 382 33 398
rect -33 348 -17 382
rect 17 348 33 382
rect -33 332 33 348
rect -15 310 15 332
rect -15 -332 15 -310
rect -33 -348 33 -332
rect -33 -382 -17 -348
rect 17 -382 33 -348
rect -33 -398 33 -382
<< polycont >>
rect -17 348 17 382
rect -17 -382 17 -348
<< locali >>
rect -175 450 -79 484
rect 79 450 175 484
rect -175 388 -141 450
rect 141 388 175 450
rect -33 348 -17 382
rect 17 348 33 382
rect -61 298 -27 314
rect -61 -314 -27 -298
rect 27 298 61 314
rect 27 -314 61 -298
rect -33 -382 -17 -348
rect 17 -382 33 -348
rect -175 -450 -141 -388
rect 141 -450 175 -388
rect -175 -484 -79 -450
rect 79 -484 175 -450
<< viali >>
rect -17 348 17 382
rect -61 -298 -27 298
rect 27 -298 61 298
rect -17 -382 17 -348
<< metal1 >>
rect -29 382 29 388
rect -29 348 -17 382
rect 17 348 29 382
rect -29 342 29 348
rect -67 298 -21 310
rect -67 -298 -61 298
rect -27 -298 -21 298
rect -67 -310 -21 -298
rect 21 298 67 310
rect 21 -298 27 298
rect 61 -298 67 298
rect 21 -310 67 -298
rect -29 -348 29 -342
rect -29 -382 -17 -348
rect 17 -382 29 -348
rect -29 -388 29 -382
<< properties >>
string FIXED_BBOX -158 -467 158 467
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.1 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
