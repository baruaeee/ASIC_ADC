magic
tech sky130A
magscale 1 2
timestamp 1706474503
<< nwell >>
rect 438 536 1266 646
<< psubdiff >>
rect 1016 -303 1050 -231
<< locali >>
rect 800 362 834 511
rect 1445 -210 1479 -131
rect 1027 -266 1052 -232
rect 1134 -244 1479 -210
rect 1802 -395 1915 -361
<< viali >>
rect 993 -266 1027 -232
rect 1915 -395 1949 -361
<< metal1 >>
rect 1190 609 1290 644
rect 860 575 1401 609
rect 556 330 614 366
rect 860 364 894 575
rect 1190 544 1290 575
rect 1367 425 1401 575
rect 544 278 550 330
rect 602 314 614 330
rect 602 278 608 314
rect 831 275 1053 309
rect 1176 302 1232 368
rect 1367 353 1433 425
rect 1859 411 1893 417
rect 1859 377 1989 411
rect 1859 357 1893 377
rect 1019 271 1053 275
rect 1465 271 1685 299
rect 1019 237 1685 271
rect 618 56 682 112
rect 708 3 742 4
rect 559 -173 625 1
rect 679 -173 742 3
rect 1019 -84 1053 237
rect 1955 130 1989 377
rect 1938 127 2038 130
rect 1481 93 2038 127
rect 1481 -16 1515 93
rect 1938 30 2038 93
rect 1481 -41 1516 -16
rect 1375 -75 1593 -41
rect 1482 -76 1516 -75
rect 1019 -85 1252 -84
rect 1019 -119 1271 -85
rect 1214 -120 1248 -119
rect 559 -424 593 -173
rect 707 -178 742 -173
rect 704 -222 742 -178
rect 1755 -211 1789 -87
rect 656 -233 742 -222
rect 987 -232 1033 -220
rect 987 -233 993 -232
rect 631 -266 993 -233
rect 1027 -233 1033 -232
rect 1027 -266 1049 -233
rect 631 -267 1049 -266
rect 1720 -245 1789 -211
rect 987 -278 1033 -267
rect 1131 -424 1165 -399
rect 1720 -401 1754 -245
rect 559 -458 1165 -424
rect 1687 -459 1754 -401
rect 1884 -361 1984 -320
rect 1884 -395 1915 -361
rect 1949 -395 1984 -361
rect 1884 -420 1984 -395
rect 862 -518 962 -504
rect 862 -570 905 -518
rect 957 -532 962 -518
rect 1233 -532 1531 -507
rect 957 -541 1531 -532
rect 957 -566 1371 -541
rect 957 -570 962 -566
rect 862 -604 962 -570
<< via1 >>
rect 550 278 602 330
rect 905 -570 957 -518
<< metal2 >>
rect 550 330 602 336
rect 550 272 602 278
rect 559 223 593 272
rect 559 189 948 223
rect 914 -518 948 189
rect 899 -570 905 -518
rect 957 -570 963 -518
use sky130_fd_pr__pfet_01v8_XGS3BL  XM0
timestamp 1706239161
transform -1 0 651 0 -1 -85
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_ZFRTVB  XM1
timestamp 1706197322
transform 1 0 1426 0 1 -428
box -446 -252 456 252
use sky130_fd_pr__pfet_01v8_XQZLDL  XM2
timestamp 1706197322
transform 0 -1 897 1 0 335
box -211 -459 211 459
use sky130_fd_pr__pfet_01v8_VZ9GC6  XM3
timestamp 1706197322
transform 1 0 1646 0 1 385
box -396 -261 396 261
use sky130_fd_pr__nfet_01v8_ATLS57  XM4
timestamp 1706197322
transform 0 -1 1508 1 0 -103
box -211 -410 211 410
<< labels >>
flabel metal1 1938 30 2038 130 0 FreeSans 256 0 0 0 V13
port 1 nsew
flabel metal1 1884 -420 1984 -320 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 1190 544 1290 644 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 862 -604 962 -504 0 FreeSans 256 0 0 0 Vin
port 2 nsew
<< end >>
