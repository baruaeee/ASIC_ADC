* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : inv01f                                       *
* Netlisted  : Sun Dec  8 22:28:22 2024                     *
* Pegasus Version: 23.11-s009 Thu Aug 31 12:45:19 PDT 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_733693291110                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_733693291110 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=6.5e-07 W=4.45e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_733693291110

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_733693291111                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_733693291111 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=6.3e-07 W=7.9e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_733693291111

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv01f                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv01f 3 4 1 2
** N=9 EP=4 FDC=2
X0 1 2 3 nfet_01v8_CDNS_733693291110 $T=295 475 0 0 $X=-110 $Y=325
X1 4 2 3 pfet_01v8_CDNS_733693291111 $T=295 2820 0 0 $X=-150 $Y=2640
.ends inv01f
