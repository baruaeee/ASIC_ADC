magic
tech sky130A
magscale 1 2
timestamp 1696298453
<< nwell >>
rect -211 -2719 211 2719
<< pmos >>
rect -15 -2500 15 2500
<< pdiff >>
rect -73 2488 -15 2500
rect -73 -2488 -61 2488
rect -27 -2488 -15 2488
rect -73 -2500 -15 -2488
rect 15 2488 73 2500
rect 15 -2488 27 2488
rect 61 -2488 73 2488
rect 15 -2500 73 -2488
<< pdiffc >>
rect -61 -2488 -27 2488
rect 27 -2488 61 2488
<< nsubdiff >>
rect -175 2649 -79 2683
rect 79 2649 175 2683
rect -175 2587 -141 2649
rect 141 2587 175 2649
rect -175 -2649 -141 -2587
rect 141 -2649 175 -2587
rect -175 -2683 -79 -2649
rect 79 -2683 175 -2649
<< nsubdiffcont >>
rect -79 2649 79 2683
rect -175 -2587 -141 2587
rect 141 -2587 175 2587
rect -79 -2683 79 -2649
<< poly >>
rect -33 2581 33 2597
rect -33 2547 -17 2581
rect 17 2547 33 2581
rect -33 2531 33 2547
rect -15 2500 15 2531
rect -15 -2531 15 -2500
rect -33 -2547 33 -2531
rect -33 -2581 -17 -2547
rect 17 -2581 33 -2547
rect -33 -2597 33 -2581
<< polycont >>
rect -17 2547 17 2581
rect -17 -2581 17 -2547
<< locali >>
rect -175 2649 -79 2683
rect 79 2649 175 2683
rect -175 2587 -141 2649
rect 141 2587 175 2649
rect -33 2547 -17 2581
rect 17 2547 33 2581
rect -61 2488 -27 2504
rect -61 -2504 -27 -2488
rect 27 2488 61 2504
rect 27 -2504 61 -2488
rect -33 -2581 -17 -2547
rect 17 -2581 33 -2547
rect -175 -2649 -141 -2587
rect 141 -2649 175 -2587
rect -175 -2683 -79 -2649
rect 79 -2683 175 -2649
<< viali >>
rect -17 2547 17 2581
rect -61 -2488 -27 2488
rect 27 -2488 61 2488
rect -17 -2581 17 -2547
<< metal1 >>
rect -32 2581 32 2596
rect -32 2547 -17 2581
rect 17 2547 32 2581
rect -32 2542 32 2547
rect -29 2541 29 2542
rect -67 2488 -21 2500
rect -67 -2488 -61 2488
rect -27 -2488 -21 2488
rect -67 -2500 -21 -2488
rect 21 2488 67 2500
rect 21 -2488 27 2488
rect 61 -2488 67 2488
rect 21 -2500 67 -2488
rect -32 -2547 32 -2540
rect -32 -2581 -17 -2547
rect 17 -2581 32 -2547
rect -32 -2594 32 -2581
<< properties >>
string FIXED_BBOX -158 -2666 158 2666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 25.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
