magic
tech sky130A
magscale 1 2
timestamp 1704501257
<< nwell >>
rect -1296 -261 1296 261
<< pmos >>
rect -1100 -42 1100 42
<< pdiff >>
rect -1158 30 -1100 42
rect -1158 -30 -1146 30
rect -1112 -30 -1100 30
rect -1158 -42 -1100 -30
rect 1100 30 1158 42
rect 1100 -30 1112 30
rect 1146 -30 1158 30
rect 1100 -42 1158 -30
<< pdiffc >>
rect -1146 -30 -1112 30
rect 1112 -30 1146 30
<< nsubdiff >>
rect -1260 191 -1164 225
rect 1164 191 1260 225
rect -1260 129 -1226 191
rect 1226 129 1260 191
rect -1260 -191 -1226 -129
rect 1226 -191 1260 -129
rect -1260 -225 -1164 -191
rect 1164 -225 1260 -191
<< nsubdiffcont >>
rect -1164 191 1164 225
rect -1260 -129 -1226 129
rect 1226 -129 1260 129
rect -1164 -225 1164 -191
<< poly >>
rect -1100 123 1100 139
rect -1100 89 -1084 123
rect 1084 89 1100 123
rect -1100 42 1100 89
rect -1100 -89 1100 -42
rect -1100 -123 -1084 -89
rect 1084 -123 1100 -89
rect -1100 -139 1100 -123
<< polycont >>
rect -1084 89 1084 123
rect -1084 -123 1084 -89
<< locali >>
rect -1260 191 -1164 225
rect 1164 191 1260 225
rect -1260 129 -1226 191
rect 1226 129 1260 191
rect -1100 89 -1084 123
rect 1084 89 1100 123
rect -1146 30 -1112 46
rect -1146 -46 -1112 -30
rect 1112 30 1146 46
rect 1112 -46 1146 -30
rect -1100 -123 -1084 -89
rect 1084 -123 1100 -89
rect -1260 -191 -1226 -129
rect 1226 -191 1260 -129
rect -1260 -225 -1164 -191
rect 1164 -225 1260 -191
<< viali >>
rect -1084 89 1084 123
rect -1146 -30 -1112 30
rect 1112 -30 1146 30
rect -1084 -123 1084 -89
<< metal1 >>
rect -1096 123 1096 129
rect -1096 89 -1084 123
rect 1084 89 1096 123
rect -1096 83 1096 89
rect -1152 30 -1106 42
rect -1152 -30 -1146 30
rect -1112 -30 -1106 30
rect -1152 -42 -1106 -30
rect 1106 30 1152 42
rect 1106 -30 1112 30
rect 1146 -30 1152 30
rect 1106 -42 1152 -30
rect -1096 -89 1096 -83
rect -1096 -123 -1084 -89
rect 1084 -123 1096 -89
rect -1096 -129 1096 -123
<< properties >>
string FIXED_BBOX -1243 -208 1243 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 11.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
