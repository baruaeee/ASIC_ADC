magic
tech sky130A
magscale 1 2
timestamp 1706392731
<< metal1 >>
rect 6910 7096 6956 7245
rect 8595 7180 8641 7299
rect 8592 7174 8644 7180
rect 8592 7116 8644 7122
rect 6901 7044 6907 7096
rect 6959 7044 6965 7096
<< via1 >>
rect 8592 7122 8644 7174
rect 6907 7044 6959 7096
<< metal2 >>
rect 8586 7171 8592 7174
rect 8460 7125 8592 7171
rect 6907 7096 6959 7102
rect 6907 7038 6959 7044
rect 6911 6825 6954 7038
rect 8460 6741 8506 7125
rect 8586 7122 8592 7125
rect 8644 7122 8650 7174
use therm  therm_0
timestamp 1706387947
transform 1 0 4297 0 1 72
box -435 1094 7123 6820
use Analog  x1
timestamp 1706392731
transform 1 0 0 0 1 7400
box 3657 -3483 10185 809
<< end >>
