magic
tech sky130A
magscale 1 2
timestamp 1704371799
<< pwell >>
rect -353 -252 353 252
<< nmos >>
rect -157 -42 157 42
<< ndiff >>
rect -215 30 -157 42
rect -215 -30 -203 30
rect -169 -30 -157 30
rect -215 -42 -157 -30
rect 157 30 215 42
rect 157 -30 169 30
rect 203 -30 215 30
rect 157 -42 215 -30
<< ndiffc >>
rect -203 -30 -169 30
rect 169 -30 203 30
<< psubdiff >>
rect -317 182 -221 216
rect 221 182 317 216
rect -317 120 -283 182
rect 283 120 317 182
rect -317 -182 -283 -120
rect 283 -182 317 -120
rect -317 -216 -221 -182
rect 221 -216 317 -182
<< psubdiffcont >>
rect -221 182 221 216
rect -317 -120 -283 120
rect 283 -120 317 120
rect -221 -216 221 -182
<< poly >>
rect -157 114 157 130
rect -157 80 -141 114
rect 141 80 157 114
rect -157 42 157 80
rect -157 -80 157 -42
rect -157 -114 -141 -80
rect 141 -114 157 -80
rect -157 -130 157 -114
<< polycont >>
rect -141 80 141 114
rect -141 -114 141 -80
<< locali >>
rect -317 182 -221 216
rect 221 182 317 216
rect -317 120 -283 182
rect 283 120 317 182
rect -157 80 -141 114
rect 141 80 157 114
rect -203 30 -169 46
rect -203 -46 -169 -30
rect 169 30 203 46
rect 169 -46 203 -30
rect -157 -114 -141 -80
rect 141 -114 157 -80
rect -317 -182 -283 -120
rect 283 -182 317 -120
rect -317 -216 -221 -182
rect 221 -216 317 -182
<< viali >>
rect -141 80 141 114
rect -203 -30 -169 30
rect 169 -30 203 30
rect -141 -114 141 -80
<< metal1 >>
rect -153 114 153 120
rect -153 80 -141 114
rect 141 80 153 114
rect -153 74 153 80
rect -209 30 -163 42
rect -209 -30 -203 30
rect -169 -30 -163 30
rect -209 -42 -163 -30
rect 163 30 209 42
rect 163 -30 169 30
rect 203 -30 209 30
rect 163 -42 209 -30
rect -153 -80 153 -74
rect -153 -114 -141 -80
rect 141 -114 153 -80
rect -153 -120 153 -114
<< properties >>
string FIXED_BBOX -300 -199 300 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 1.57 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
