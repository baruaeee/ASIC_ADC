* NGSPICE file created from th15.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_MYW2PY a_n73_n48# a_n33_n145# a_15_n48# w_n211_n267#
+ VSUBS
X0 a_15_n48# a_n33_n145# a_n73_n48# w_n211_n267# sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.54 as=0.139 ps=1.54 w=0.48 l=0.15
C0 a_15_n48# w_n211_n267# 0.05f
C1 a_15_n48# a_n33_n145# 0.0197f
C2 a_15_n48# a_n73_n48# 0.0795f
C3 a_n33_n145# w_n211_n267# 0.237f
C4 a_n73_n48# w_n211_n267# 0.05f
C5 a_n33_n145# a_n73_n48# 0.0197f
C6 a_15_n48# VSUBS 0.0287f
C7 a_n73_n48# VSUBS 0.0287f
C8 a_n33_n145# VSUBS 0.115f
C9 w_n211_n267# VSUBS 1.05f
.ends

.subckt sky130_fd_pr__nfet_01v8_JRGCPP a_n1108_n42# a_1050_n42# a_n1210_n216# a_n1050_n130#
X0 a_1050_n42# a_n1050_n130# a_n1108_n42# a_n1210_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=10.5
C0 a_n1108_n42# a_n1050_n130# 0.0251f
C1 a_1050_n42# a_n1050_n130# 0.0251f
C2 a_1050_n42# a_n1210_n216# 0.0931f
C3 a_n1108_n42# a_n1210_n216# 0.0931f
C4 a_n1050_n130# a_n1210_n216# 5.94f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJ78MR a_n73_n1050# w_n211_n1269# a_15_n1050# a_n33_n1147#
+ VSUBS
X0 a_15_n1050# a_n33_n1147# a_n73_n1050# w_n211_n1269# sky130_fd_pr__pfet_01v8 ad=3.05 pd=21.6 as=3.05 ps=21.6 w=10.5 l=0.15
C0 a_15_n1050# w_n211_n1269# 0.661f
C1 a_15_n1050# a_n33_n1147# 0.065f
C2 a_15_n1050# a_n73_n1050# 1.67f
C3 a_n33_n1147# w_n211_n1269# 0.242f
C4 a_n73_n1050# w_n211_n1269# 0.661f
C5 a_n33_n1147# a_n73_n1050# 0.065f
C6 a_15_n1050# VSUBS 0.434f
C7 a_n73_n1050# VSUBS 0.434f
C8 a_n33_n1147# VSUBS 0.129f
C9 w_n211_n1269# VSUBS 4.56f
.ends

.subckt sky130_fd_pr__pfet_01v8_6M437L a_n1108_n42# a_1050_n42# a_n1050_n139# w_n1246_n261#
+ VSUBS
X0 a_1050_n42# a_n1050_n139# a_n1108_n42# w_n1246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=10.5
C0 a_1050_n42# w_n1246_n261# 0.0498f
C1 a_1050_n42# a_n1050_n139# 0.0251f
C2 a_n1050_n139# w_n1246_n261# 3.36f
C3 a_n1108_n42# w_n1246_n261# 0.0498f
C4 a_n1050_n139# a_n1108_n42# 0.0251f
C5 a_1050_n42# VSUBS 0.0428f
C6 a_n1108_n42# VSUBS 0.0428f
C7 a_n1050_n139# VSUBS 2.7f
C8 w_n1246_n261# VSUBS 5.27f
.ends

.subckt sky130_fd_pr__nfet_01v8_A5ES5P a_n73_n1000# a_15_n1000# a_n33_n1088# a_n175_n1174#
X0 a_15_n1000# a_n33_n1088# a_n73_n1000# a_n175_n1174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.6 as=2.9 ps=20.6 w=10 l=0.15
C0 a_n73_n1000# a_n33_n1088# 0.0649f
C1 a_15_n1000# a_n33_n1088# 0.0649f
C2 a_n73_n1000# a_15_n1000# 1.59f
C3 a_15_n1000# a_n175_n1174# 1.04f
C4 a_n73_n1000# a_n175_n1174# 1.04f
C5 a_n33_n1088# a_n175_n1174# 0.359f
.ends

.subckt th15 Vp Vout Vin Vn
XXM0 m1_915_n714# Vn Vn Vp Vn sky130_fd_pr__pfet_01v8_MYW2PY
XXM1 m1_1074_6# m1_915_n714# Vn Vin sky130_fd_pr__nfet_01v8_JRGCPP
XXM2 v1 m1_1074_6# Vn Vin sky130_fd_pr__nfet_01v8_JRGCPP
XXM3 v1 Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_XJ78MR
XXM4 Vp m1_4024_602# v1 Vp Vn sky130_fd_pr__pfet_01v8_6M437L
XXM5 Vn Vout v1 Vn sky130_fd_pr__nfet_01v8_A5ES5P
XXM7 m1_4024_602# Vout v1 Vp Vn sky130_fd_pr__pfet_01v8_6M437L
C0 Vn m1_4024_602# -4.17e-25
C1 Vn Vout 0.0294f
C2 m1_1074_6# v1 0.0103f
C3 Vn Vp 1.35f
C4 Vin Vn 0.17f
C5 m1_1074_6# Vp 0.0774f
C6 m1_1074_6# Vin 1.03f
C7 v1 m1_4024_602# 0.999f
C8 Vn m1_915_n714# 0.388f
C9 Vout v1 0.214f
C10 Vp v1 1.22f
C11 Vout m1_4024_602# 0.00816f
C12 m1_1074_6# m1_915_n714# 0.0137f
C13 Vin v1 0.641f
C14 Vp m1_4024_602# 0.404f
C15 Vp Vout 0.129f
C16 Vin m1_4024_602# 1.79e-19
C17 Vin Vp 0.222f
C18 m1_915_n714# v1 3.02e-20
C19 m1_1074_6# Vn 0.201f
C20 m1_915_n714# Vp 0.596f
C21 Vin m1_915_n714# 0.378f
C22 Vn v1 0.15f
C23 Vin 0 11.3f
C24 m1_4024_602# 0 0.411f
C25 Vout 0 1.43f
C26 v1 0 6.08f
C27 m1_1074_6# 0 0.643f
C28 Vn 0 1.59f
C29 m1_915_n714# 0 0.787f
C30 Vp 0 17.1f
.ends

