** sch_path: /home/exotic/Desktop/ASIC_ADC/xschem/Vth_sch/Pre_layout/th11.sch
**.subckt th11 Vin Vout
*.ipin Vin
*.opin Vout
VDD VDD GND 1.8
Vin Vin GND pulse(0 0.2 0ns 1ns 1ns 5ns 10ns)
V_logic_high V_LH GND 1.25
V_logic_low V_LL GND 0.5
x1 VDD Vout Vin GND th11
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.save all





.dc Vin 0 1.8 0.01
*.tran 1n 30n
.control
run
set color0=white
set color1=black
plot Vin Vout V_LH V_LL
set xbrushwidth=3
.save all
.endc
.end


**** end user architecture code
**.ends

* NGSPICE file created from th11.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_XGAKDL a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
+ VSUBS
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_15_n200# a_n73_n200# 0.321f
C1 w_n211_n419# a_n73_n200# 0.143f
C2 a_n33_n297# a_n73_n200# 0.0293f
C3 w_n211_n419# a_15_n200# 0.143f
C4 a_n33_n297# a_15_n200# 0.0293f
C5 w_n211_n419# a_n33_n297# 0.24f
C6 a_15_n200# VSUBS 0.0902f
C7 a_n73_n200# VSUBS 0.0902f
C8 a_n33_n297# VSUBS 0.119f
C9 w_n211_n419# VSUBS 1.58f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFH27D a_50_n42# a_n210_n216# a_n108_n42# a_n50_n130#
X0 a_50_n42# a_n50_n130# a_n108_n42# a_n210_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 a_n50_n130# a_50_n42# 0.00909f
C1 a_n108_n42# a_50_n42# 0.0391f
C2 a_n50_n130# a_n108_n42# 0.00909f
C3 a_50_n42# a_n210_n216# 0.0801f
C4 a_n108_n42# a_n210_n216# 0.0801f
C5 a_n50_n130# a_n210_n216# 0.439f
.ends

.subckt sky130_fd_pr__pfet_01v8_E7ZT25 a_15_n43# w_n211_n262# a_n73_n43# a_n33_n140#
+ VSUBS
X0 a_15_n43# a_n33_n140# a_n73_n43# w_n211_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.15
C0 a_15_n43# a_n73_n43# 0.0715f
C1 w_n211_n262# a_n73_n43# 0.0469f
C2 a_n33_n140# a_n73_n43# 0.0193f
C3 w_n211_n262# a_15_n43# 0.0469f
C4 a_n33_n140# a_15_n43# 0.0193f
C5 w_n211_n262# a_n33_n140# 0.236f
C6 a_15_n43# VSUBS 0.0267f
C7 a_n73_n43# VSUBS 0.0267f
C8 a_n33_n140# VSUBS 0.115f
C9 w_n211_n262# VSUBS 1.03f
.ends

.subckt sky130_fd_pr__pfet_01v8_JM8GTH a_50_n42# w_n246_n261# a_n50_n139# a_n108_n42#
+ VSUBS
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 a_50_n42# a_n108_n42# 0.0391f
C1 w_n246_n261# a_n108_n42# 0.0499f
C2 a_n50_n139# a_n108_n42# 0.00909f
C3 w_n246_n261# a_50_n42# 0.0499f
C4 a_n50_n139# a_50_n42# 0.00909f
C5 w_n246_n261# a_n50_n139# 0.279f
C6 a_50_n42# VSUBS 0.0298f
C7 a_n108_n42# VSUBS 0.0298f
C8 a_n50_n139# VSUBS 0.175f
C9 w_n246_n261# VSUBS 1.18f
.ends

.subckt sky130_fd_pr__nfet_01v8_L9ESAD a_n175_n224# a_n73_n50# a_n33_n138# a_15_n50#
X0 a_15_n50# a_n33_n138# a_n73_n50# a_n175_n224# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_n33_n138# a_15_n50# 0.0216f
C1 a_n73_n50# a_15_n50# 0.0826f
C2 a_n33_n138# a_n73_n50# 0.0216f
C3 a_15_n50# a_n175_n224# 0.081f
C4 a_n73_n50# a_n175_n224# 0.081f
C5 a_n33_n138# a_n175_n224# 0.339f
.ends

.subckt th11 Vp V11 Vin Vn
XXM0 m1_717_301# Vp Vn Vn Vn sky130_fd_pr__pfet_01v8_XGAKDL
XXM1 m1_717_301# Vn m1_509_303# Vin sky130_fd_pr__nfet_01v8_ZFH27D
XXM2 m1_509_303# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_E7ZT25
XXM3 V11 Vp m1_509_303# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM4 Vn Vn m1_509_303# V11 sky130_fd_pr__nfet_01v8_L9ESAD
C0 Vin m1_509_303# 0.248f
C1 m1_717_301# Vp 0.0487f
C2 V11 m1_717_301# 1.71e-20
C3 V11 Vp 0.0686f
C4 m1_717_301# m1_509_303# 0.0301f
C5 m1_509_303# Vp 0.352f
C6 V11 m1_509_303# 0.0742f
C7 m1_717_301# Vin 0.0345f
C8 Vin Vp 0.258f
C9 V11 Vin 0.00112f
C10 Vin Vn 0.856f
C11 m1_509_303# Vn 0.717f
C12 Vp Vn 4.47f
C13 V11 Vn 0.485f
C14 m1_717_301# Vn 0.299f
.ends


.GLOBAL VDD
.GLOBAL GND
.GLOBAL V_LH
.GLOBAL V_LL
.end
