magic
tech sky130A
magscale 1 2
timestamp 1702941826
<< checkpaint >>
rect 14342 2099 17284 2118
rect 10103 -925 17284 2099
rect 14342 -978 17284 -925
<< error_s >>
rect 10807 5723 10865 5729
rect 10807 5689 10819 5723
rect 10807 5683 10865 5689
rect 10977 4726 11011 4744
rect 10977 4690 11047 4726
rect 10994 4656 11065 4690
rect 5268 999 5303 1033
rect 10661 1016 10695 1034
rect 5269 980 5303 999
rect 5288 583 5303 980
rect 5322 946 5357 980
rect 5322 583 5356 946
rect 5322 549 5337 583
rect 10625 530 10695 1016
rect 10807 613 10865 619
rect 10807 579 10819 613
rect 10807 573 10865 579
rect 10625 494 10678 530
rect 10994 477 11064 4656
rect 11176 4588 11234 4594
rect 11176 4554 11188 4588
rect 11176 4548 11234 4554
rect 11176 560 11234 566
rect 11176 526 11188 560
rect 11176 520 11234 526
rect 10994 441 11047 477
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_XJP7MR  XM1
timestamp 0
transform 1 0 11205 0 1 2557
box -211 -2169 211 2169
use sky130_fd_pr__pfet_01v8_MSU6BZ  XM2
timestamp 0
transform 1 0 15813 0 1 570
box -211 -288 211 288
use sky130_fd_pr__nfet_01v8_DJ4NP4  XM3
timestamp 0
transform 1 0 13509 0 1 587
box -2146 -252 2146 252
use sky130_fd_pr__pfet_01v8_KVC9YE  XM7
timestamp 0
transform 1 0 2643 0 1 808
box -2696 -261 2696 261
use sky130_fd_pr__pfet_01v8_KVC9YE  XM9
timestamp 0
transform 1 0 7982 0 1 755
box -2696 -261 2696 261
use sky130_fd_pr__nfet_01v8_3STNDZ  XM10
timestamp 0
transform 1 0 10836 0 1 3151
box -211 -2710 211 2710
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
