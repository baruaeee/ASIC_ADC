* NGSPICE file created from analog_therm.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_JLSX9N a_n317_n216# a_n157_n130# a_n215_n42# a_157_n42#
X0 a_157_n42# a_n157_n130# a_n215_n42# a_n317_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.57
C0 a_n157_n130# a_157_n42# 0.0179f
C1 a_n215_n42# a_157_n42# 0.0166f
C2 a_n215_n42# a_n157_n130# 0.0179f
C3 a_157_n42# a_n317_n216# 0.0832f
C4 a_n215_n42# a_n317_n216# 0.0832f
C5 a_n157_n130# a_n317_n216# 1.03f
.ends

.subckt sky130_fd_pr__pfet_01v8_XYZSMQ a_n33_n255# a_15_n158# w_n211_n377# a_n73_n158#
+ VSUBS
X0 a_15_n158# a_n33_n255# a_n73_n158# w_n211_n377# sky130_fd_pr__pfet_01v8 ad=0.458 pd=3.74 as=0.458 ps=3.74 w=1.58 l=0.15
C0 w_n211_n377# a_n33_n255# 0.24f
C1 a_15_n158# a_n33_n255# 0.0271f
C2 w_n211_n377# a_n73_n158# 0.117f
C3 a_15_n158# a_n73_n158# 0.254f
C4 a_15_n158# w_n211_n377# 0.117f
C5 a_n33_n255# a_n73_n158# 0.0271f
C6 a_15_n158# VSUBS 0.0732f
C7 a_n73_n158# VSUBS 0.0732f
C8 a_n33_n255# VSUBS 0.118f
C9 w_n211_n377# VSUBS 1.43f
.ends

.subckt sky130_fd_pr__pfet_01v8_AZD9DW w_n353_n261# a_n157_n139# a_n215_n42# a_157_n42#
+ VSUBS
X0 a_157_n42# a_n157_n139# a_n215_n42# w_n353_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.57
C0 w_n353_n261# a_n157_n139# 0.611f
C1 a_157_n42# a_n157_n139# 0.0179f
C2 w_n353_n261# a_n215_n42# 0.0498f
C3 a_157_n42# a_n215_n42# 0.0166f
C4 a_157_n42# w_n353_n261# 0.0498f
C5 a_n157_n139# a_n215_n42# 0.0179f
C6 a_157_n42# VSUBS 0.0329f
C7 a_n215_n42# VSUBS 0.0329f
C8 a_n157_n139# VSUBS 0.446f
C9 w_n353_n261# VSUBS 1.62f
.ends

.subckt sky130_fd_pr__nfet_01v8_T8HSQ7 a_15_n157# a_n175_n331# a_n33_n245# a_n73_n157#
X0 a_15_n157# a_n33_n245# a_n73_n157# a_n175_n331# sky130_fd_pr__nfet_01v8 ad=0.455 pd=3.72 as=0.455 ps=3.72 w=1.57 l=0.15
C0 a_n33_n245# a_n73_n157# 0.0289f
C1 a_n33_n245# a_15_n157# 0.0289f
C2 a_n73_n157# a_15_n157# 0.253f
C3 a_15_n157# a_n175_n331# 0.19f
C4 a_n73_n157# a_n175_n331# 0.19f
C5 a_n33_n245# a_n175_n331# 0.346f
.ends

.subckt th09 V09 Vin m1_891_n977# Vp m1_1725_85# Vn
XXM0 Vn Vin Vn m1_891_n977# sky130_fd_pr__nfet_01v8_JLSX9N
XXM1 Vin Vp Vp m1_891_n977# Vn sky130_fd_pr__pfet_01v8_XYZSMQ
XXM2 Vp m1_891_n977# Vp m1_1725_85# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM3 Vp m1_891_n977# V09 m1_1725_85# Vn sky130_fd_pr__pfet_01v8_AZD9DW
XXM4 V09 Vn m1_891_n977# Vn sky130_fd_pr__nfet_01v8_T8HSQ7
C0 m1_891_n977# Vp 0.469f
C1 m1_891_n977# m1_1725_85# 0.0672f
C2 m1_891_n977# V09 0.291f
C3 Vin Vp 0.162f
C4 Vin m1_1725_85# 9.1e-19
C5 Vin V09 0.00135f
C6 Vp m1_1725_85# 0.14f
C7 Vp V09 0.131f
C8 V09 m1_1725_85# 0.0153f
C9 Vin m1_891_n977# 0.208f
C10 Vin Vn 1.36f
C11 m1_891_n977# Vn 1.29f
C12 V09 Vn 0.467f
C13 Vp Vn 4.41f
C14 m1_1725_85# Vn 0.13f
.ends

.subckt sky130_fd_pr__pfet_01v8_FP437E w_n521_n261# a_n383_n42# a_n325_n139# a_325_n42#
+ VSUBS
X0 a_325_n42# a_n325_n139# a_n383_n42# w_n521_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=3.25
C0 a_n325_n139# w_n521_n261# 1.13f
C1 a_n325_n139# a_n383_n42# 0.0222f
C2 a_325_n42# a_n325_n139# 0.0222f
C3 a_n383_n42# w_n521_n261# 0.0498f
C4 a_325_n42# w_n521_n261# 0.0498f
C5 a_325_n42# a_n383_n42# 0.00865f
C6 a_325_n42# VSUBS 0.0355f
C7 a_n383_n42# VSUBS 0.0355f
C8 a_n325_n139# VSUBS 0.87f
C9 w_n521_n261# VSUBS 2.3f
.ends

.subckt sky130_fd_pr__nfet_01v8_L7T3GD a_n33_n130# a_15_n42# a_n175_n216# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n42# a_n33_n130# 0.0209f
C1 a_n73_n42# a_15_n42# 0.0699f
C2 a_15_n42# a_n33_n130# 0.0209f
C3 a_15_n42# a_n175_n216# 0.0729f
C4 a_n73_n42# a_n175_n216# 0.0729f
C5 a_n33_n130# a_n175_n216# 0.338f
.ends

.subckt preamp Vp Vin Vn Vpamp
XXM0 Vpamp Vpamp Vin Vn Vpamp sky130_fd_pr__pfet_01v8_FP437E
XXM1 Vin Vpamp Vpamp Vp sky130_fd_pr__nfet_01v8_L7T3GD
C0 Vin Vn 0.0405f
C1 Vn Vpamp 0.0667f
C2 Vin Vp 0.116f
C3 Vin Vpamp 0.665f
C4 Vpamp Vp 0.116f
C5 Vin 0 1.35f
C6 Vpamp 0 2.29f
C7 Vp 0 0.324f
C8 Vn 0 0.123f
.ends

.subckt sky130_fd_pr__pfet_01v8_3QB9EZ a_n296_n139# a_n354_n42# a_296_n42# w_n492_n261#
+ VSUBS
X0 a_296_n42# a_n296_n139# a_n354_n42# w_n492_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.96
C0 a_n296_n139# w_n492_n261# 1.04f
C1 a_n296_n139# a_296_n42# 0.0218f
C2 w_n492_n261# a_296_n42# 0.0498f
C3 a_n296_n139# a_n354_n42# 0.0218f
C4 w_n492_n261# a_n354_n42# 0.0498f
C5 a_296_n42# a_n354_n42# 0.00943f
C6 a_296_n42# VSUBS 0.0352f
C7 a_n354_n42# VSUBS 0.0352f
C8 a_n296_n139# VSUBS 0.797f
C9 w_n492_n261# VSUBS 2.19f
.ends

.subckt sky130_fd_pr__nfet_01v8_J2SMPG a_n33_n398# a_15_n310# a_n175_n484# a_n73_n310#
X0 a_15_n310# a_n33_n398# a_n73_n310# a_n175_n484# sky130_fd_pr__nfet_01v8 ad=0.899 pd=6.78 as=0.899 ps=6.78 w=3.1 l=0.15
C0 a_n73_n310# a_n33_n398# 0.0365f
C1 a_n73_n310# a_15_n310# 0.496f
C2 a_n33_n398# a_15_n310# 0.0365f
C3 a_15_n310# a_n175_n484# 0.345f
C4 a_n73_n310# a_n175_n484# 0.345f
C5 a_n33_n398# a_n175_n484# 0.349f
.ends

.subckt sky130_fd_pr__nfet_01v8_G45C34 a_297_n48# a_n297_n136# a_n457_n222# a_n355_n48#
X0 a_297_n48# a_n297_n136# a_n355_n48# a_n457_n222# sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.54 as=0.139 ps=1.54 w=0.48 l=2.97
C0 a_n355_n48# a_n297_n136# 0.0239f
C1 a_n355_n48# a_297_n48# 0.0107f
C2 a_n297_n136# a_297_n48# 0.0239f
C3 a_297_n48# a_n457_n222# 0.0929f
C4 a_n355_n48# a_n457_n222# 0.0929f
C5 a_n297_n136# a_n457_n222# 1.8f
.ends

.subckt sky130_fd_pr__pfet_01v8_XA2NHL a_15_n310# w_n211_n529# a_n73_n310# a_n33_n407#
+ VSUBS
X0 a_15_n310# a_n33_n407# a_n73_n310# w_n211_n529# sky130_fd_pr__pfet_01v8 ad=0.899 pd=6.78 as=0.899 ps=6.78 w=3.1 l=0.15
C0 w_n211_n529# a_n73_n310# 0.21f
C1 a_15_n310# a_n73_n310# 0.496f
C2 a_n73_n310# a_n33_n407# 0.0346f
C3 w_n211_n529# a_15_n310# 0.21f
C4 w_n211_n529# a_n33_n407# 0.241f
C5 a_15_n310# a_n33_n407# 0.0346f
C6 a_15_n310# VSUBS 0.135f
C7 a_n73_n310# VSUBS 0.135f
C8 a_n33_n407# VSUBS 0.121f
C9 w_n211_n529# VSUBS 1.97f
.ends

.subckt th01 Vp Vin Vout m1_931_n929# Vn
XXM2 Vin Vp m1_931_n929# Vp Vn sky130_fd_pr__pfet_01v8_3QB9EZ
XXM3 Vin m1_931_n929# Vn Vn sky130_fd_pr__nfet_01v8_J2SMPG
XXM4 Vn m1_931_n929# Vn Vout sky130_fd_pr__nfet_01v8_G45C34
XXM5 Vp Vp Vout m1_931_n929# Vn sky130_fd_pr__pfet_01v8_XA2NHL
C0 m1_931_n929# Vp 0.324f
C1 Vin m1_931_n929# 0.206f
C2 Vp Vout 0.0877f
C3 Vin Vout 5.64e-20
C4 m1_931_n929# Vout 0.202f
C5 Vin Vp 0.391f
C6 Vin Vn 1.12f
C7 m1_931_n929# Vn 2.31f
C8 Vp Vn 4.35f
C9 Vout Vn 0.405f
.ends

.subckt sky130_fd_pr__pfet_01v8_NZD9V2 w_n243_n261# a_47_n42# a_n47_n139# a_n105_n42#
+ VSUBS
X0 a_47_n42# a_n47_n139# a_n105_n42# w_n243_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.47
C0 a_47_n42# a_n105_n42# 0.0406f
C1 a_n105_n42# a_n47_n139# 0.00866f
C2 w_n243_n261# a_n105_n42# 0.0499f
C3 a_47_n42# a_n47_n139# 0.00866f
C4 a_47_n42# w_n243_n261# 0.0499f
C5 w_n243_n261# a_n47_n139# 0.27f
C6 a_47_n42# VSUBS 0.0297f
C7 a_n105_n42# VSUBS 0.0297f
C8 a_n47_n139# VSUBS 0.168f
C9 w_n243_n261# VSUBS 1.17f
.ends

.subckt sky130_fd_pr__pfet_01v8_3PDS9J a_n102_n42# a_44_n42# a_n44_n139# w_n240_n261#
+ VSUBS
X0 a_44_n42# a_n44_n139# a_n102_n42# w_n240_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.44
C0 a_44_n42# a_n102_n42# 0.0423f
C1 a_n102_n42# a_n44_n139# 0.00823f
C2 w_n240_n261# a_n102_n42# 0.0499f
C3 a_44_n42# a_n44_n139# 0.00823f
C4 a_44_n42# w_n240_n261# 0.0499f
C5 w_n240_n261# a_n44_n139# 0.261f
C6 a_44_n42# VSUBS 0.0296f
C7 a_n102_n42# VSUBS 0.0296f
C8 a_n44_n139# VSUBS 0.16f
C9 w_n240_n261# VSUBS 1.15f
.ends

.subckt sky130_fd_pr__nfet_01v8_97T34Z a_n73_n46# a_n175_n220# a_n33_n134# a_15_n46#
X0 a_15_n46# a_n33_n134# a_n73_n46# a_n175_n220# sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.5 as=0.133 ps=1.5 w=0.46 l=0.15
C0 a_15_n46# a_n73_n46# 0.0763f
C1 a_n33_n134# a_15_n46# 0.0212f
C2 a_n33_n134# a_n73_n46# 0.0212f
C3 a_15_n46# a_n175_n220# 0.0769f
C4 a_n73_n46# a_n175_n220# 0.0769f
C5 a_n33_n134# a_n175_n220# 0.338f
.ends

.subckt th06 Vp Vin V06 m1_528_n874# Vn
XXM0 Vin m1_528_n874# Vn Vn sky130_fd_pr__nfet_01v8_L7T3GD
XXM1 Vp m1_528_n874# Vin Vp Vn sky130_fd_pr__pfet_01v8_NZD9V2
XXM2 Vp V06 m1_528_n874# Vp Vn sky130_fd_pr__pfet_01v8_3PDS9J
XXM3 Vn Vn m1_528_n874# V06 sky130_fd_pr__nfet_01v8_97T34Z
C0 Vp V06 0.109f
C1 Vin m1_528_n874# 0.224f
C2 V06 Vin 2.39e-21
C3 V06 m1_528_n874# 0.135f
C4 Vp Vin 0.192f
C5 Vp m1_528_n874# 0.467f
C6 V06 Vn 0.353f
C7 m1_528_n874# Vn 0.971f
C8 Vin Vn 0.726f
C9 Vp Vn 2.62f
.ends

.subckt sky130_fd_pr__nfet_01v8_VGVEGU a_n74_n42# a_n33_n130# a_n176_n216# a_16_n42#
X0 a_16_n42# a_n33_n130# a_n74_n42# a_n176_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.16
C0 a_n33_n130# a_16_n42# 0.0191f
C1 a_16_n42# a_n74_n42# 0.0684f
C2 a_n33_n130# a_n74_n42# 0.0191f
C3 a_16_n42# a_n176_n216# 0.0737f
C4 a_n74_n42# a_n176_n216# 0.0737f
C5 a_n33_n130# a_n176_n216# 0.338f
.ends

.subckt sky130_fd_pr__pfet_01v8_EDPLE3 a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 w_n211_n261# a_n73_n42# 0.0463f
C1 a_15_n42# a_n33_n139# 0.0192f
C2 a_n73_n42# a_n33_n139# 0.0192f
C3 w_n211_n261# a_n33_n139# 0.236f
C4 a_15_n42# a_n73_n42# 0.0699f
C5 a_15_n42# w_n211_n261# 0.0463f
C6 a_15_n42# VSUBS 0.0263f
C7 a_n73_n42# VSUBS 0.0263f
C8 a_n33_n139# VSUBS 0.115f
C9 w_n211_n261# VSUBS 1.03f
.ends

.subckt th07 Vin V07 Vp m1_400_n1066# Vn
XXM0 m1_400_n1066# Vin Vn Vn sky130_fd_pr__nfet_01v8_VGVEGU
XXM1 m1_400_n1066# Vp Vin Vp Vn sky130_fd_pr__pfet_01v8_EDPLE3
XXM2 Vp V07 m1_400_n1066# Vp Vn sky130_fd_pr__pfet_01v8_NZD9V2
XXM3 Vn Vn m1_400_n1066# V07 sky130_fd_pr__nfet_01v8_97T34Z
C0 Vp V07 0.102f
C1 Vp m1_400_n1066# 0.32f
C2 m1_400_n1066# V07 0.167f
C3 Vin Vp 0.212f
C4 Vin V07 6.52e-19
C5 Vin m1_400_n1066# 0.436f
C6 Vin Vn 0.75f
C7 m1_400_n1066# Vn 0.943f
C8 V07 Vn 0.395f
C9 Vp Vn 2.43f
.ends

.subckt sky130_fd_pr__nfet_01v8_LNCAWD a_n67_n130# a_n125_n42# a_67_n42# a_n227_n216#
X0 a_67_n42# a_n67_n130# a_n125_n42# a_n227_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.67
C0 a_n67_n130# a_67_n42# 0.0112f
C1 a_n67_n130# a_n125_n42# 0.0112f
C2 a_67_n42# a_n125_n42# 0.0322f
C3 a_67_n42# a_n227_n216# 0.0807f
C4 a_n125_n42# a_n227_n216# 0.0807f
C5 a_n67_n130# a_n227_n216# 0.533f
.ends

.subckt sky130_fd_pr__pfet_01v8_M6KFPY a_n73_n67# a_n33_n164# a_15_n67# w_n211_n286#
+ VSUBS
X0 a_15_n67# a_n33_n164# a_n73_n67# w_n211_n286# sky130_fd_pr__pfet_01v8 ad=0.194 pd=1.92 as=0.194 ps=1.92 w=0.67 l=0.15
C0 a_15_n67# w_n211_n286# 0.0616f
C1 w_n211_n286# a_n73_n67# 0.0616f
C2 a_15_n67# a_n73_n67# 0.11f
C3 w_n211_n286# a_n33_n164# 0.238f
C4 a_15_n67# a_n33_n164# 0.0213f
C5 a_n73_n67# a_n33_n164# 0.0213f
C6 a_15_n67# VSUBS 0.0364f
C7 a_n73_n67# VSUBS 0.0364f
C8 a_n33_n164# VSUBS 0.116f
C9 w_n211_n286# VSUBS 1.11f
.ends

.subckt sky130_fd_pr__nfet_01v8_NCP4B2 a_n73_n47# a_n175_n221# a_n33_n135# a_15_n47#
X0 a_15_n47# a_n33_n135# a_n73_n47# a_n175_n221# sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.52 as=0.136 ps=1.52 w=0.47 l=0.15
C0 a_n33_n135# a_15_n47# 0.0213f
C1 a_n33_n135# a_n73_n47# 0.0213f
C2 a_15_n47# a_n73_n47# 0.0779f
C3 a_15_n47# a_n175_n221# 0.0779f
C4 a_n73_n47# a_n175_n221# 0.0779f
C5 a_n33_n135# a_n175_n221# 0.338f
.ends

.subckt th08 V08 Vin m1_451_n1105# Vp Vn
XXM0 Vin m1_451_n1105# Vn Vn sky130_fd_pr__nfet_01v8_LNCAWD
XXM1 m1_451_n1105# Vin Vp Vp Vn sky130_fd_pr__pfet_01v8_M6KFPY
XXM2 Vp V08 m1_451_n1105# Vp Vn sky130_fd_pr__pfet_01v8_NZD9V2
XXM3 Vn Vn m1_451_n1105# V08 sky130_fd_pr__nfet_01v8_NCP4B2
C0 V08 Vp 0.0989f
C1 Vin m1_451_n1105# 0.365f
C2 m1_451_n1105# V08 0.175f
C3 Vin V08 2.59e-19
C4 m1_451_n1105# Vp 0.176f
C5 Vin Vp 0.125f
C6 m1_451_n1105# Vn 0.838f
C7 Vin Vn 0.981f
C8 V08 Vn 0.403f
C9 Vp Vn 2.37f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n73_n100# a_n33_n197# 0.0281f
C1 a_n73_n100# a_15_n100# 0.162f
C2 a_15_n100# a_n33_n197# 0.0262f
C3 a_n73_n100# w_n211_n319# 0.0813f
C4 a_n33_n197# w_n211_n319# 0.246f
C5 a_15_n100# w_n211_n319# 0.0815f
C6 a_15_n100# VSUBS 0.0492f
C7 a_n73_n100# VSUBS 0.0487f
C8 a_n33_n197# VSUBS 0.129f
C9 w_n211_n319# VSUBS 1.23f
.ends

.subckt sky130_fd_pr__pfet_01v8_QPDSQG a_n87_n42# w_n225_n261# a_n33_n139# a_29_n42#
+ VSUBS
X0 a_29_n42# a_n33_n139# a_n87_n42# w_n225_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.29
C0 a_n87_n42# a_n33_n139# 0.00625f
C1 a_n87_n42# a_29_n42# 0.0532f
C2 a_29_n42# a_n33_n139# 0.00625f
C3 a_n87_n42# w_n225_n261# 0.0499f
C4 a_n33_n139# w_n225_n261# 0.229f
C5 a_29_n42# w_n225_n261# 0.0499f
C6 a_29_n42# VSUBS 0.029f
C7 a_n87_n42# VSUBS 0.029f
C8 a_n33_n139# VSUBS 0.128f
C9 w_n225_n261# VSUBS 1.09f
.ends

.subckt sky130_fd_pr__pfet_01v8_M479BZ a_15_n42# w_n211_n261# a_n33_n139# a_n73_n42#
+ VSUBS
X0 a_15_n42# a_n33_n139# a_n73_n42# w_n211_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n73_n42# a_n33_n139# 0.0192f
C1 a_n73_n42# a_15_n42# 0.0699f
C2 a_15_n42# a_n33_n139# 0.0192f
C3 a_n73_n42# w_n211_n261# 0.0463f
C4 a_n33_n139# w_n211_n261# 0.236f
C5 a_15_n42# w_n211_n261# 0.0463f
C6 a_15_n42# VSUBS 0.0263f
C7 a_n73_n42# VSUBS 0.0263f
C8 a_n33_n139# VSUBS 0.115f
C9 w_n211_n261# VSUBS 1.03f
.ends

.subckt th10 V10 Vin m1_718_n418# Vp Vn m1_878_n414#
XXM0 Vn m1_878_n414# Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Vin m1_878_n414# Vn m1_718_n418# sky130_fd_pr__nfet_01v8_L7T3GD
XXM2 Vp Vp Vin m1_718_n418# Vn sky130_fd_pr__pfet_01v8_QPDSQG
XXM3 V10 Vp m1_718_n418# Vp Vn sky130_fd_pr__pfet_01v8_M479BZ
XXM4 m1_718_n418# V10 Vn Vn sky130_fd_pr__nfet_01v8_L7T3GD
C0 m1_878_n414# V10 9.3e-21
C1 Vn Vp 0.468f
C2 Vin V10 1.33e-19
C3 Vn m1_718_n418# 0.14f
C4 m1_878_n414# Vp 0.0409f
C5 m1_878_n414# m1_718_n418# 0.0145f
C6 Vin Vp 0.301f
C7 Vn m1_878_n414# 0.157f
C8 Vin m1_718_n418# 0.308f
C9 Vp V10 0.0825f
C10 Vn Vin 0.0481f
C11 m1_718_n418# V10 0.191f
C12 Vn V10 0.0667f
C13 Vin m1_878_n414# 0.0391f
C14 Vp m1_718_n418# 0.272f
C15 Vin 0 0.692f
C16 m1_718_n418# 0 0.567f
C17 V10 0 0.319f
C18 Vn 0 0.208f
C19 Vp 0 3.6f
C20 m1_878_n414# 0 0.16f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGAKDL a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
+ VSUBS
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n33_n297# a_15_n200# 0.0293f
C1 a_15_n200# w_n211_n419# 0.143f
C2 a_n73_n200# a_15_n200# 0.321f
C3 a_n33_n297# w_n211_n419# 0.24f
C4 a_n33_n297# a_n73_n200# 0.0293f
C5 a_n73_n200# w_n211_n419# 0.143f
C6 a_15_n200# VSUBS 0.0902f
C7 a_n73_n200# VSUBS 0.0902f
C8 a_n33_n297# VSUBS 0.119f
C9 w_n211_n419# VSUBS 1.58f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFH27D a_50_n42# a_n210_n216# a_n108_n42# a_n50_n130#
X0 a_50_n42# a_n50_n130# a_n108_n42# a_n210_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 a_n108_n42# a_n50_n130# 0.00909f
C1 a_n108_n42# a_50_n42# 0.0391f
C2 a_50_n42# a_n50_n130# 0.00909f
C3 a_50_n42# a_n210_n216# 0.0801f
C4 a_n108_n42# a_n210_n216# 0.0801f
C5 a_n50_n130# a_n210_n216# 0.439f
.ends

.subckt sky130_fd_pr__pfet_01v8_E7ZT25 a_15_n43# w_n211_n262# a_n73_n43# a_n33_n140#
+ VSUBS
X0 a_15_n43# a_n33_n140# a_n73_n43# w_n211_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.15
C0 a_n33_n140# a_15_n43# 0.0193f
C1 a_15_n43# w_n211_n262# 0.0469f
C2 a_n73_n43# a_15_n43# 0.0715f
C3 a_n33_n140# w_n211_n262# 0.236f
C4 a_n33_n140# a_n73_n43# 0.0193f
C5 a_n73_n43# w_n211_n262# 0.0469f
C6 a_15_n43# VSUBS 0.0267f
C7 a_n73_n43# VSUBS 0.0267f
C8 a_n33_n140# VSUBS 0.115f
C9 w_n211_n262# VSUBS 1.03f
.ends

.subckt sky130_fd_pr__pfet_01v8_JM8GTH a_50_n42# w_n246_n261# a_n50_n139# a_n108_n42#
+ VSUBS
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 a_n50_n139# a_50_n42# 0.00909f
C1 a_50_n42# w_n246_n261# 0.0499f
C2 a_n108_n42# a_50_n42# 0.0391f
C3 a_n50_n139# w_n246_n261# 0.279f
C4 a_n50_n139# a_n108_n42# 0.00909f
C5 a_n108_n42# w_n246_n261# 0.0499f
C6 a_50_n42# VSUBS 0.0298f
C7 a_n108_n42# VSUBS 0.0298f
C8 a_n50_n139# VSUBS 0.175f
C9 w_n246_n261# VSUBS 1.18f
.ends

.subckt sky130_fd_pr__nfet_01v8_L9ESAD a_n175_n224# a_n73_n50# a_n33_n138# a_15_n50#
X0 a_15_n50# a_n33_n138# a_n73_n50# a_n175_n224# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_n73_n50# a_n33_n138# 0.0216f
C1 a_n73_n50# a_15_n50# 0.0826f
C2 a_15_n50# a_n33_n138# 0.0216f
C3 a_15_n50# a_n175_n224# 0.081f
C4 a_n73_n50# a_n175_n224# 0.081f
C5 a_n33_n138# a_n175_n224# 0.339f
.ends

.subckt th11 V11 Vin Vp m1_717_301# m1_509_303# Vn
XXM0 m1_717_301# Vp Vn Vn Vn sky130_fd_pr__pfet_01v8_XGAKDL
XXM1 m1_717_301# Vn m1_509_303# Vin sky130_fd_pr__nfet_01v8_ZFH27D
XXM2 m1_509_303# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_E7ZT25
XXM3 V11 Vp m1_509_303# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM4 Vn Vn m1_509_303# V11 sky130_fd_pr__nfet_01v8_L9ESAD
C0 Vin Vp 0.258f
C1 m1_717_301# Vp 0.0487f
C2 Vin m1_509_303# 0.248f
C3 m1_509_303# m1_717_301# 0.0301f
C4 V11 Vp 0.0686f
C5 Vin m1_717_301# 0.0345f
C6 m1_509_303# V11 0.0742f
C7 Vin V11 0.00112f
C8 m1_717_301# V11 1.71e-20
C9 m1_509_303# Vp 0.352f
C10 Vin Vn 0.856f
C11 m1_509_303# Vn 0.717f
C12 V11 Vn 0.485f
C13 Vp Vn 4.47f
C14 m1_717_301# Vn 0.299f
.ends

.subckt sky130_fd_pr__pfet_01v8_P28Q2U a_n33_n232# a_15_n135# w_n211_n354# a_n73_n135#
+ VSUBS
X0 a_15_n135# a_n33_n232# a_n73_n135# w_n211_n354# sky130_fd_pr__pfet_01v8 ad=0.391 pd=3.28 as=0.391 ps=3.28 w=1.35 l=0.15
C0 a_15_n135# a_n33_n232# 0.0258f
C1 a_n73_n135# a_n33_n232# 0.0258f
C2 a_15_n135# w_n211_n354# 0.103f
C3 w_n211_n354# a_n73_n135# 0.103f
C4 w_n211_n354# a_n33_n232# 0.24f
C5 a_15_n135# a_n73_n135# 0.218f
C6 a_15_n135# VSUBS 0.0639f
C7 a_n73_n135# VSUBS 0.0639f
C8 a_n33_n232# VSUBS 0.118f
C9 w_n211_n354# VSUBS 1.35f
.ends

.subckt sky130_fd_pr__nfet_01v8_HZA4VB a_n360_n216# a_n200_n130# a_200_n42# a_n258_n42#
X0 a_200_n42# a_n200_n130# a_n258_n42# a_n360_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_200_n42# a_n258_n42# 0.0134f
C1 a_n200_n130# a_200_n42# 0.0196f
C2 a_n200_n130# a_n258_n42# 0.0196f
C3 a_200_n42# a_n360_n216# 0.0841f
C4 a_n258_n42# a_n360_n216# 0.0841f
C5 a_n200_n130# a_n360_n216# 1.26f
.ends

.subckt sky130_fd_pr__pfet_01v8_WV9GCW a_n158_n42# w_n296_n261# a_n100_n139# a_100_n42#
+ VSUBS
X0 a_100_n42# a_n100_n139# a_n158_n42# w_n296_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1
C0 a_100_n42# a_n100_n139# 0.0144f
C1 a_n158_n42# a_n100_n139# 0.0144f
C2 a_100_n42# w_n296_n261# 0.0499f
C3 w_n296_n261# a_n158_n42# 0.0499f
C4 w_n296_n261# a_n100_n139# 0.434f
C5 a_100_n42# a_n158_n42# 0.024f
C6 a_100_n42# VSUBS 0.0315f
C7 a_n158_n42# VSUBS 0.0315f
C8 a_n100_n139# VSUBS 0.302f
C9 w_n296_n261# VSUBS 1.38f
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_15_n100# a_n73_n100# 0.162f
C1 a_n33_n188# a_15_n100# 0.0254f
C2 a_n33_n188# a_n73_n100# 0.0254f
C3 a_15_n100# a_n175_n274# 0.132f
C4 a_n73_n100# a_n175_n274# 0.132f
C5 a_n33_n188# a_n175_n274# 0.343f
.ends

.subckt th12 Vout Vin m1_532_n361# Vp m1_773_n853# Vn
XXM0 Vn m1_773_n853# Vp Vn Vn sky130_fd_pr__pfet_01v8_P28Q2U
XXM1 Vn Vin m1_773_n853# m1_532_n361# sky130_fd_pr__nfet_01v8_HZA4VB
XXM2 m1_532_n361# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM3 Vp Vp m1_532_n361# Vout Vn sky130_fd_pr__pfet_01v8_WV9GCW
XXM4 Vn m1_532_n361# Vout Vn sky130_fd_pr__nfet_01v8_648S5X
C0 Vin Vp 0.435f
C1 Vout Vin 4.83e-19
C2 m1_773_n853# Vin 0.102f
C3 m1_532_n361# Vin 0.399f
C4 Vout Vp 0.0968f
C5 m1_773_n853# Vp 0.0827f
C6 Vout m1_773_n853# 0.00284f
C7 m1_532_n361# Vp 0.226f
C8 Vout m1_532_n361# 0.181f
C9 m1_773_n853# m1_532_n361# 0.0208f
C10 m1_532_n361# Vn 1.04f
C11 Vout Vn 0.478f
C12 Vp Vn 4.59f
C13 Vin Vn 1.62f
C14 m1_773_n853# Vn 0.44f
.ends

.subckt sky130_fd_pr__nfet_01v8_L6G859 a_n288_n42# a_230_n42# a_n390_n216# a_n230_n130#
X0 a_230_n42# a_n230_n130# a_n288_n42# a_n390_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2.3
C0 a_n230_n130# a_230_n42# 0.0204f
C1 a_n230_n130# a_n288_n42# 0.0204f
C2 a_230_n42# a_n288_n42# 0.0119f
C3 a_230_n42# a_n390_n216# 0.0846f
C4 a_n288_n42# a_n390_n216# 0.0846f
C5 a_n230_n130# a_n390_n216# 1.43f
.ends

.subckt sky130_fd_pr__pfet_01v8_XW9KDL a_n73_n230# a_n33_n327# a_15_n230# w_n211_n449#
+ VSUBS
X0 a_15_n230# a_n33_n327# a_n73_n230# w_n211_n449# sky130_fd_pr__pfet_01v8 ad=0.667 pd=5.18 as=0.667 ps=5.18 w=2.3 l=0.15
C0 a_n73_n230# a_15_n230# 0.369f
C1 w_n211_n449# a_n73_n230# 0.161f
C2 a_n33_n327# a_15_n230# 0.0338f
C3 w_n211_n449# a_n33_n327# 0.246f
C4 w_n211_n449# a_15_n230# 0.161f
C5 a_n73_n230# a_n33_n327# 0.0338f
C6 a_15_n230# VSUBS 0.102f
C7 a_n73_n230# VSUBS 0.102f
C8 a_n33_n327# VSUBS 0.129f
C9 w_n211_n449# VSUBS 1.69f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GC6 a_200_n42# w_n396_n261# a_n200_n139# a_n258_n42#
+ VSUBS
X0 a_200_n42# a_n200_n139# a_n258_n42# w_n396_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=2
C0 a_n258_n42# a_200_n42# 0.0134f
C1 w_n396_n261# a_n258_n42# 0.0498f
C2 a_n200_n139# a_200_n42# 0.0196f
C3 w_n396_n261# a_n200_n139# 0.743f
C4 w_n396_n261# a_200_n42# 0.0498f
C5 a_n258_n42# a_n200_n139# 0.0196f
C6 a_200_n42# VSUBS 0.0338f
C7 a_n258_n42# VSUBS 0.0338f
C8 a_n200_n139# VSUBS 0.554f
C9 w_n396_n261# VSUBS 1.79f
.ends

.subckt sky130_fd_pr__nfet_01v8_ATLS57 a_15_n200# a_n175_n374# a_n73_n200# a_n33_n288#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n175_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n33_n288# a_15_n200# 0.0357f
C1 a_n33_n288# a_n73_n200# 0.0336f
C2 a_15_n200# a_n73_n200# 0.321f
C3 a_15_n200# a_n175_n374# 0.232f
C4 a_n73_n200# a_n175_n374# 0.232f
C5 a_n33_n288# a_n175_n374# 0.358f
.ends

.subckt th13 Vout Vin m1_724_n958# m1_546_n454# Vp Vn
XXM0 m1_724_n958# Vn Vp Vn Vn sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 m1_546_n454# m1_724_n958# Vn Vin sky130_fd_pr__nfet_01v8_L6G859
XXM2 m1_546_n454# Vin Vp Vp Vn sky130_fd_pr__pfet_01v8_XW9KDL
XXM3 Vout Vp m1_546_n454# Vp Vn sky130_fd_pr__pfet_01v8_VZ9GC6
XXM4 Vout Vn Vn m1_546_n454# sky130_fd_pr__nfet_01v8_ATLS57
C0 m1_724_n958# Vin 0.14f
C1 Vin Vn 0.126f
C2 m1_724_n958# Vout 0.00247f
C3 m1_724_n958# Vp 0.312f
C4 Vout Vn 0.147f
C5 Vp Vn 0.589f
C6 m1_724_n958# m1_546_n454# 0.0214f
C7 m1_546_n454# Vn 0.331f
C8 Vout Vin 0.00172f
C9 Vp Vin 0.151f
C10 m1_546_n454# Vin 0.349f
C11 Vp Vout 0.346f
C12 m1_724_n958# Vn 0.0967f
C13 m1_546_n454# Vout 0.546f
C14 m1_546_n454# Vp 0.574f
C15 Vout 0 0.513f
C16 Vn 0 0.573f
C17 m1_546_n454# 0 1.54f
C18 Vp 0 4.74f
C19 Vin 0 1.66f
C20 m1_724_n958# 0 0.188f
.ends

.subckt sky130_fd_pr__nfet_01v8_9GNSAK a_n33_n550# a_n125_n550# a_n227_n724# a_63_n550#
+ a_n63_n576#
X0 a_63_n550# a_n63_n576# a_n33_n550# a_n227_n724# sky130_fd_pr__nfet_01v8 ad=1.71 pd=11.6 as=0.908 ps=5.83 w=5.5 l=0.15
X1 a_n33_n550# a_n63_n576# a_n125_n550# a_n227_n724# sky130_fd_pr__nfet_01v8 ad=0.908 pd=5.83 as=1.71 ps=11.6 w=5.5 l=0.15
C0 a_63_n550# a_n33_n550# 0.809f
C1 a_n33_n550# a_n63_n576# 0.0599f
C2 a_63_n550# a_n63_n576# 0.0319f
C3 a_n125_n550# a_n33_n550# 0.809f
C4 a_n125_n550# a_n63_n576# 0.0232f
C5 a_63_n550# a_n227_n724# 0.596f
C6 a_n33_n550# a_n227_n724# 0.0778f
C7 a_n125_n550# a_n227_n724# 0.597f
C8 a_n63_n576# a_n227_n724# 0.3f
.ends

.subckt sky130_fd_pr__pfet_01v8_UTD9YE w_n1296_n261# a_n1158_n42# a_n1100_n139# a_1100_n42#
+ VSUBS
X0 a_1100_n42# a_n1100_n139# a_n1158_n42# w_n1296_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=11
C0 a_n1158_n42# w_n1296_n261# 0.0498f
C1 a_1100_n42# w_n1296_n261# 0.0498f
C2 a_n1100_n139# a_n1158_n42# 0.0251f
C3 a_n1100_n139# a_1100_n42# 0.0251f
C4 a_n1100_n139# w_n1296_n261# 3.52f
C5 a_1100_n42# VSUBS 0.0428f
C6 a_n1158_n42# VSUBS 0.0428f
C7 a_n1100_n139# VSUBS 2.83f
C8 w_n1296_n261# VSUBS 5.47f
.ends

.subckt sky130_fd_pr__nfet_01v8_VZ7MP4 a_n1158_n42# a_n1260_n216# a_n1100_n130# a_1100_n42#
X0 a_1100_n42# a_n1100_n130# a_n1158_n42# a_n1260_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=11
C0 a_1100_n42# a_n1100_n130# 0.0251f
C1 a_n1158_n42# a_n1100_n130# 0.0251f
C2 a_1100_n42# a_n1260_n216# 0.0931f
C3 a_n1158_n42# a_n1260_n216# 0.0931f
C4 a_n1100_n130# a_n1260_n216# 6.21f
.ends

.subckt sky130_fd_pr__pfet_01v8_UGSTRG a_n33_n1197# a_n76_n1100# w_n214_n1319# a_18_n1100#
+ VSUBS
X0 a_18_n1100# a_n33_n1197# a_n76_n1100# w_n214_n1319# sky130_fd_pr__pfet_01v8 ad=3.19 pd=22.6 as=3.19 ps=22.6 w=11 l=0.18
C0 a_18_n1100# a_n76_n1100# 1.64f
C1 a_n76_n1100# w_n214_n1319# 0.693f
C2 a_18_n1100# w_n214_n1319# 0.693f
C3 a_n33_n1197# a_n76_n1100# 0.0705f
C4 a_n33_n1197# a_18_n1100# 0.0705f
C5 a_n33_n1197# w_n214_n1319# 0.239f
C6 a_18_n1100# VSUBS 0.46f
C7 a_n76_n1100# VSUBS 0.46f
C8 a_n33_n1197# VSUBS 0.133f
C9 w_n214_n1319# VSUBS 4.79f
.ends

.subckt th02 Vout Vn Vp m1_4146_502# Vin m1_1199_9#
XXM0 Vn m1_4146_502# Vn m1_4146_502# Vin sky130_fd_pr__nfet_01v8_9GNSAK
XXM1 Vp m1_1199_9# Vin m1_4146_502# Vn sky130_fd_pr__pfet_01v8_UTD9YE
XXM2 m1_1199_9# Vn Vp Vp sky130_fd_pr__nfet_01v8_VZ7MP4
XXM3 m1_4146_502# Vout Vp Vp Vn sky130_fd_pr__pfet_01v8_UGSTRG
XXM4 Vn Vn m1_4146_502# Vout sky130_fd_pr__nfet_01v8_VZ7MP4
C0 m1_1199_9# m1_4146_502# 4.98e-19
C1 Vin Vp 0.3f
C2 Vin Vout 0.0111f
C3 Vout Vp 0.202f
C4 Vin m1_4146_502# 0.58f
C5 Vp m1_4146_502# 0.374f
C6 Vout m1_4146_502# 0.328f
C7 m1_1199_9# Vin 0.0993f
C8 m1_1199_9# Vp 0.155f
C9 Vout Vn 0.554f
C10 m1_4146_502# Vn 9.06f
C11 m1_1199_9# Vn 0.445f
C12 Vp Vn 16.7f
C13 Vin Vn 2.92f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJ7SDL a_15_n450# w_n211_n669# a_n73_n450# a_n33_n547#
+ VSUBS
X0 a_15_n450# a_n33_n547# a_n73_n450# w_n211_n669# sky130_fd_pr__pfet_01v8 ad=1.3 pd=9.58 as=1.3 ps=9.58 w=4.5 l=0.15
C0 a_n73_n450# w_n211_n669# 0.295f
C1 a_n33_n547# a_15_n450# 0.0407f
C2 a_n73_n450# a_15_n450# 0.718f
C3 w_n211_n669# a_15_n450# 0.295f
C4 a_n73_n450# a_n33_n547# 0.0407f
C5 w_n211_n669# a_n33_n547# 0.242f
C6 a_15_n450# VSUBS 0.191f
C7 a_n73_n450# VSUBS 0.191f
C8 a_n33_n547# VSUBS 0.122f
C9 w_n211_n669# VSUBS 2.46f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFMUVB a_n608_n42# a_550_n42# a_n710_n216# a_n550_n130#
X0 a_550_n42# a_n550_n130# a_n608_n42# a_n710_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=5.5
C0 a_550_n42# a_n550_n130# 0.0242f
C1 a_550_n42# a_n608_n42# 0.00526f
C2 a_n550_n130# a_n608_n42# 0.0242f
C3 a_550_n42# a_n710_n216# 0.0873f
C4 a_n608_n42# a_n710_n216# 0.0873f
C5 a_n550_n130# a_n710_n216# 3.19f
.ends

.subckt sky130_fd_pr__pfet_01v8_UJPVTG w_n211_n769# a_n73_n550# a_n33_n647# a_15_n550#
+ VSUBS
X0 a_15_n550# a_n33_n647# a_n73_n550# w_n211_n769# sky130_fd_pr__pfet_01v8 ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.15
C0 a_n73_n550# w_n211_n769# 0.356f
C1 a_n33_n647# a_15_n550# 0.0449f
C2 a_n73_n550# a_15_n550# 0.877f
C3 w_n211_n769# a_15_n550# 0.356f
C4 a_n73_n550# a_n33_n647# 0.0449f
C5 w_n211_n769# a_n33_n647# 0.242f
C6 a_15_n550# VSUBS 0.232f
C7 a_n73_n550# VSUBS 0.232f
C8 a_n33_n647# VSUBS 0.122f
C9 w_n211_n769# VSUBS 2.81f
.ends

.subckt sky130_fd_pr__pfet_01v8_VZ9GTR a_n608_n42# a_550_n42# w_n746_n261# a_n550_n139#
+ VSUBS
X0 a_550_n42# a_n550_n139# a_n608_n42# w_n746_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=5.5
C0 a_n608_n42# w_n746_n261# 0.0498f
C1 a_n550_n139# a_550_n42# 0.0242f
C2 a_n608_n42# a_550_n42# 0.00526f
C3 w_n746_n261# a_550_n42# 0.0498f
C4 a_n608_n42# a_n550_n139# 0.0242f
C5 w_n746_n261# a_n550_n139# 1.82f
C6 a_550_n42# VSUBS 0.037f
C7 a_n608_n42# VSUBS 0.037f
C8 a_n550_n139# VSUBS 1.44f
C9 w_n746_n261# VSUBS 3.22f
.ends

.subckt sky130_fd_pr__nfet_01v8_9GNSAM a_n73_n550# a_n175_n724# a_15_n550# a_n33_n638#
X0 a_15_n550# a_n33_n638# a_n73_n550# a_n175_n724# sky130_fd_pr__nfet_01v8 ad=1.6 pd=11.6 as=1.6 ps=11.6 w=5.5 l=0.15
C0 a_15_n550# a_n33_n638# 0.0468f
C1 a_15_n550# a_n73_n550# 0.877f
C2 a_n33_n638# a_n73_n550# 0.0468f
C3 a_15_n550# a_n175_n724# 0.588f
C4 a_n73_n550# a_n175_n724# 0.588f
C5 a_n33_n638# a_n175_n724# 0.352f
.ends

.subckt th14 Vin m1_1594_n962# Vout Vp m1_710_n388# m1_2498_n384# Vn
XXM0 m1_1594_n962# Vp Vn Vn Vn sky130_fd_pr__pfet_01v8_XJ7SDL
XXM1 m1_710_n388# m1_1594_n962# Vn Vin sky130_fd_pr__nfet_01v8_ZFMUVB
XXM2 Vp m1_710_n388# Vin Vp Vn sky130_fd_pr__pfet_01v8_UJPVTG
XXM3 Vp m1_2498_n384# Vp m1_710_n388# Vn sky130_fd_pr__pfet_01v8_VZ9GTR
XXM4 m1_2498_n384# Vout Vp m1_710_n388# Vn sky130_fd_pr__pfet_01v8_VZ9GTR
XXM5 Vn Vn Vout m1_710_n388# sky130_fd_pr__nfet_01v8_9GNSAM
C0 m1_710_n388# Vn 0.459f
C1 Vn m1_2498_n384# 3.34e-24
C2 Vp m1_710_n388# 0.755f
C3 Vp m1_2498_n384# 0.276f
C4 m1_710_n388# Vout 0.191f
C5 Vout m1_2498_n384# 0.0142f
C6 Vp Vn 0.876f
C7 Vn Vout 0.0354f
C8 Vp Vout 0.125f
C9 m1_710_n388# m1_1594_n962# 0.00647f
C10 m1_710_n388# Vin 0.365f
C11 m1_2498_n384# Vin 1.46e-19
C12 Vn m1_1594_n962# 0.111f
C13 Vn Vin 0.0583f
C14 Vp m1_1594_n962# 0.237f
C15 Vp Vin 0.214f
C16 Vin m1_1594_n962# 0.166f
C17 m1_710_n388# m1_2498_n384# 0.768f
C18 Vin 0 3.4f
C19 Vout 0 0.854f
C20 Vn 0 0.831f
C21 m1_710_n388# 0 3.52f
C22 m1_2498_n384# 0 0.297f
C23 Vp 0 11.9f
C24 m1_1594_n962# 0 0.292f
.ends

.subckt sky130_fd_pr__nfet_01v8_8X7S4D a_15_n130# a_n33_n218# a_n73_n130# a_n175_n304#
X0 a_15_n130# a_n33_n218# a_n73_n130# a_n175_n304# sky130_fd_pr__nfet_01v8 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=0.15
C0 a_n73_n130# a_n33_n218# 0.0274f
C1 a_n73_n130# a_15_n130# 0.21f
C2 a_15_n130# a_n33_n218# 0.0274f
C3 a_15_n130# a_n175_n304# 0.162f
C4 a_n73_n130# a_n175_n304# 0.162f
C5 a_n33_n218# a_n175_n304# 0.345f
.ends

.subckt sky130_fd_pr__pfet_01v8_GZD9X3 a_n139_n139# a_139_n42# w_n335_n261# a_n197_n42#
+ VSUBS
X0 a_139_n42# a_n139_n139# a_n197_n42# w_n335_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.39
C0 a_n197_n42# a_139_n42# 0.0184f
C1 a_n139_n139# w_n335_n261# 0.555f
C2 a_n139_n139# a_n197_n42# 0.017f
C3 a_n197_n42# w_n335_n261# 0.0498f
C4 a_n139_n139# a_139_n42# 0.017f
C5 a_139_n42# w_n335_n261# 0.0498f
C6 a_139_n42# VSUBS 0.0325f
C7 a_n197_n42# VSUBS 0.0325f
C8 a_n139_n139# VSUBS 0.4f
C9 w_n335_n261# VSUBS 1.54f
.ends

.subckt sky130_fd_pr__nfet_01v8_LH5FDA a_n310_n216# a_n150_n130# a_n208_n42# a_150_n42#
X0 a_150_n42# a_n150_n130# a_n208_n42# a_n310_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.5
C0 a_n208_n42# a_n150_n130# 0.0176f
C1 a_n208_n42# a_150_n42# 0.0172f
C2 a_150_n42# a_n150_n130# 0.0176f
C3 a_150_n42# a_n310_n216# 0.0831f
C4 a_n208_n42# a_n310_n216# 0.0831f
C5 a_n150_n130# a_n310_n216# 0.99f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJP3BL a_15_n150# w_n211_n369# a_n73_n150# a_n33_n247#
+ VSUBS
X0 a_15_n150# a_n33_n247# a_n73_n150# w_n211_n369# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.15
C0 a_n73_n150# a_15_n150# 0.242f
C1 a_n33_n247# w_n211_n369# 0.24f
C2 a_n33_n247# a_n73_n150# 0.0267f
C3 a_n73_n150# w_n211_n369# 0.112f
C4 a_n33_n247# a_15_n150# 0.0267f
C5 a_15_n150# w_n211_n369# 0.112f
C6 a_15_n150# VSUBS 0.07f
C7 a_n73_n150# VSUBS 0.07f
C8 a_n33_n247# VSUBS 0.118f
C9 w_n211_n369# VSUBS 1.41f
.ends

.subckt th03 Vp Vout Vin m1_782_n682# Vn li_1010_10# m1_522_n210#
XXM0 m1_782_n682# Vin Vn Vn sky130_fd_pr__nfet_01v8_8X7S4D
XXM1 Vin m1_782_n682# li_1010_10# m1_522_n210# Vn sky130_fd_pr__pfet_01v8_GZD9X3
XXM2 Vn Vp m1_522_n210# Vp sky130_fd_pr__nfet_01v8_LH5FDA
XXM3 Vout li_1010_10# Vp m1_782_n682# Vn sky130_fd_pr__pfet_01v8_XJP3BL
XXM4 Vn m1_782_n682# Vn Vout sky130_fd_pr__nfet_01v8_LH5FDA
C0 m1_522_n210# Vp 0.041f
C1 li_1010_10# Vin 0.0791f
C2 Vin m1_782_n682# 0.212f
C3 Vout Vp 3.29e-19
C4 m1_522_n210# li_1010_10# 0.0635f
C5 m1_522_n210# m1_782_n682# 0.0254f
C6 m1_522_n210# Vin 0.0482f
C7 Vout li_1010_10# 0.132f
C8 li_1010_10# Vp 0.0961f
C9 Vout m1_782_n682# 0.0652f
C10 m1_782_n682# Vp 0.143f
C11 Vout Vin 5.05e-19
C12 Vin Vp 0.0439f
C13 m1_522_n210# Vout 0.00126f
C14 li_1010_10# m1_782_n682# 0.263f
C15 Vout Vn 0.462f
C16 m1_782_n682# Vn 1.57f
C17 Vp Vn 1.26f
C18 li_1010_10# Vn 3.06f
C19 m1_522_n210# Vn 0.278f
C20 Vin Vn 0.853f
.ends

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPB A3 0.0268f
C1 C1 VGND 0.0181f
C2 VPB a_75_199# 0.0486f
C3 A2 VGND 0.0119f
C4 A2 a_315_47# 0.00335f
C5 A1 VPB 0.0306f
C6 VPWR VPB 0.0749f
C7 A2 a_208_47# 0.00102f
C8 a_201_297# VPB 0.00186f
C9 X VPB 0.0107f
C10 a_75_199# A3 0.163f
C11 B1 VPB 0.0292f
C12 VPWR A3 0.0181f
C13 A1 a_75_199# 0.0696f
C14 VPWR a_75_199# 0.109f
C15 VGND VPB 0.00772f
C16 a_201_297# A3 0.00642f
C17 X A3 0.00317f
C18 a_201_297# a_75_199# 0.16f
C19 VPWR A1 0.0151f
C20 X a_75_199# 0.0959f
C21 a_201_297# A1 0.011f
C22 VPWR a_201_297# 0.211f
C23 A1 X 1.2e-19
C24 C1 VPB 0.0394f
C25 B1 a_75_199# 0.102f
C26 VPWR X 0.0676f
C27 A2 VPB 0.0376f
C28 VGND A3 0.0161f
C29 a_201_297# X 0.0131f
C30 B1 A1 0.0716f
C31 VPWR B1 0.0125f
C32 VGND a_75_199# 0.362f
C33 a_201_297# B1 0.00594f
C34 a_544_297# a_75_199# 0.0176f
C35 a_315_47# a_75_199# 0.0202f
C36 a_208_47# A3 3.65e-19
C37 B1 X 7.79e-20
C38 VGND A1 0.0113f
C39 VPWR VGND 0.0735f
C40 a_208_47# a_75_199# 0.0159f
C41 a_315_47# A1 0.00313f
C42 A2 A3 0.0747f
C43 VPWR a_544_297# 0.0105f
C44 VPWR a_315_47# 0.00154f
C45 a_201_297# VGND 0.00403f
C46 C1 a_75_199# 0.0628f
C47 A2 a_75_199# 0.0621f
C48 VGND X 0.0609f
C49 VPWR a_208_47# 8.35e-19
C50 a_201_297# a_544_297# 0.00702f
C51 a_544_297# X 2.35e-19
C52 C1 A1 3.21e-19
C53 A2 A1 0.0689f
C54 VPWR C1 0.0146f
C55 VPWR A2 0.0174f
C56 B1 VGND 0.0171f
C57 a_208_47# X 1.91e-19
C58 B1 a_544_297# 1.13e-19
C59 C1 a_201_297# 0.00243f
C60 A2 a_201_297# 0.0112f
C61 C1 X 5.14e-20
C62 A2 X 3.01e-19
C63 VGND a_544_297# 0.00256f
C64 VGND a_315_47# 0.00427f
C65 C1 B1 0.066f
C66 VGND a_208_47# 0.00302f
C67 VGND VNB 0.437f
C68 VPWR VNB 0.365f
C69 X VNB 0.0906f
C70 C1 VNB 0.148f
C71 B1 VNB 0.0947f
C72 A1 VNB 0.101f
C73 A2 VNB 0.11f
C74 A3 VNB 0.0908f
C75 VPB VNB 0.782f
C76 a_201_297# VNB 0.00345f
C77 a_75_199# VNB 0.205f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_181_47# C 0.00151f
C1 a_27_47# VPWR 0.145f
C2 VPWR C 0.00464f
C3 a_27_47# C 0.186f
C4 a_109_47# A 6.45e-19
C5 B A 0.0869f
C6 B X 0.00111f
C7 VGND A 0.0154f
C8 VPB A 0.0426f
C9 VGND X 0.0708f
C10 VPB X 0.0121f
C11 VGND a_109_47# 0.00123f
C12 B VGND 0.00714f
C13 B VPB 0.0836f
C14 VPWR A 0.0185f
C15 VGND VPB 0.00604f
C16 VPWR X 0.0766f
C17 VGND a_181_47# 0.00261f
C18 VPWR a_109_47# 3.29e-19
C19 B VPWR 0.128f
C20 a_27_47# A 0.157f
C21 VGND VPWR 0.0475f
C22 a_27_47# X 0.087f
C23 VPWR VPB 0.0795f
C24 X C 0.0149f
C25 a_27_47# a_109_47# 0.00517f
C26 B a_27_47# 0.0625f
C27 a_181_47# VPWR 3.97e-19
C28 B C 0.0746f
C29 a_27_47# VGND 0.134f
C30 a_27_47# VPB 0.0501f
C31 VGND C 0.0703f
C32 VPB C 0.0347f
C33 a_27_47# a_181_47# 0.00401f
C34 VGND VNB 0.3f
C35 X VNB 0.0923f
C36 C VNB 0.12f
C37 A VNB 0.174f
C38 VPWR VNB 0.274f
C39 B VNB 0.102f
C40 VPB VNB 0.516f
C41 a_27_47# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
C0 VGND VPB 0.0797f
C1 VPWR VPB 0.0625f
C2 VGND VPWR 0.353f
C3 VPWR VNB 0.47f
C4 VGND VNB 0.427f
C5 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VGND VPB 0.116f
C1 VPWR VPB 0.0787f
C2 VGND VPWR 0.546f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
C0 VPWR a_81_21# 0.146f
C1 VGND A1 0.0786f
C2 VPB B1 0.0387f
C3 A1 a_81_21# 0.0568f
C4 VGND B1 0.0181f
C5 VGND VPB 0.00713f
C6 B1 a_81_21# 0.148f
C7 VPB a_81_21# 0.0593f
C8 VGND a_81_21# 0.173f
C9 a_384_47# a_299_297# 1.48e-19
C10 A2 a_299_297# 0.0468f
C11 VPWR a_299_297# 0.202f
C12 A1 a_299_297# 0.0585f
C13 VPWR X 0.0847f
C14 a_384_47# VPWR 4.08e-19
C15 B1 a_299_297# 0.00863f
C16 VPB a_299_297# 0.0111f
C17 VPWR A2 0.0201f
C18 A1 a_384_47# 0.00884f
C19 B1 X 3.04e-20
C20 A1 A2 0.0921f
C21 VGND a_299_297# 0.00772f
C22 VPB X 0.0108f
C23 a_299_297# a_81_21# 0.0821f
C24 A1 VPWR 0.0209f
C25 VGND X 0.0512f
C26 X a_81_21# 0.112f
C27 VPB A2 0.0373f
C28 VPWR B1 0.0196f
C29 VGND a_384_47# 0.00366f
C30 VPWR VPB 0.068f
C31 VGND A2 0.0495f
C32 a_384_47# a_81_21# 0.00138f
C33 A1 B1 0.0817f
C34 A1 VPB 0.0264f
C35 A2 a_81_21# 7.47e-19
C36 VGND VPWR 0.0579f
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 A Y 0.0894f
C1 VPWR VGND 0.0423f
C2 VPB VGND 0.00649f
C3 Y VGND 0.155f
C4 VPWR VPB 0.0521f
C5 VPWR Y 0.209f
C6 A VGND 0.0638f
C7 VPWR A 0.0631f
C8 VPB Y 0.0061f
C9 A VPB 0.0742f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 a_111_297# A 0.00223f
C1 B VPWR 0.147f
C2 VPB A 0.0377f
C3 B X 6.52e-19
C4 B a_29_53# 0.121f
C5 a_183_297# A 0.00239f
C6 B VGND 0.0152f
C7 X VPWR 0.0885f
C8 B C 0.0802f
C9 a_29_53# VPWR 0.0833f
C10 a_29_53# X 0.0991f
C11 VGND VPWR 0.0459f
C12 B VPB 0.0962f
C13 VGND X 0.036f
C14 C VPWR 0.00457f
C15 a_111_297# VPWR 5.94e-19
C16 VGND a_29_53# 0.217f
C17 C a_29_53# 0.0857f
C18 VPB VPWR 0.0649f
C19 a_111_297# a_29_53# 0.005f
C20 VGND C 0.0161f
C21 B A 0.0787f
C22 VPB X 0.0109f
C23 VGND a_111_297# 3.96e-19
C24 VPB a_29_53# 0.0491f
C25 a_183_297# VPWR 8.13e-19
C26 VGND VPB 0.00724f
C27 VPWR A 0.00936f
C28 VPB C 0.0396f
C29 X A 0.00127f
C30 a_183_297# a_29_53# 0.00868f
C31 a_29_53# A 0.242f
C32 a_183_297# VGND 5.75e-19
C33 VGND A 0.0187f
C34 C A 0.0343f
C35 VGND VNB 0.306f
C36 X VNB 0.0882f
C37 A VNB 0.117f
C38 C VNB 0.16f
C39 B VNB 0.117f
C40 VPWR VNB 0.253f
C41 VPB VNB 0.516f
C42 a_29_53# VNB 0.18f
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
C0 VGND VPB 0.161f
C1 VPWR VPB 0.0858f
C2 VGND VPWR 0.903f
C3 VPWR VNB 0.867f
C4 VGND VNB 0.761f
C5 VPB VNB 0.605f
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 Y B 0.0877f
C1 A B 0.0584f
C2 A Y 0.0471f
C3 VPWR a_109_297# 0.00638f
C4 Y a_109_297# 0.0113f
C5 VPB VGND 0.00456f
C6 VPWR VPB 0.0449f
C7 VPWR VGND 0.0314f
C8 VPB B 0.0367f
C9 VPB Y 0.0139f
C10 VPB A 0.0415f
C11 VGND B 0.0451f
C12 Y VGND 0.154f
C13 A VGND 0.0486f
C14 VPWR B 0.0148f
C15 VPWR Y 0.0995f
C16 VGND a_109_297# 0.00128f
C17 VPWR A 0.0528f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
C0 X A2 0.00157f
C1 a_109_297# B2 0.0133f
C2 a_193_297# VGND 0.00438f
C3 VPWR A2 0.0209f
C4 VPWR X 0.0897f
C5 VGND B2 0.0174f
C6 a_193_297# A2 0.00683f
C7 a_193_297# X 0.00367f
C8 VPB B1 0.0321f
C9 a_193_297# VPWR 0.169f
C10 X B2 6.77e-20
C11 VPB a_27_47# 0.0512f
C12 VPWR B2 0.00842f
C13 VPB A1 0.0343f
C14 a_193_297# B2 0.00126f
C15 VPB C1 0.0367f
C16 VPB a_109_297# 0.00421f
C17 a_27_47# B1 0.112f
C18 VGND VPB 0.00844f
C19 A1 B1 0.0609f
C20 a_205_47# a_27_47# 0.00762f
C21 VPB A2 0.027f
C22 C1 B1 6.46e-19
C23 VPB X 0.0113f
C24 A1 a_27_47# 0.0984f
C25 VPB VPWR 0.0799f
C26 a_109_297# B1 0.00736f
C27 C1 a_27_47# 0.0792f
C28 a_193_297# VPB 0.00774f
C29 VGND B1 0.0133f
C30 a_109_297# a_27_47# 0.0961f
C31 A1 C1 1.77e-20
C32 VPB B2 0.0256f
C33 VGND a_27_47# 0.395f
C34 a_205_47# VGND 0.00156f
C35 A1 a_109_297# 1.05e-19
C36 X B1 9.58e-20
C37 a_465_47# a_27_47# 0.013f
C38 VPWR B1 0.00982f
C39 a_109_297# C1 0.00739f
C40 VGND A1 0.0126f
C41 A2 a_27_47# 0.153f
C42 X a_27_47# 0.0921f
C43 VGND C1 0.0196f
C44 A1 a_465_47# 7.06e-19
C45 a_193_297# B1 0.00869f
C46 VPWR a_27_47# 0.099f
C47 a_205_47# VPWR 1.62e-19
C48 A1 A2 0.0692f
C49 A1 X 2.77e-19
C50 B1 B2 0.0784f
C51 VGND a_109_297# 0.00284f
C52 a_193_297# a_27_47# 0.144f
C53 A1 VPWR 0.0161f
C54 C1 A2 9.03e-21
C55 X C1 5.03e-20
C56 a_27_47# B2 0.0959f
C57 VPWR C1 0.0139f
C58 a_109_297# X 3.99e-19
C59 a_193_297# A1 0.0109f
C60 VGND a_465_47# 0.00257f
C61 a_109_297# VPWR 0.15f
C62 VGND A2 0.0168f
C63 VGND X 0.061f
C64 C1 B2 0.0726f
C65 VGND VPWR 0.0722f
C66 a_465_47# X 1.56e-19
C67 a_193_297# a_109_297# 0.0927f
C68 a_465_47# VPWR 5.05e-19
C69 VGND VNB 0.437f
C70 X VNB 0.0919f
C71 VPWR VNB 0.364f
C72 A2 VNB 0.0896f
C73 A1 VNB 0.106f
C74 B1 VNB 0.108f
C75 B2 VNB 0.0887f
C76 C1 VNB 0.139f
C77 VPB VNB 0.782f
C78 a_193_297# VNB 0.0011f
C79 a_109_297# VNB 7.11e-19
C80 a_27_47# VNB 0.216f
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
C0 A2 a_93_21# 0.0747f
C1 A1 VPB 0.0296f
C2 A1 B2 3.14e-19
C3 VPB a_93_21# 0.0485f
C4 VPWR X 0.0849f
C5 A1 a_346_47# 0.00465f
C6 B2 a_93_21# 0.0147f
C7 A3 a_93_21# 0.124f
C8 VPWR a_250_297# 0.313f
C9 a_346_47# a_93_21# 0.0119f
C10 a_584_47# a_93_21# 0.00278f
C11 B1 VPWR 0.01f
C12 A1 a_93_21# 0.0641f
C13 VPWR a_256_47# 9.47e-19
C14 a_250_297# X 5.42e-19
C15 VPWR VGND 0.076f
C16 VPWR A2 0.0133f
C17 B1 X 3.83e-20
C18 B1 a_250_297# 0.0125f
C19 VPB VPWR 0.0756f
C20 VPWR B2 0.0108f
C21 VPWR A3 0.0158f
C22 VGND X 0.06f
C23 VPWR a_346_47# 0.00109f
C24 VGND a_250_297# 0.0072f
C25 A2 X 1.19e-19
C26 B1 a_256_47# 2.07e-20
C27 VPWR a_584_47# 9.47e-19
C28 A2 a_250_297# 0.0129f
C29 VPB X 0.0108f
C30 B1 VGND 0.0344f
C31 A1 VPWR 0.016f
C32 VPB a_250_297# 0.00616f
C33 X A3 2.45e-19
C34 B1 A2 1.44e-20
C35 a_256_47# VGND 0.00394f
C36 VPWR a_93_21# 0.0907f
C37 B2 a_250_297# 0.0344f
C38 a_250_297# A3 0.00602f
C39 B1 VPB 0.0276f
C40 a_256_47# A2 0.00256f
C41 B1 B2 0.0823f
C42 B1 A3 7.88e-22
C43 a_584_47# a_250_297# 2.43e-19
C44 A2 VGND 0.0114f
C45 A1 X 6.03e-20
C46 B1 a_346_47# 5.39e-20
C47 VPB VGND 0.00788f
C48 a_256_47# A3 4.42e-19
C49 A1 a_250_297# 0.0129f
C50 X a_93_21# 0.0841f
C51 B1 a_584_47# 0.00143f
C52 B2 VGND 0.0469f
C53 VGND A3 0.00974f
C54 a_250_297# a_93_21# 0.188f
C55 VPB A2 0.0287f
C56 B1 A1 0.0965f
C57 VGND a_346_47# 0.00514f
C58 A2 B2 1.46e-19
C59 A2 A3 0.0788f
C60 a_584_47# VGND 0.00683f
C61 B1 a_93_21# 0.0774f
C62 A2 a_346_47# 0.00252f
C63 VPB B2 0.0355f
C64 VPB A3 0.0291f
C65 A1 VGND 0.0133f
C66 a_256_47# a_93_21# 0.0114f
C67 B2 A3 9.12e-20
C68 VGND a_93_21# 0.251f
C69 A1 A2 0.0971f
C70 VGND VNB 0.465f
C71 VPWR VNB 0.365f
C72 X VNB 0.0937f
C73 B2 VNB 0.14f
C74 B1 VNB 0.101f
C75 A1 VNB 0.0951f
C76 A2 VNB 0.0921f
C77 A3 VNB 0.0929f
C78 VPB VNB 0.782f
C79 a_250_297# VNB 0.0278f
C80 a_93_21# VNB 0.151f
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 a_27_297# D 0.054f
C1 VGND X 0.0354f
C2 B D 0.00287f
C3 VPB C 0.0338f
C4 a_109_297# VGND 7.58e-19
C5 VGND D 0.0517f
C6 VPB A 0.033f
C7 VPB VPWR 0.075f
C8 VPB a_27_297# 0.0517f
C9 a_205_297# C 0.00261f
C10 A C 0.028f
C11 VPB B 0.106f
C12 VPB X 0.0109f
C13 VPWR C 0.00723f
C14 VPB VGND 0.00796f
C15 a_27_297# C 0.158f
C16 a_205_297# VPWR 5.16e-19
C17 a_205_297# a_27_297# 0.00412f
C18 A VPWR 0.00769f
C19 VPB D 0.0405f
C20 a_277_297# C 5.54e-19
C21 C B 0.0917f
C22 A a_27_297# 0.163f
C23 VGND C 0.0191f
C24 a_27_297# VPWR 0.084f
C25 A a_277_297# 2.28e-19
C26 A B 0.0639f
C27 a_109_297# C 0.00356f
C28 a_205_297# VGND 3.36e-19
C29 A X 0.00133f
C30 a_277_297# VPWR 7.48e-19
C31 VPWR B 0.193f
C32 C D 0.0954f
C33 A VGND 0.016f
C34 VPWR X 0.0878f
C35 a_27_297# a_277_297# 0.00876f
C36 a_27_297# B 0.159f
C37 VGND VPWR 0.0546f
C38 a_27_297# X 0.0991f
C39 a_27_297# VGND 0.235f
C40 a_109_297# VPWR 9.23e-19
C41 A D 2.13e-19
C42 a_277_297# B 2.29e-19
C43 VPWR D 0.00503f
C44 a_277_297# X 6.43e-20
C45 X B 6.42e-19
C46 a_109_297# a_27_297# 0.00695f
C47 a_277_297# VGND 4.65e-19
C48 VGND B 0.0159f
C49 VGND VNB 0.367f
C50 X VNB 0.0883f
C51 A VNB 0.109f
C52 C VNB 0.105f
C53 D VNB 0.175f
C54 B VNB 0.115f
C55 VPWR VNB 0.29f
C56 VPB VNB 0.605f
C57 a_27_297# VNB 0.163f
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
C0 VGND VPB 0.35f
C1 VPWR VPB 0.137f
C2 VGND VPWR 1.57f
C3 VPWR VNB 1.67f
C4 VGND VNB 1.47f
C5 VPB VNB 1.14f
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
C0 B a_27_47# 0.0794f
C1 C VPB 0.0742f
C2 C VPWR 0.0182f
C3 VPB a_27_47# 0.092f
C4 VGND X 0.0588f
C5 C a_369_47# 0.00448f
C6 VPWR a_27_47# 0.106f
C7 A_N a_27_47# 0.237f
C8 VGND a_193_413# 0.0915f
C9 C a_469_47# 0.00202f
C10 D VGND 0.0372f
C11 VGND a_297_47# 0.00183f
C12 a_193_413# X 0.108f
C13 D X 0.0168f
C14 VGND B 0.037f
C15 D a_193_413# 0.155f
C16 VPB VGND 0.0123f
C17 VGND VPWR 0.0727f
C18 a_297_47# a_193_413# 0.00137f
C19 VGND A_N 0.0205f
C20 VGND a_369_47# 0.00505f
C21 VGND a_469_47# 0.00551f
C22 B a_193_413# 0.144f
C23 VPB X 0.0108f
C24 C VGND 0.0395f
C25 VPB a_193_413# 0.0644f
C26 VPWR X 0.0586f
C27 VGND a_27_47# 0.103f
C28 VPWR a_193_413# 0.281f
C29 a_193_413# A_N 0.00151f
C30 D VPB 0.0763f
C31 a_297_47# B 0.00353f
C32 a_369_47# a_193_413# 0.00181f
C33 a_469_47# X 0.001f
C34 D VPWR 0.0186f
C35 a_469_47# a_193_413# 0.00109f
C36 C X 0.00479f
C37 a_297_47# VPWR 2.82e-19
C38 C a_193_413# 0.0389f
C39 D a_469_47# 0.00183f
C40 a_193_413# a_27_47# 0.125f
C41 VPB B 0.089f
C42 D C 0.183f
C43 B VPWR 0.0186f
C44 B a_369_47# 0.00129f
C45 VPB VPWR 0.0818f
C46 VPB A_N 0.0832f
C47 VPWR A_N 0.02f
C48 VPWR a_369_47# 6.65e-19
C49 C B 0.164f
C50 VPWR a_469_47# 7.77e-19
C51 VGND VNB 0.456f
C52 X VNB 0.0934f
C53 VPWR VNB 0.368f
C54 D VNB 0.123f
C55 C VNB 0.108f
C56 B VNB 0.12f
C57 A_N VNB 0.198f
C58 VPB VNB 0.782f
C59 a_193_413# VNB 0.136f
C60 a_27_47# VNB 0.224f
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
C0 a_109_93# B 0.0802f
C1 a_209_311# a_368_53# 0.0026f
C2 a_209_311# VPWR 0.155f
C3 a_209_311# VGND 0.131f
C4 VPWR B 0.131f
C5 VPB C 0.0339f
C6 VGND B 0.00796f
C7 VPB X 0.0119f
C8 a_209_311# B 0.0609f
C9 VPB A_N 0.111f
C10 VPB a_109_93# 0.0652f
C11 X C 0.0176f
C12 VPB VPWR 0.104f
C13 VPB VGND 0.00909f
C14 A_N C 7.6e-19
C15 a_109_93# C 3.91e-20
C16 a_209_311# VPB 0.0515f
C17 a_296_53# a_109_93# 1.84e-19
C18 X A_N 1.44e-19
C19 VPB B 0.0914f
C20 a_368_53# C 0.00415f
C21 C VPWR 0.005f
C22 VGND C 0.0678f
C23 a_296_53# VPWR 1.15e-19
C24 a_109_93# A_N 0.117f
C25 a_296_53# VGND 6.07e-19
C26 X VPWR 0.0732f
C27 a_209_311# C 0.19f
C28 X VGND 0.0647f
C29 A_N VPWR 0.0513f
C30 C B 0.0671f
C31 a_296_53# a_209_311# 0.0049f
C32 A_N VGND 0.045f
C33 a_109_93# VPWR 0.0984f
C34 a_109_93# VGND 0.0784f
C35 a_209_311# X 0.0877f
C36 a_209_311# A_N 0.00515f
C37 X B 0.00119f
C38 a_368_53# VPWR 4.26e-19
C39 A_N B 2.03e-19
C40 a_368_53# VGND 0.0031f
C41 VGND VPWR 0.0657f
C42 a_209_311# a_109_93# 0.168f
C43 VGND VNB 0.44f
C44 X VNB 0.0925f
C45 C VNB 0.114f
C46 B VNB 0.101f
C47 VPWR VNB 0.342f
C48 A_N VNB 0.197f
C49 VPB VNB 0.693f
C50 a_209_311# VNB 0.143f
C51 a_109_93# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
C0 X A 0.014f
C1 VPWR A 0.022f
C2 VPWR X 0.317f
C3 VGND a_27_47# 0.148f
C4 A a_27_47# 0.195f
C5 X a_27_47# 0.328f
C6 VPWR a_27_47# 0.219f
C7 VGND VPB 0.00583f
C8 VPB A 0.0321f
C9 VPB X 0.0122f
C10 VPB VPWR 0.0632f
C11 VPB a_27_47# 0.139f
C12 VGND A 0.0431f
C13 VGND X 0.216f
C14 VGND VPWR 0.057f
C15 VGND VNB 0.358f
C16 X VNB 0.067f
C17 VPWR VNB 0.308f
C18 A VNB 0.148f
C19 VPB VNB 0.605f
C20 a_27_47# VNB 0.543f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
C0 A VPB 0.0806f
C1 VGND a_59_75# 0.116f
C2 VPWR VPB 0.0729f
C3 VPWR A 0.0362f
C4 B a_59_75# 0.143f
C5 X a_59_75# 0.109f
C6 VPB a_59_75# 0.0563f
C7 A a_59_75# 0.0809f
C8 VPWR a_59_75# 0.15f
C9 VGND a_145_75# 0.00468f
C10 a_145_75# X 5.76e-19
C11 VPWR a_145_75# 6.31e-19
C12 a_145_75# a_59_75# 0.00658f
C13 B VGND 0.0115f
C14 VGND X 0.0993f
C15 VGND VPB 0.008f
C16 VGND A 0.0147f
C17 B X 0.00276f
C18 VGND VPWR 0.0461f
C19 B VPB 0.0629f
C20 B A 0.0971f
C21 B VPWR 0.0117f
C22 VPB X 0.0127f
C23 A X 1.68e-19
C24 VPWR X 0.111f
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_191_297# B 0.00223f
C1 D VPB 0.0376f
C2 a_191_297# VGND 9.29e-19
C3 B A 0.11f
C4 D Y 0.108f
C5 VGND A 0.0526f
C6 D VPWR 0.0128f
C7 Y VPB 0.0127f
C8 D C 0.0523f
C9 a_297_297# Y 1.24e-19
C10 VPWR VPB 0.0524f
C11 VPWR Y 0.0561f
C12 C VPB 0.0299f
C13 D VGND 0.0456f
C14 C Y 0.125f
C15 a_297_297# VPWR 0.00317f
C16 a_109_297# Y 0.0122f
C17 VPB B 0.0304f
C18 VPWR C 0.0509f
C19 Y B 0.0403f
C20 VGND VPB 0.0048f
C21 VPWR a_109_297# 0.00576f
C22 VGND Y 0.151f
C23 a_297_297# B 0.0132f
C24 a_109_297# C 0.0062f
C25 a_297_297# VGND 8.1e-19
C26 VPWR B 0.0887f
C27 a_191_297# Y 0.00142f
C28 VPB A 0.041f
C29 VPWR VGND 0.0492f
C30 C B 0.173f
C31 Y A 0.0175f
C32 C VGND 0.0184f
C33 a_297_297# A 3.16e-19
C34 a_109_297# VGND 0.00181f
C35 a_191_297# VPWR 0.0049f
C36 a_191_297# C 0.0195f
C37 VPWR A 0.0483f
C38 C A 0.00268f
C39 VGND B 0.0191f
C40 VGND VNB 0.322f
C41 VPWR VNB 0.276f
C42 Y VNB 0.0645f
C43 A VNB 0.174f
C44 B VNB 0.0968f
C45 C VNB 0.0911f
C46 D VNB 0.159f
C47 VPB VNB 0.516f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 VPWR A 0.0217f
C1 X A 8.48e-19
C2 X VPWR 0.0896f
C3 VGND a_75_212# 0.105f
C4 A a_75_212# 0.178f
C5 VPWR a_75_212# 0.134f
C6 X a_75_212# 0.107f
C7 VGND VPB 0.00507f
C8 VPB A 0.0525f
C9 VPB VPWR 0.0355f
C10 VPB X 0.0128f
C11 VPB a_75_212# 0.0571f
C12 VGND A 0.0184f
C13 VGND VPWR 0.0289f
C14 VGND X 0.0545f
C15 VGND VNB 0.207f
C16 VPWR VNB 0.176f
C17 X VNB 0.0942f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_75_212# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 X A 8.48e-19
C1 VPWR A 0.0215f
C2 VPWR X 0.0897f
C3 VGND a_27_47# 0.105f
C4 A a_27_47# 0.181f
C5 X a_27_47# 0.107f
C6 VPWR a_27_47# 0.135f
C7 VGND VPB 0.00505f
C8 VPB A 0.0524f
C9 VPB X 0.0128f
C10 VPB VPWR 0.0355f
C11 VPB a_27_47# 0.0592f
C12 VGND A 0.0184f
C13 VGND X 0.0546f
C14 VGND VPWR 0.029f
C15 VGND VNB 0.207f
C16 X VNB 0.0941f
C17 VPWR VNB 0.175f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_27_47# VNB 0.208f
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
C0 X a_62_47# 0.156f
C1 VPWR VPB 0.103f
C2 a_841_47# a_664_47# 0.134f
C3 VPWR A 0.0174f
C4 VPB a_62_47# 0.0515f
C5 VPWR a_664_47# 0.131f
C6 A a_62_47# 0.244f
C7 VPWR a_841_47# 0.0614f
C8 VPWR a_62_47# 0.149f
C9 VGND a_381_47# 0.125f
C10 a_558_47# a_381_47# 0.16f
C11 VGND a_558_47# 0.0816f
C12 X a_381_47# 0.318f
C13 VPB a_381_47# 0.0447f
C14 VGND X 0.106f
C15 a_381_47# A 5.42e-19
C16 VGND VPB 0.008f
C17 a_558_47# X 0.0144f
C18 VGND A 0.0176f
C19 VPB a_558_47# 0.115f
C20 VGND a_664_47# 0.125f
C21 VPWR a_381_47# 0.134f
C22 VGND a_841_47# 0.0585f
C23 a_558_47# a_664_47# 0.314f
C24 VPB X 0.126f
C25 VGND VPWR 0.0902f
C26 a_558_47# a_841_47# 0.00368f
C27 X A 0.0142f
C28 VGND a_62_47# 0.144f
C29 X a_664_47# 6.67e-19
C30 VPWR a_558_47# 0.084f
C31 VPB A 0.105f
C32 VPB a_664_47# 0.043f
C33 VPB a_841_47# 0.0108f
C34 VPWR X 0.108f
C35 VGND VNB 0.537f
C36 VPWR VNB 0.439f
C37 X VNB 0.163f
C38 A VNB 0.198f
C39 VPB VNB 0.959f
C40 a_841_47# VNB 0.0929f
C41 a_664_47# VNB 0.13f
C42 a_558_47# VNB 0.164f
C43 a_381_47# VNB 0.11f
C44 a_62_47# VNB 0.169f
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 a_47_47# VPWR 0.273f
C1 a_285_47# VPWR 0.00255f
C2 A VPWR 0.0349f
C3 VPB Y 0.00878f
C4 VPB VGND 0.00568f
C5 a_377_297# VPWR 0.00559f
C6 VPB B 0.0643f
C7 VPB a_47_47# 0.0444f
C8 VPB a_285_47# 5.53e-19
C9 VGND Y 0.0381f
C10 VPB A 0.0822f
C11 B Y 0.00334f
C12 a_129_47# VGND 0.00547f
C13 a_47_47# Y 0.143f
C14 a_129_47# B 0.00236f
C15 a_129_47# a_47_47# 0.00369f
C16 VGND B 0.0389f
C17 VPB VPWR 0.0718f
C18 a_285_47# Y 0.0439f
C19 Y A 0.00181f
C20 VGND a_47_47# 0.104f
C21 a_47_47# B 0.356f
C22 VGND a_285_47# 0.211f
C23 VGND A 0.0635f
C24 a_377_297# Y 0.00188f
C25 a_285_47# B 0.067f
C26 B A 0.236f
C27 Y VPWR 0.107f
C28 a_47_47# a_285_47# 0.0175f
C29 a_47_47# A 0.0307f
C30 a_129_47# VPWR 9.47e-19
C31 a_377_297# VGND 0.00125f
C32 a_377_297# B 0.00254f
C33 VGND VPWR 0.0665f
C34 a_285_47# A 0.0353f
C35 B VPWR 0.0408f
C36 a_377_297# a_47_47# 0.00899f
C37 VGND VNB 0.4f
C38 Y VNB 0.0783f
C39 VPWR VNB 0.352f
C40 A VNB 0.217f
C41 B VNB 0.212f
C42 VPB VNB 0.693f
C43 a_285_47# VNB 0.0174f
C44 a_47_47# VNB 0.199f
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
C0 B1 a_80_21# 0.0964f
C1 C1 VPWR 0.0137f
C2 A2 a_80_21# 0.128f
C3 VPWR a_80_21# 0.119f
C4 A1 a_80_21# 0.111f
C5 C1 VPB 0.0379f
C6 a_300_47# a_80_21# 0.00997f
C7 VPB a_80_21# 0.0661f
C8 C1 a_80_21# 0.079f
C9 a_217_297# VGND 0.00342f
C10 X VGND 0.0654f
C11 X a_217_297# 0.00271f
C12 a_472_297# VGND 0.00188f
C13 a_472_297# a_217_297# 0.00517f
C14 B1 VGND 0.0175f
C15 X a_472_297# 2.6e-19
C16 B1 a_217_297# 0.00651f
C17 A2 VGND 0.0191f
C18 A2 a_217_297# 0.0135f
C19 VPWR VGND 0.0665f
C20 VGND A1 0.0147f
C21 X B1 1.18e-19
C22 VPWR a_217_297# 0.197f
C23 a_217_297# A1 0.0124f
C24 a_300_47# VGND 0.00536f
C25 VPB VGND 0.00775f
C26 X A2 6.82e-19
C27 a_472_297# B1 1.87e-19
C28 VPB a_217_297# 0.00494f
C29 X VPWR 0.0884f
C30 X A1 3.62e-19
C31 C1 VGND 0.0176f
C32 X a_300_47# 5.31e-19
C33 X VPB 0.0118f
C34 a_472_297# VPWR 0.00703f
C35 C1 a_217_297# 0.00262f
C36 VGND a_80_21# 0.293f
C37 a_217_297# a_80_21# 0.127f
C38 X C1 7.15e-20
C39 B1 VPWR 0.0129f
C40 B1 A1 0.0834f
C41 X a_80_21# 0.118f
C42 B1 VPB 0.0267f
C43 A2 VPWR 0.0161f
C44 A2 A1 0.0881f
C45 a_472_297# a_80_21# 0.0164f
C46 VPWR A1 0.0149f
C47 A2 VPB 0.0384f
C48 VPWR a_300_47# 8.53e-19
C49 a_300_47# A1 5.95e-19
C50 VPWR VPB 0.0754f
C51 C1 B1 0.0846f
C52 VPB A1 0.0266f
C53 VGND VNB 0.385f
C54 VPWR VNB 0.325f
C55 X VNB 0.0899f
C56 C1 VNB 0.144f
C57 B1 VNB 0.0899f
C58 A1 VNB 0.0905f
C59 A2 VNB 0.108f
C60 VPB VNB 0.693f
C61 a_217_297# VNB 0.00117f
C62 a_80_21# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_27_47# C 0.0516f
C1 VGND X 0.0903f
C2 a_109_47# B 0.00153f
C3 a_303_47# C 0.00527f
C4 B C 0.161f
C5 VPB D 0.0782f
C6 a_109_47# VGND 0.00223f
C7 VGND C 0.0408f
C8 a_109_47# C 1.72e-20
C9 VPB VPWR 0.077f
C10 VPB A 0.0907f
C11 VPB a_27_47# 0.082f
C12 VPB B 0.0643f
C13 VPWR D 0.0207f
C14 VPB X 0.0111f
C15 a_197_47# VPWR 5.24e-19
C16 VPB VGND 0.00852f
C17 a_27_47# D 0.107f
C18 a_197_47# a_27_47# 0.00167f
C19 VPWR A 0.044f
C20 VPB C 0.0609f
C21 a_303_47# D 0.00119f
C22 VPWR a_27_47# 0.326f
C23 X D 0.00746f
C24 a_197_47# B 0.00623f
C25 VGND D 0.0898f
C26 a_27_47# A 0.153f
C27 VPWR a_303_47# 4.83e-19
C28 VPWR B 0.0231f
C29 a_197_47# VGND 0.00387f
C30 VPWR X 0.0945f
C31 A B 0.0839f
C32 D C 0.18f
C33 VPWR VGND 0.0662f
C34 a_27_47# a_303_47# 0.00119f
C35 a_27_47# B 0.13f
C36 VGND A 0.0151f
C37 a_197_47# C 0.00123f
C38 a_27_47# X 0.0754f
C39 a_109_47# VPWR 4.66e-19
C40 a_27_47# VGND 0.132f
C41 VPWR C 0.021f
C42 a_109_47# a_27_47# 0.00578f
C43 a_303_47# VGND 0.00381f
C44 VGND B 0.0453f
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
C0 B1 a_76_199# 0.00185f
C1 X VPB 0.0113f
C2 X A1_N 0.00211f
C3 VPB a_76_199# 0.0817f
C4 VGND A2_N 0.0174f
C5 A1_N a_76_199# 0.119f
C6 B2 a_76_199# 0.0626f
C7 VGND a_226_47# 0.149f
C8 a_226_297# a_76_199# 0.00354f
C9 VPWR VGND 0.0743f
C10 a_556_47# a_76_199# 0.0017f
C11 VGND a_489_413# 0.0058f
C12 X a_76_199# 0.0995f
C13 a_226_47# A2_N 0.141f
C14 VGND B1 0.0471f
C15 VPWR A2_N 0.00449f
C16 VPWR a_226_47# 0.0187f
C17 VPB VGND 0.0128f
C18 VGND A1_N 0.0261f
C19 a_489_413# a_226_47# 0.00579f
C20 VGND B2 0.0335f
C21 VGND a_226_297# 5.63e-19
C22 VPWR a_489_413# 0.143f
C23 VGND a_556_47# 0.00639f
C24 VPB A2_N 0.0327f
C25 X VGND 0.0627f
C26 VPB a_226_47# 0.111f
C27 A1_N A2_N 0.11f
C28 VPWR B1 0.0188f
C29 VGND a_76_199# 0.108f
C30 A1_N a_226_47# 0.0209f
C31 a_226_47# B2 0.0975f
C32 VPWR VPB 0.0951f
C33 a_489_413# B1 0.0382f
C34 a_226_297# a_226_47# 0.00128f
C35 VPWR A1_N 0.00672f
C36 VPWR B2 0.0161f
C37 VPB a_489_413# 0.015f
C38 X A2_N 2.55e-19
C39 VPWR a_226_297# 8.54e-19
C40 a_489_413# B2 0.0541f
C41 X a_226_47# 0.0108f
C42 A2_N a_76_199# 0.0125f
C43 VPWR a_556_47# 7.24e-19
C44 a_226_47# a_76_199# 0.188f
C45 VPB B1 0.0803f
C46 VPWR X 0.0589f
C47 B1 B2 0.182f
C48 VPWR a_76_199# 0.2f
C49 VPB A1_N 0.0339f
C50 VPB B2 0.0645f
C51 a_489_413# a_76_199# 0.0473f
C52 A1_N a_226_297# 0.00184f
C53 a_556_47# B2 0.00291f
C54 VGND VNB 0.462f
C55 A2_N VNB 0.103f
C56 A1_N VNB 0.111f
C57 VPWR VNB 0.369f
C58 X VNB 0.0975f
C59 B1 VNB 0.206f
C60 B2 VNB 0.106f
C61 VPB VNB 0.782f
C62 a_489_413# VNB 0.0254f
C63 a_226_47# VNB 0.162f
C64 a_76_199# VNB 0.141f
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
C0 X D 0.0193f
C1 a_27_47# A_N 0.0906f
C2 a_223_47# VGND 0.199f
C3 VPWR D 0.0143f
C4 VPWR X 0.0582f
C5 a_223_47# a_429_93# 0.00492f
C6 VGND A_N 0.0146f
C7 a_223_47# VPB 0.0799f
C8 a_223_47# D 4.03e-19
C9 VPB A_N 0.0848f
C10 a_223_47# VPWR 0.114f
C11 VPWR A_N 0.0318f
C12 a_343_93# a_615_93# 0.00103f
C13 a_615_93# C 0.00407f
C14 a_223_47# A_N 0.00833f
C15 a_343_93# a_515_93# 0.00115f
C16 a_343_93# B_N 0.00112f
C17 VGND a_615_93# 0.0044f
C18 C a_515_93# 0.00389f
C19 C B_N 9.56e-20
C20 a_615_93# D 0.00564f
C21 a_343_93# C 0.0397f
C22 a_615_93# VPWR 8.49e-19
C23 a_27_47# B_N 0.138f
C24 VGND a_515_93# 0.00408f
C25 VGND B_N 0.0427f
C26 a_343_93# a_27_47# 0.0406f
C27 B_N VPB 0.0646f
C28 a_343_93# VGND 0.0548f
C29 D B_N 6.67e-20
C30 VPWR a_515_93# 7.86e-19
C31 X B_N 4.64e-20
C32 a_343_93# a_429_93# 0.00484f
C33 a_343_93# VPB 0.0857f
C34 VPWR B_N 0.0168f
C35 VGND C 0.025f
C36 a_223_47# a_515_93# 0.00482f
C37 a_343_93# D 0.114f
C38 a_343_93# X 0.126f
C39 C VPB 0.0686f
C40 a_223_47# B_N 0.0431f
C41 a_343_93# VPWR 0.255f
C42 C D 0.163f
C43 B_N A_N 0.117f
C44 VGND a_27_47# 0.0715f
C45 a_343_93# a_223_47# 0.269f
C46 C VPWR 0.012f
C47 a_27_47# VPB 0.154f
C48 a_223_47# C 0.151f
C49 VGND a_429_93# 0.00122f
C50 VGND VPB 0.0167f
C51 a_27_47# VPWR 0.0897f
C52 VGND D 0.0414f
C53 VGND X 0.0609f
C54 VGND VPWR 0.0906f
C55 D VPB 0.081f
C56 a_223_47# a_27_47# 0.267f
C57 X VPB 0.0103f
C58 a_429_93# VPWR 5.19e-19
C59 VPWR VPB 0.106f
C60 VGND VNB 0.553f
C61 X VNB 0.0908f
C62 VPWR VNB 0.453f
C63 D VNB 0.124f
C64 C VNB 0.107f
C65 B_N VNB 0.134f
C66 A_N VNB 0.144f
C67 VPB VNB 0.959f
C68 a_343_93# VNB 0.172f
C69 a_223_47# VNB 0.141f
C70 a_27_47# VNB 0.259f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VPWR a_35_297# 0.096f
C1 X B 0.0149f
C2 X A 0.00166f
C3 B a_35_297# 0.203f
C4 X a_285_47# 0.00206f
C5 A a_35_297# 0.0633f
C6 X VPB 0.0154f
C7 a_285_47# a_35_297# 0.00723f
C8 VPB a_35_297# 0.0699f
C9 X a_35_297# 0.166f
C10 VGND a_117_297# 0.00177f
C11 VGND a_285_297# 0.00394f
C12 VPWR a_117_297# 0.00852f
C13 B a_117_297# 0.00777f
C14 VGND VPWR 0.0643f
C15 VGND B 0.0304f
C16 a_285_297# VPWR 0.246f
C17 VGND A 0.0325f
C18 B a_285_297# 0.0553f
C19 VGND a_285_47# 0.00552f
C20 VGND VPB 0.00696f
C21 a_285_297# A 0.00749f
C22 X a_117_297# 2.25e-19
C23 a_285_297# VPB 0.0133f
C24 a_117_297# a_35_297# 0.00641f
C25 B VPWR 0.0703f
C26 VGND X 0.173f
C27 VPWR A 0.0348f
C28 VGND a_35_297# 0.177f
C29 VPWR a_285_47# 8.6e-19
C30 VPWR VPB 0.0689f
C31 X a_285_297# 0.0712f
C32 B A 0.221f
C33 a_285_297# a_35_297# 0.025f
C34 B a_285_47# 3.98e-19
C35 B VPB 0.0697f
C36 X VPWR 0.0537f
C37 VPB A 0.051f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 VGND A 0.0158f
C1 a_215_297# B 0.159f
C2 X A 0.00127f
C3 X VGND 0.0359f
C4 a_109_53# VPWR 0.0418f
C5 a_109_53# A 1.19e-19
C6 VPWR B 0.255f
C7 a_109_53# VGND 0.118f
C8 A B 0.0666f
C9 VGND B 0.0161f
C10 X B 6.65e-19
C11 a_109_53# B 0.0246f
C12 C a_465_297# 6.89e-19
C13 VPB D_N 0.0461f
C14 a_215_297# a_465_297# 0.00827f
C15 a_297_297# C 0.00375f
C16 a_215_297# D_N 3.19e-19
C17 a_465_297# VPWR 7.08e-19
C18 a_297_297# a_215_297# 0.00659f
C19 C VPB 0.0337f
C20 D_N VPWR 0.0412f
C21 A a_465_297# 5.42e-19
C22 VGND a_465_297# 5.02e-19
C23 C a_215_297# 0.161f
C24 VGND D_N 0.0531f
C25 a_297_297# VPWR 8.59e-19
C26 a_215_297# VPB 0.0508f
C27 a_297_297# VGND 6.5e-19
C28 C a_392_297# 0.00267f
C29 C VPWR 0.00753f
C30 a_109_53# D_N 0.0889f
C31 C A 0.0281f
C32 VPB VPWR 0.122f
C33 C VGND 0.0202f
C34 a_297_297# a_109_53# 7.06e-21
C35 VPB A 0.0325f
C36 VGND VPB 0.0115f
C37 a_215_297# a_392_297# 0.00419f
C38 a_215_297# VPWR 0.0871f
C39 X VPB 0.011f
C40 a_215_297# A 0.157f
C41 a_215_297# VGND 0.237f
C42 a_109_53# C 0.0984f
C43 a_215_297# X 0.0991f
C44 a_109_53# VPB 0.0547f
C45 C B 0.0893f
C46 a_392_297# VPWR 5.29e-19
C47 VPB B 0.116f
C48 A VPWR 0.0073f
C49 a_392_297# VGND 3.44e-19
C50 a_109_53# a_215_297# 0.0807f
C51 VGND VPWR 0.075f
C52 X VPWR 0.0885f
C53 VGND VNB 0.469f
C54 X VNB 0.0884f
C55 A VNB 0.108f
C56 C VNB 0.101f
C57 D_N VNB 0.185f
C58 B VNB 0.101f
C59 VPWR VNB 0.399f
C60 VPB VNB 0.782f
C61 a_109_53# VNB 0.159f
C62 a_215_297# VNB 0.142f
.ends

.subckt therm b[0] b[1] b[2] b[3] p[0] p[10] p[11] p[12] p[13] p[14] p[1] p[2] p[3]
+ p[4] p[5] p[6] p[7] p[8] net7 _04_ net19 net15 net14 _31_/a_35_297# input7/a_27_47#
+ _27_/a_27_297# input1/a_75_212# input5/a_62_47# net2 input5/a_841_47# _19_ net8
+ _17_ _01_ _44_/a_250_297# p[9] input15/a_27_47# _20_ _14_ net1 _16_ net9 VPWR net5
+ VGND _29_/a_29_53#
X_49_ net7 _02_ _19_ _20_ _21_ VGND VGND VPWR VPWR net17 _49_/a_208_47# _49_/a_75_199#
+ _49_/a_544_297# _49_/a_315_47# _49_/a_201_297# sky130_fd_sc_hd__a311o_1
X_48_ net11 _02_ _07_ VGND VGND VPWR VPWR _21_ _48_/a_181_47# _48_/a_109_47# _48_/a_27_47#
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ net5 _12_ _17_ VGND VGND VPWR VPWR _20_ _47_/a_384_47# _47_/a_81_21# _47_/a_299_297#
+ sky130_fd_sc_hd__a21o_1
X_46_ _04_ VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__inv_2
X_29_ net11 net13 net12 VGND VGND VPWR VPWR _03_ _29_/a_29_53# _29_/a_183_297# _29_/a_111_297#
+ sky130_fd_sc_hd__or3_1
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28_ _00_ _01_ VGND VGND VPWR VPWR _02_ _28_/a_109_297# sky130_fd_sc_hd__nor2_1
X_45_ _02_ _09_ _12_ _13_ _18_ VGND VGND VPWR VPWR net16 _45_/a_193_297# _45_/a_465_47#
+ _45_/a_205_47# _45_/a_109_297# _45_/a_27_47# sky130_fd_sc_hd__a221o_1
X_44_ net14 _14_ _15_ _17_ net2 VGND VGND VPWR VPWR _18_ _44_/a_256_47# _44_/a_584_47#
+ _44_/a_93_21# _44_/a_250_297# _44_/a_346_47# sky130_fd_sc_hd__a32o_1
X_27_ net14 net15 net3 net2 VGND VGND VPWR VPWR _01_ _27_/a_277_297# _27_/a_205_297#
+ _27_/a_27_297# _27_/a_109_297# sky130_fd_sc_hd__or4_1
XFILLER_0_7_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_26_ net5 net4 net6 VGND VGND VPWR VPWR _00_ _26_/a_29_53# _26_/a_183_297# _26_/a_111_297#
+ sky130_fd_sc_hd__or3_1
X_43_ _00_ _06_ _10_ _16_ VGND VGND VPWR VPWR _17_ _43_/a_369_47# _43_/a_469_47# _43_/a_297_47#
+ _43_/a_193_413# _43_/a_27_47# sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_42_ net3 net15 net14 VGND VGND VPWR VPWR _16_ _42_/a_109_93# _42_/a_368_53# _42_/a_209_311#
+ _42_/a_296_53# sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_3_Left_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND VPWR VPWR b[0] output16/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_41_ _06_ _10_ VGND VGND VPWR VPWR _15_ _41_/a_145_75# _41_/a_59_75# sky130_fd_sc_hd__and2_1
Xoutput17 net17 VGND VGND VPWR VPWR b[1] output17/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_40_ net15 net3 net2 _00_ VGND VGND VPWR VPWR _14_ _40_/a_297_297# _40_/a_191_297#
+ _40_/a_109_297# sky130_fd_sc_hd__nor4_1
Xoutput18 net18 VGND VGND VPWR VPWR b[2] output18/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR b[3] output19/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_7_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 p[0] VGND VGND VPWR VPWR net1 input1/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput2 p[10] VGND VGND VPWR VPWR net2 input2/a_27_47# sky130_fd_sc_hd__buf_1
Xinput3 p[11] VGND VGND VPWR VPWR net3 input3/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 p[12] VGND VGND VPWR VPWR net4 input4/a_75_212# sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 p[13] VGND VGND VPWR VPWR net5 input5/a_664_47# input5/a_841_47# input5/a_381_47#
+ input5/a_62_47# input5/a_558_47# sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_1_Left_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 p[14] VGND VGND VPWR VPWR net6 input6/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 p[1] VGND VGND VPWR VPWR net7 input7/a_27_47# sky130_fd_sc_hd__buf_1
Xinput10 p[4] VGND VGND VPWR VPWR net10 input10/a_27_47# sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 p[2] VGND VGND VPWR VPWR net8 input8/a_27_47# sky130_fd_sc_hd__buf_1
Xinput11 p[5] VGND VGND VPWR VPWR net11 input11/a_27_47# sky130_fd_sc_hd__buf_1
X_39_ net5 net6 VGND VGND VPWR VPWR _13_ _39_/a_129_47# _39_/a_47_47# _39_/a_285_47#
+ _39_/a_377_297# sky130_fd_sc_hd__xnor2_1
Xinput9 p[3] VGND VGND VPWR VPWR net9 input9/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput12 p[6] VGND VGND VPWR VPWR net12 input12/a_27_47# sky130_fd_sc_hd__buf_1
X_55_ _14_ _15_ _20_ _22_ VGND VGND VPWR VPWR net19 _55_/a_472_297# _55_/a_80_21#
+ _55_/a_300_47# _55_/a_217_297# sky130_fd_sc_hd__a211o_1
X_38_ net4 _06_ _10_ _11_ VGND VGND VPWR VPWR _12_ _38_/a_109_47# _38_/a_197_47# _38_/a_303_47#
+ _38_/a_27_47# sky130_fd_sc_hd__and4_1
X_54_ _25_ VGND VGND VPWR VPWR net18 _54_/a_75_212# sky130_fd_sc_hd__clkbuf_1
Xinput13 p[7] VGND VGND VPWR VPWR net13 input13/a_27_47# sky130_fd_sc_hd__buf_1
X_37_ net14 net15 net3 net2 VGND VGND VPWR VPWR _11_ _37_/a_109_47# _37_/a_197_47#
+ _37_/a_303_47# _37_/a_27_47# sky130_fd_sc_hd__and4_1
X_53_ _21_ _22_ _24_ VGND VGND VPWR VPWR _25_ _53_/a_29_53# _53_/a_183_297# _53_/a_111_297#
+ sky130_fd_sc_hd__or3_1
Xinput14 p[8] VGND VGND VPWR VPWR net14 input14/a_27_47# sky130_fd_sc_hd__buf_1
X_36_ net11 net10 net13 net12 VGND VGND VPWR VPWR _10_ _36_/a_109_47# _36_/a_197_47#
+ _36_/a_303_47# _36_/a_27_47# sky130_fd_sc_hd__and4_1
X_52_ _02_ _06_ _23_ _12_ net5 VGND VGND VPWR VPWR _24_ _52_/a_256_47# _52_/a_584_47#
+ _52_/a_93_21# _52_/a_250_297# _52_/a_346_47# sky130_fd_sc_hd__a32o_1
X_35_ _04_ _05_ _07_ _08_ VGND VGND VPWR VPWR _09_ _35_/a_489_413# _35_/a_226_47#
+ _35_/a_556_47# _35_/a_226_297# _35_/a_76_199# sky130_fd_sc_hd__a2bb2o_1
Xinput15 p[9] VGND VGND VPWR VPWR net15 input15/a_27_47# sky130_fd_sc_hd__buf_1
X_51_ _03_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__inv_2
X_34_ net11 net12 VGND VGND VPWR VPWR _08_ _34_/a_129_47# _34_/a_47_47# _34_/a_285_47#
+ _34_/a_377_297# sky130_fd_sc_hd__xnor2_1
X_33_ net13 _06_ net10 VGND VGND VPWR VPWR _07_ _33_/a_109_93# _33_/a_368_53# _33_/a_209_311#
+ _33_/a_296_53# sky130_fd_sc_hd__and3b_1
X_50_ net5 net6 _15_ _11_ VGND VGND VPWR VPWR _22_ _50_/a_515_93# _50_/a_223_47# _50_/a_615_93#
+ _50_/a_343_93# _50_/a_429_93# _50_/a_27_47# sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ net7 net1 net9 net8 VGND VGND VPWR VPWR _06_ _32_/a_109_47# _32_/a_197_47# _32_/a_303_47#
+ _32_/a_27_47# sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_5_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31_ net7 net8 VGND VGND VPWR VPWR _05_ _31_/a_117_297# _31_/a_285_297# _31_/a_285_47#
+ _31_/a_35_297# sky130_fd_sc_hd__xor2_1
X_30_ net9 net10 _03_ net1 VGND VGND VPWR VPWR _04_ _30_/a_465_297# _30_/a_297_297#
+ _30_/a_215_297# _30_/a_392_297# _30_/a_109_53# sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
C0 _13_ _09_ 0.0927f
C1 net9 _30_/a_109_53# 0.0193f
C2 net9 _50_/a_223_47# 2e-19
C3 _38_/a_27_47# net5 1.76e-19
C4 _11_ _17_ 0.197f
C5 input2/a_27_47# _30_/a_109_53# 1.54e-20
C6 input9/a_75_212# _03_ 9.32e-20
C7 net1 _02_ 0.00251f
C8 output19/a_27_47# _42_/a_109_93# 1.56e-20
C9 input3/a_27_47# _44_/a_250_297# 2.07e-19
C10 _11_ net9 5.39e-19
C11 _55_/a_300_47# _02_ 0.00371f
C12 _15_ p[12] 0.0162f
C13 net7 net17 0.2f
C14 _30_/a_215_297# _05_ 0.0453f
C15 _50_/a_429_93# net4 4.16e-19
C16 _50_/a_343_93# net6 0.00214f
C17 _23_ b[2] 2.87e-20
C18 _21_ net16 1.89e-19
C19 input5/a_62_47# net5 0.00329f
C20 _33_/a_296_53# net10 8.22e-20
C21 _50_/a_223_47# _26_/a_29_53# 0.00124f
C22 net10 net4 8.28e-22
C23 _39_/a_285_47# _17_ 7.36e-21
C24 _20_ _03_ 0.0794f
C25 _42_/a_109_93# net14 0.00351f
C26 p[11] p[10] 0.00241f
C27 _37_/a_27_47# net3 0.094f
C28 _43_/a_27_47# _00_ 0.0431f
C29 _13_ net10 4.52e-21
C30 _40_/a_109_297# net3 3.14e-19
C31 net2 _40_/a_191_297# 0.00143f
C32 VPWR _12_ 0.28f
C33 net5 _30_/a_215_297# 8.27e-21
C34 _11_ _26_/a_29_53# 1.09e-19
C35 VPWR _36_/a_27_47# -0.00832f
C36 p[2] _49_/a_201_297# 4.58e-20
C37 net18 _03_ 2.07e-21
C38 _44_/a_93_21# _16_ 0.00354f
C39 VPWR _14_ 0.186f
C40 net15 _49_/a_201_297# 1.41e-19
C41 _01_ _32_/a_303_47# 8.58e-19
C42 VPWR _09_ 0.297f
C43 p[12] net6 0.0941f
C44 input7/a_27_47# net1 0.0383f
C45 net9 _29_/a_111_297# 8.06e-21
C46 net16 _02_ 8.94e-19
C47 input6/a_27_47# output19/a_27_47# 0.107f
C48 b[3] _42_/a_209_311# 3.71e-19
C49 _44_/a_93_21# net15 0.00573f
C50 _35_/a_489_413# _07_ 0.00429f
C51 _18_ _03_ 7.25e-23
C52 net1 _32_/a_27_47# 0.0211f
C53 _37_/a_27_47# input15/a_27_47# 3.27e-19
C54 net9 _28_/a_109_297# 3.7e-19
C55 input5/a_381_47# net2 0.0138f
C56 _21_ _23_ 0.0217f
C57 input6/a_27_47# net14 7.05e-19
C58 _16_ net15 0.214f
C59 net13 _34_/a_47_47# 1.68e-19
C60 input5/a_381_47# net19 0.00173f
C61 _50_/a_429_93# VPWR -3.61e-19
C62 _25_ _12_ 1.23e-20
C63 p[0] VPWR 0.0839f
C64 p[10] net14 3.02e-19
C65 _03_ _07_ 0.0113f
C66 _42_/a_109_93# _27_/a_27_297# 1.35e-20
C67 _55_/a_472_297# VPWR 0.00488f
C68 _25_ _36_/a_27_47# 2.34e-20
C69 _15_ _42_/a_209_311# 0.0521f
C70 _25_ _09_ 1.49e-19
C71 input8/a_27_47# _31_/a_285_297# 1.04e-19
C72 VPWR net10 0.362f
C73 _17_ _42_/a_109_93# 7.83e-20
C74 _43_/a_193_413# _43_/a_369_47# -1.25e-19
C75 _37_/a_197_47# _15_ 3.02e-19
C76 _00_ _12_ 0.00396f
C77 _35_/a_489_413# _10_ 3.41e-19
C78 _14_ _00_ 0.133f
C79 net13 _19_ 4.45e-20
C80 b[3] input5/a_62_47# 0.00324f
C81 _50_/a_343_93# _20_ 0.00826f
C82 net13 p[3] 9.49e-19
C83 _00_ _09_ 9.35e-21
C84 _55_/a_217_297# _20_ 0.0013f
C85 _02_ p[13] 7.58e-20
C86 _02_ _23_ 0.0641f
C87 _52_/a_256_47# _23_ 6.66e-19
C88 _43_/a_193_413# p[9] 1.09e-19
C89 _22_ _35_/a_76_199# 6.58e-21
C90 net9 input5/a_841_47# 2.7e-19
C91 _53_/a_29_53# b[2] 6.22e-19
C92 p[1] input5/a_558_47# 1.61e-21
C93 _05_ _31_/a_285_297# 6.12e-19
C94 input5/a_664_47# net1 2.41e-19
C95 _10_ _03_ 0.00244f
C96 net13 _33_/a_368_53# 2.1e-20
C97 _15_ _27_/a_205_297# 5.5e-20
C98 _42_/a_209_311# net6 1.32e-20
C99 _36_/a_109_47# _06_ 0.00168f
C100 _33_/a_109_93# _52_/a_250_297# 5.17e-22
C101 net13 net6 0.00188f
C102 _14_ _26_/a_183_297# 6.98e-22
C103 _25_ net10 2.02e-19
C104 p[10] _27_/a_27_297# 6.35e-19
C105 input6/a_27_47# _17_ 7.13e-22
C106 _50_/a_223_47# _47_/a_299_297# 2.74e-20
C107 _38_/a_303_47# _12_ 0.00153f
C108 _50_/a_343_93# _47_/a_81_21# 0.00282f
C109 _38_/a_109_47# net4 7.32e-19
C110 input5/a_62_47# _19_ 0.00159f
C111 _50_/a_343_93# _18_ 0.0276f
C112 _11_ _47_/a_299_297# 0.00738f
C113 input12/a_27_47# net10 0.00182f
C114 net7 _31_/a_285_47# 0.00132f
C115 net11 net1 1.13e-19
C116 input10/a_27_47# net10 0.00321f
C117 net1 _35_/a_226_47# 1.3e-20
C118 _43_/a_193_413# _01_ 8.16e-19
C119 p[10] input2/a_27_47# 0.00924f
C120 _43_/a_469_47# net15 7.41e-19
C121 b[1] net8 0.00195f
C122 net1 _06_ 0.0115f
C123 p[3] _30_/a_215_297# 2.01e-19
C124 net2 _22_ 1.93e-20
C125 _12_ _05_ 2.52e-19
C126 _22_ net19 2.17e-19
C127 _36_/a_27_47# _05_ 3.67e-21
C128 _53_/a_29_53# _21_ 0.00959f
C129 _55_/a_300_47# _06_ 2.5e-20
C130 _12_ _45_/a_465_47# 0.00211f
C131 p[12] _18_ 3.95e-21
C132 _10_ _41_/a_145_75# 5.18e-19
C133 input14/a_27_47# p[8] 0.0159f
C134 _32_/a_27_47# p[13] 6.49e-20
C135 _09_ _05_ 0.0683f
C136 _22_ _45_/a_193_297# 0.0234f
C137 _53_/a_111_297# _10_ 2.06e-19
C138 net6 _30_/a_215_297# 3.3e-21
C139 VPWR _42_/a_296_53# -6.37e-20
C140 p[2] _49_/a_75_199# 1.06e-19
C141 net13 input9/a_75_212# 4.4e-19
C142 net12 p[4] 5.33e-19
C143 _10_ _30_/a_297_297# 1.25e-20
C144 _09_ _45_/a_465_47# 2.77e-19
C145 _50_/a_343_93# _10_ 0.0284f
C146 net15 _49_/a_75_199# 5.13e-20
C147 _44_/a_256_47# net14 0.00379f
C148 _14_ p[14] 1.66e-20
C149 _37_/a_303_47# VPWR -3.13e-19
C150 _39_/a_47_47# _03_ 1.47e-19
C151 _01_ _31_/a_35_297# 4.27e-19
C152 _55_/a_217_297# _10_ 1.43e-19
C153 _12_ net5 0.983f
C154 _14_ net5 3.89e-19
C155 _36_/a_27_47# net5 0.0163f
C156 net11 net16 4.43e-22
C157 _38_/a_109_47# VPWR -4.66e-19
C158 p[1] net2 5.99e-20
C159 input3/a_27_47# _42_/a_109_93# 0.00249f
C160 _09_ net5 5.18e-19
C161 _42_/a_209_311# _20_ 1.66e-20
C162 _53_/a_29_53# _02_ 0.0388f
C163 net1 net3 4.25e-20
C164 VPWR net17 0.0371f
C165 net13 _20_ 5.95e-19
C166 net14 _03_ 1.5e-19
C167 VPWR _44_/a_584_47# -2.28e-19
C168 net12 _50_/a_27_47# 7.99e-21
C169 net16 _06_ 0.0511f
C170 VPWR _27_/a_277_297# -3.63e-19
C171 input5/a_558_47# net8 0.00357f
C172 net10 _05_ 0.457f
C173 _24_ b[2] 1.85e-19
C174 p[12] _10_ 0.0993f
C175 _49_/a_315_47# _03_ 9.22e-19
C176 _34_/a_285_47# net10 0.0454f
C177 _22_ b[2] 0.0043f
C178 input5/a_664_47# p[13] 8.06e-19
C179 input14/a_27_47# net3 9.36e-19
C180 p[7] net9 8.26e-19
C181 _15_ _43_/a_27_47# 8.96e-20
C182 net18 _38_/a_27_47# 0.00997f
C183 input9/a_75_212# _30_/a_215_297# 6.24e-21
C184 net10 net5 0.0316f
C185 _42_/a_209_311# _18_ 3.21e-19
C186 net7 net1 0.0712f
C187 net13 _18_ 1.06e-20
C188 _11_ p[9] 1.01e-19
C189 p[5] VPWR 0.092f
C190 p[8] p[13] 0.00172f
C191 _03_ _34_/a_377_297# 3.13e-20
C192 net11 _23_ 0.0461f
C193 _19_ _31_/a_285_297# 1.34e-19
C194 _27_/a_27_297# _03_ 2.68e-19
C195 _52_/a_250_297# _35_/a_76_199# 3.4e-21
C196 net13 _07_ 0.00686f
C197 _20_ _30_/a_215_297# 6.08e-19
C198 net12 _29_/a_29_53# 0.0132f
C199 _50_/a_27_47# _29_/a_29_53# 1.44e-20
C200 _35_/a_226_47# _23_ 4.21e-19
C201 _37_/a_27_47# VPWR -0.0178f
C202 VPWR _40_/a_109_297# -4.23e-19
C203 b[3] _14_ 1.92e-19
C204 _23_ _06_ 0.218f
C205 _11_ _39_/a_377_297# 2.57e-20
C206 _43_/a_27_47# net6 9.07e-20
C207 _21_ _24_ 0.0388f
C208 _33_/a_109_93# _35_/a_76_199# 3.08e-19
C209 _21_ _22_ 0.00314f
C210 _11_ _41_/a_59_75# 8.7e-19
C211 net9 _03_ 0.15f
C212 _21_ p[6] 0.00203f
C213 _50_/a_343_93# net14 1.07e-20
C214 _38_/a_197_47# _06_ 4.32e-19
C215 input2/a_27_47# _03_ 2.71e-19
C216 _55_/a_217_297# net14 2.1e-19
C217 _55_/a_80_21# _01_ 0.0121f
C218 p[12] output19/a_27_47# 1.78e-19
C219 _39_/a_47_47# p[12] 3.32e-19
C220 net13 _10_ 0.00151f
C221 _15_ _12_ 0.00833f
C222 _08_ _34_/a_129_47# 3.29e-19
C223 _49_/a_75_199# _29_/a_29_53# 1.28e-19
C224 _42_/a_368_53# net3 3.82e-19
C225 _15_ _14_ 0.148f
C226 _04_ _22_ 1.76e-20
C227 net19 net8 1.15e-19
C228 net2 net8 0.0525f
C229 _26_/a_29_53# _03_ 7.93e-21
C230 _38_/a_27_47# _10_ 0.0133f
C231 _24_ _02_ 0.023f
C232 net3 p[13] 3.65e-19
C233 b[3] _55_/a_472_297# 1.51e-19
C234 _22_ _02_ 0.552f
C235 input12/a_27_47# p[5] 0.00359f
C236 _14_ _19_ 2.71e-21
C237 p[5] input10/a_27_47# 0.0172f
C238 _19_ _09_ 4.8e-21
C239 _37_/a_27_47# _00_ 6.15e-20
C240 net6 _12_ 0.0891f
C241 input13/a_27_47# p[7] 0.0167f
C242 net17 _05_ 0.0111f
C243 net6 _36_/a_27_47# 5.1e-19
C244 _15_ _50_/a_429_93# 6.82e-19
C245 _11_ _45_/a_27_47# 0.0703f
C246 _14_ net6 2.11e-19
C247 p[1] _04_ 1.74e-21
C248 VPWR _31_/a_285_47# -2.91e-19
C249 _35_/a_556_47# VPWR -7.24e-19
C250 net10 _34_/a_47_47# 0.0507f
C251 _15_ _55_/a_472_297# 0.00626f
C252 _50_/a_343_93# _17_ 0.0015f
C253 net6 _09_ 5.43e-20
C254 _40_/a_191_297# _06_ 5.84e-19
C255 p[11] _37_/a_197_47# 1.59e-19
C256 _44_/a_93_21# _43_/a_193_413# 0.0161f
C257 net7 p[13] 1.91e-19
C258 net9 _30_/a_297_297# 7.83e-19
C259 net9 _50_/a_343_93# 6.64e-19
C260 _10_ _30_/a_215_297# 5.66e-20
C261 _53_/a_29_53# net11 8.31e-19
C262 _43_/a_27_47# _20_ 0.0124f
C263 net5 net17 4.21e-21
C264 _53_/a_29_53# _06_ 0.0709f
C265 p[3] net10 8.58e-19
C266 _16_ _43_/a_193_413# 0.0261f
C267 _52_/a_250_297# b[2] 1.6e-19
C268 net2 b[1] 0.0191f
C269 _50_/a_429_93# net6 6.18e-19
C270 _49_/a_201_297# _31_/a_35_297# 5.52e-20
C271 _43_/a_193_413# net15 0.00169f
C272 _33_/a_368_53# net10 0.00171f
C273 p[11] input5/a_62_47# 0.00153f
C274 _44_/a_93_21# _44_/a_250_297# -6.97e-22
C275 _50_/a_343_93# _26_/a_29_53# 2.61e-19
C276 input6/a_27_47# p[9] 0.0762f
C277 input5/a_381_47# _06_ 1.6e-19
C278 _42_/a_209_311# net14 0.0238f
C279 _22_ _32_/a_27_47# 1.76e-19
C280 _53_/a_29_53# _48_/a_27_47# 3.14e-21
C281 net10 net6 1.35e-20
C282 net13 net14 2.21e-21
C283 _40_/a_191_297# net3 1.89e-19
C284 _37_/a_197_47# net14 7e-19
C285 net2 _40_/a_297_297# 0.00101f
C286 VPWR _36_/a_109_47# -4.66e-19
C287 _44_/a_250_297# _16_ 3.25e-19
C288 _43_/a_27_47# _18_ 0.0201f
C289 p[1] input7/a_27_47# 0.0164f
C290 p[2] _31_/a_35_297# 0.00264f
C291 _44_/a_250_297# net15 8.86e-20
C292 _52_/a_93_21# _23_ 0.0166f
C293 _37_/a_27_47# p[14] 1.37e-19
C294 _49_/a_544_297# _03_ 0.00568f
C295 _20_ _12_ 3.9e-19
C296 _20_ _36_/a_27_47# 0.00148f
C297 _37_/a_27_47# net5 1.13e-20
C298 _14_ _20_ 0.144f
C299 _27_/a_205_297# net14 3.63e-19
C300 _21_ net8 0.00656f
C301 _20_ _09_ 7.11e-19
C302 net4 net16 0.155f
C303 VPWR _30_/a_465_297# -4.57e-19
C304 input5/a_558_47# net2 5.99e-21
C305 input5/a_558_47# net19 2.24e-20
C306 input5/a_381_47# net3 0.0299f
C307 input5/a_62_47# net14 5.28e-20
C308 net18 _12_ 8.24e-19
C309 _25_ _36_/a_109_47# 3.76e-21
C310 _13_ net16 0.0198f
C311 p[10] _01_ 7.94e-20
C312 _42_/a_209_311# _27_/a_27_297# 4.7e-20
C313 _15_ _42_/a_296_53# 1.28e-19
C314 net1 VPWR 1.17f
C315 input9/a_75_212# net10 0.00699f
C316 _04_ net8 0.02f
C317 _17_ _42_/a_209_311# 1.22e-19
C318 b[3] _44_/a_584_47# 0.00109f
C319 _10_ _43_/a_27_47# 0.0279f
C320 net18 _09_ 1.97e-21
C321 _04_ _52_/a_250_297# 3.98e-21
C322 _33_/a_109_93# _21_ 1.62e-20
C323 _55_/a_300_47# VPWR -4.61e-19
C324 _44_/a_346_47# _10_ 9.13e-21
C325 _47_/a_81_21# _12_ 0.00158f
C326 _37_/a_197_47# _17_ 9.19e-21
C327 _47_/a_81_21# _14_ 6.24e-20
C328 _02_ net8 0.334f
C329 _18_ _12_ 0.0115f
C330 net13 net9 0.035f
C331 net11 _22_ 6.82e-21
C332 _18_ _36_/a_27_47# 5.46e-20
C333 _55_/a_472_297# _20_ 0.00212f
C334 _52_/a_250_297# _02_ 0.0128f
C335 input14/a_27_47# VPWR 0.0735f
C336 net11 p[6] 0.0099f
C337 input2/a_27_47# _42_/a_209_311# 1e-22
C338 _14_ _18_ 0.243f
C339 net10 _20_ 3.23e-19
C340 p[1] input5/a_664_47# 1.21e-20
C341 net7 input5/a_381_47# 4.91e-19
C342 _33_/a_109_93# _04_ 0.0299f
C343 _22_ _35_/a_226_47# 1.39e-20
C344 _12_ _07_ 2.94e-23
C345 _18_ _09_ 7.01e-21
C346 _24_ _06_ 0.113f
C347 _05_ _31_/a_285_47# 5.61e-19
C348 p[6] _06_ 2.62e-19
C349 _22_ _06_ 0.124f
C350 _19_ net17 0.0211f
C351 _09_ _07_ 0.0405f
C352 _33_/a_109_93# _02_ 1.54e-21
C353 _22_ _26_/a_111_297# 0.00137f
C354 net13 _26_/a_29_53# 2.23e-20
C355 _11_ _44_/a_93_21# 4.78e-20
C356 VPWR net16 0.518f
C357 net1 _00_ 9.43e-19
C358 _13_ _23_ 2.08e-20
C359 input12/a_27_47# net1 7.44e-20
C360 p[6] _48_/a_27_47# 2.22e-19
C361 _55_/a_80_21# _16_ 0.0143f
C362 _11_ _16_ 4.42e-20
C363 net9 input5/a_62_47# 3.12e-19
C364 _38_/a_197_47# net4 7.64e-19
C365 _11_ _47_/a_384_47# 7.23e-20
C366 _10_ _12_ 0.19f
C367 input7/a_27_47# net8 2.03e-21
C368 _04_ b[1] 5.79e-19
C369 _14_ _10_ 0.0571f
C370 _36_/a_197_47# _06_ 6.18e-19
C371 _10_ _36_/a_27_47# 0.00109f
C372 _53_/a_29_53# _52_/a_93_21# 0.00116f
C373 net10 _18_ 1.47e-21
C374 _55_/a_80_21# net15 0.00759f
C375 _49_/a_75_199# _31_/a_35_297# 6.24e-19
C376 _10_ _09_ 0.0222f
C377 net9 _30_/a_215_297# 0.0458f
C378 _22_ net3 9.39e-20
C379 _11_ net15 0.145f
C380 net10 _07_ 0.057f
C381 net2 net19 0.599f
C382 input2/a_27_47# _30_/a_215_297# 3.51e-20
C383 _29_/a_183_297# _03_ 7.36e-19
C384 _32_/a_27_47# net8 0.0275f
C385 _37_/a_27_47# _15_ 1.11e-19
C386 _25_ net16 1.16e-19
C387 _53_/a_183_297# _10_ 2.86e-19
C388 _43_/a_27_47# net14 4.87e-20
C389 VPWR _42_/a_368_53# -3.03e-19
C390 input8/a_27_47# net1 0.0347f
C391 net12 _08_ 0.0269f
C392 _14_ _43_/a_297_47# 9.11e-19
C393 _50_/a_429_93# _10_ 0.00167f
C394 _44_/a_346_47# net14 0.00464f
C395 VPWR p[13] 0.183f
C396 _55_/a_472_297# _10_ 7.35e-21
C397 _36_/a_109_47# net5 0.00144f
C398 VPWR _23_ -0.00374f
C399 _10_ net10 4.45e-19
C400 p[11] _14_ 7.85e-20
C401 input3/a_27_47# _42_/a_209_311# 1.56e-19
C402 net13 input13/a_27_47# 0.00139f
C403 net7 _22_ 2.73e-20
C404 _39_/a_129_47# b[0] 2.6e-20
C405 _38_/a_197_47# VPWR -5.24e-19
C406 _37_/a_27_47# net6 4.3e-20
C407 _40_/a_109_297# net6 2.53e-20
C408 input5/a_558_47# _04_ 1.25e-20
C409 net1 _05_ 0.151f
C410 net12 _30_/a_109_53# 4.25e-20
C411 _16_ _28_/a_109_297# 1.26e-19
C412 _01_ _03_ 2.85e-19
C413 _50_/a_27_47# _50_/a_223_47# 5.68e-32
C414 input5/a_664_47# net8 0.0116f
C415 _39_/a_47_47# _12_ 0.0317f
C416 _14_ output19/a_27_47# 1.43e-19
C417 _44_/a_93_21# _42_/a_109_93# 1.25e-19
C418 net12 _11_ 3.82e-21
C419 _11_ _50_/a_27_47# 0.0592f
C420 _03_ _49_/a_208_47# 3.86e-19
C421 _21_ _35_/a_76_199# 0.0175f
C422 _53_/a_29_53# net4 3.26e-19
C423 _20_ net17 4e-20
C424 _35_/a_489_413# _45_/a_27_47# 3.89e-21
C425 _25_ _23_ 0.00465f
C426 _38_/a_303_47# net16 6.47e-19
C427 _39_/a_47_47# _09_ 7.7e-21
C428 _53_/a_29_53# _13_ 9.05e-19
C429 net13 _49_/a_544_297# 3.43e-19
C430 net1 net5 0.0772f
C431 p[1] net7 0.00514f
C432 _17_ _43_/a_27_47# 0.00131f
C433 _04_ _35_/a_76_199# 0.0269f
C434 _44_/a_346_47# _17_ 7.2e-19
C435 input3/a_27_47# input5/a_62_47# 0.00179f
C436 _14_ net14 0.184f
C437 net11 net8 1.5e-19
C438 _16_ input5/a_841_47# 8.62e-19
C439 _45_/a_27_47# _03_ 2.06e-20
C440 net11 _52_/a_250_297# 1.2e-19
C441 _42_/a_109_93# net15 4.62e-19
C442 _52_/a_93_21# _24_ 0.0211f
C443 _52_/a_250_297# _35_/a_226_47# 2.63e-20
C444 _06_ net8 0.00282f
C445 _22_ _52_/a_93_21# 0.0347f
C446 _35_/a_76_199# _02_ 5.73e-19
C447 _49_/a_315_47# _09_ 1.11e-20
C448 net12 _29_/a_111_297# 1.21e-19
C449 _29_/a_29_53# _30_/a_109_53# 0.0103f
C450 net15 input5/a_841_47# 0.00585f
C451 _50_/a_223_47# _29_/a_29_53# 1.45e-20
C452 _52_/a_250_297# _06_ 0.0058f
C453 input6/a_27_47# _44_/a_93_21# 8.53e-19
C454 p[12] input4/a_75_212# 0.02f
C455 p[12] p[9] 1.4e-19
C456 _39_/a_47_47# net10 4.72e-22
C457 VPWR _40_/a_191_297# -6.82e-19
C458 _50_/a_343_93# _41_/a_59_75# 6.13e-22
C459 input7/a_27_47# input5/a_558_47# 1.22e-20
C460 net11 _33_/a_109_93# 5.14e-19
C461 _33_/a_109_93# _35_/a_226_47# 4.9e-19
C462 _33_/a_209_311# _35_/a_76_199# 9.95e-21
C463 _50_/a_429_93# net14 6.04e-21
C464 _50_/a_343_93# _01_ 0.0131f
C465 _55_/a_217_297# _01_ 0.00112f
C466 _33_/a_109_93# _06_ 9.13e-19
C467 _53_/a_29_53# VPWR 0.00821f
C468 net16 net5 0.00461f
C469 _40_/a_109_297# _20_ 2.35e-20
C470 p[5] net18 1.98e-19
C471 _04_ net19 2.07e-20
C472 net2 _04_ 0.158f
C473 _14_ _27_/a_27_297# 1.66e-21
C474 input6/a_27_47# net15 0.00115f
C475 _17_ _12_ 0.0109f
C476 p[12] _41_/a_59_75# 0.0547f
C477 _14_ _17_ 0.489f
C478 net3 net8 9.23e-19
C479 p[10] net15 0.01f
C480 _54_/a_75_212# _02_ 6.6e-20
C481 input5/a_381_47# VPWR 8.33e-19
C482 _38_/a_109_47# _10_ 5.44e-19
C483 net9 _12_ 4.39e-22
C484 net19 _02_ 0.0474f
C485 net9 _36_/a_27_47# 0.00493f
C486 _10_ _44_/a_584_47# 1.14e-20
C487 net9 _09_ 2.62e-19
C488 _02_ _45_/a_193_297# 0.00988f
C489 _53_/a_29_53# _25_ 0.00146f
C490 _11_ _45_/a_109_297# 0.00168f
C491 net4 _24_ 8.65e-20
C492 _37_/a_27_47# _18_ 3.31e-20
C493 b[3] input14/a_27_47# 0.0211f
C494 net10 _34_/a_377_297# 1.62e-19
C495 _22_ net4 0.0866f
C496 _21_ b[2] 2.14e-19
C497 _42_/a_209_311# p[9] 5.51e-21
C498 _13_ _24_ 2.47e-19
C499 _26_/a_29_53# _12_ 0.00243f
C500 p[11] _37_/a_303_47# 1.04e-19
C501 net5 p[13] 0.0069f
C502 _26_/a_29_53# _36_/a_27_47# 1.6e-19
C503 _13_ _22_ 0.00309f
C504 _40_/a_297_297# _06_ 1.64e-19
C505 net7 net8 0.295f
C506 _14_ _26_/a_29_53# 3.67e-19
C507 _23_ net5 0.0052f
C508 net9 _30_/a_392_297# 9.92e-19
C509 _55_/a_300_47# _15_ 1.42e-20
C510 net1 _19_ 2.86e-19
C511 p[3] net1 6.54e-19
C512 input7/a_27_47# net2 3.24e-19
C513 net9 net10 0.111f
C514 output16/a_27_47# net4 0.00706f
C515 input2/a_27_47# net10 1.17e-20
C516 _02_ b[2] 2.69e-19
C517 _13_ output16/a_27_47# 4.58e-19
C518 _44_/a_93_21# _44_/a_256_47# -6.6e-20
C519 input5/a_558_47# _06_ 3.55e-19
C520 _42_/a_296_53# net14 2.18e-19
C521 _42_/a_209_311# _01_ 1.58e-19
C522 net13 _01_ 0.00228f
C523 VPWR _24_ 0.0129f
C524 _40_/a_297_297# net3 2.54e-19
C525 _26_/a_29_53# net10 3.48e-22
C526 _49_/a_201_297# _03_ 0.00842f
C527 _37_/a_303_47# net14 0.00112f
C528 VPWR _22_ 1.4f
C529 VPWR p[6] 0.0738f
C530 p[10] _49_/a_75_199# 2.29e-20
C531 _52_/a_93_21# _52_/a_250_297# -6.97e-22
C532 net7 b[1] 0.005f
C533 net11 _35_/a_76_199# 4e-19
C534 net14 net17 5.43e-19
C535 _21_ _04_ 0.39f
C536 _35_/a_556_47# _07_ 0.00128f
C537 _44_/a_584_47# net14 7.2e-19
C538 b[3] p[13] 0.165f
C539 _35_/a_76_199# _06_ 0.00425f
C540 input13/a_27_47# _09_ 1.27e-21
C541 p[7] p[4] 7.8e-20
C542 p[11] _37_/a_27_47# 4.41e-19
C543 _27_/a_277_297# net14 5.1e-19
C544 VPWR _36_/a_197_47# -5.24e-19
C545 _33_/a_109_93# _52_/a_93_21# 2.89e-21
C546 input5/a_558_47# net3 0.0137f
C547 _21_ _02_ 0.397f
C548 net6 net16 8.27e-20
C549 VPWR output16/a_27_47# 0.122f
C550 input5/a_664_47# net19 1.38e-21
C551 input5/a_664_47# net2 8.11e-20
C552 p[1] VPWR 0.08f
C553 input9/a_75_212# net1 0.002f
C554 net15 _03_ 4.26e-20
C555 _25_ _22_ 5.39e-19
C556 _04_ _02_ 0.0541f
C557 _42_/a_109_93# output17/a_27_47# 8.6e-21
C558 _55_/a_80_21# _43_/a_193_413# 2.54e-19
C559 net12 p[7] 0.0343f
C560 _37_/a_303_47# _17_ 1.23e-20
C561 _22_ _00_ 0.477f
C562 _11_ _43_/a_193_413# 5.45e-19
C563 _47_/a_299_297# _12_ 0.00805f
C564 net11 _54_/a_75_212# 0.00956f
C565 _49_/a_544_297# _09_ 2.56e-20
C566 input12/a_27_47# p[6] 0.0166f
C567 _27_/a_27_297# net17 0.00181f
C568 input5/a_381_47# net5 0.0546f
C569 input13/a_27_47# net10 8.86e-20
C570 net1 _20_ 0.363f
C571 _52_/a_256_47# _02_ 0.00344f
C572 input10/a_27_47# p[6] 0.00214f
C573 _54_/a_75_212# _06_ 0.00727f
C574 net19 p[8] 0.0268f
C575 net2 p[8] 0.00102f
C576 _33_/a_209_311# _04_ 0.00133f
C577 net7 input5/a_558_47# 0.00358f
C578 _25_ _36_/a_197_47# 2.37e-21
C579 _37_/a_27_47# net14 0.0584f
C580 net2 _06_ 0.0108f
C581 net19 _06_ 0.00522f
C582 _30_/a_109_53# _31_/a_35_297# 2.89e-20
C583 _35_/a_226_47# _45_/a_193_297# 8.15e-21
C584 _35_/a_489_413# net12 3.97e-20
C585 _55_/a_80_21# _31_/a_35_297# 5.9e-21
C586 net4 _52_/a_250_297# 0.00136f
C587 _22_ _26_/a_183_297# 0.00184f
C588 net9 net17 1.26e-20
C589 _45_/a_193_297# _06_ 0.00201f
C590 p[0] input1/a_75_212# 0.0172f
C591 input2/a_27_47# net17 0.0398f
C592 net6 _23_ 2.13e-19
C593 net11 _36_/a_303_47# 7.63e-20
C594 _13_ _52_/a_250_297# 5.43e-19
C595 p[10] output17/a_27_47# 0.118f
C596 net12 _03_ 0.0268f
C597 _55_/a_217_297# _16_ 0.0017f
C598 net1 _47_/a_81_21# 1.58e-21
C599 _21_ _32_/a_27_47# 8.95e-19
C600 net7 _35_/a_76_199# 1.79e-20
C601 _36_/a_303_47# _06_ 5.3e-19
C602 _55_/a_217_297# net15 7.79e-19
C603 net1 _07_ 6.08e-22
C604 _04_ _32_/a_27_47# 1.43e-19
C605 net11 b[2] 1.46e-19
C606 net19 net3 0.611f
C607 net2 net3 0.519f
C608 _22_ _05_ 3.33e-21
C609 net18 net16 0.00585f
C610 _49_/a_75_199# _03_ 0.0849f
C611 b[2] _06_ 0.0116f
C612 _40_/a_109_297# _17_ 9.67e-19
C613 _37_/a_27_47# _17_ 0.00277f
C614 _34_/a_285_47# p[6] 8.31e-20
C615 _32_/a_27_47# _02_ 0.00247f
C616 input8/a_27_47# p[1] 5.13e-20
C617 _43_/a_27_47# _01_ 9.77e-20
C618 _53_/a_29_53# _34_/a_47_47# 5.88e-22
C619 VPWR net8 0.703f
C620 p[12] net15 2.99e-19
C621 _14_ _43_/a_369_47# 0.00135f
C622 VPWR _52_/a_250_297# 0.019f
C623 _01_ _31_/a_285_297# 1.92e-19
C624 input5/a_664_47# _21_ 9.42e-22
C625 _24_ net5 5.83e-20
C626 _03_ _29_/a_29_53# 0.0414f
C627 net1 _10_ 4.34e-19
C628 input4/a_75_212# _12_ 2.09e-20
C629 _22_ net5 0.405f
C630 _27_/a_109_297# _03_ 1.97e-20
C631 _18_ net16 8.17e-21
C632 net2 input15/a_27_47# 0.00296f
C633 _14_ p[9] 2.62e-21
C634 net19 input15/a_27_47# 0.00236f
C635 p[5] input11/a_27_47# 0.0433f
C636 net7 net2 0.00234f
C637 _52_/a_93_21# _35_/a_76_199# 6.83e-21
C638 _39_/a_285_47# b[0] 1.88e-19
C639 input5/a_664_47# _04_ 6.73e-21
C640 _33_/a_109_93# VPWR -0.00817f
C641 _40_/a_191_297# net6 1.16e-20
C642 _29_/a_183_297# _09_ 4.51e-20
C643 net12 _30_/a_297_297# 7.14e-21
C644 net13 _49_/a_201_297# 3.31e-19
C645 _39_/a_377_297# _12_ 6.77e-19
C646 net11 _21_ 0.586f
C647 _44_/a_250_297# _42_/a_109_93# 6.38e-19
C648 _44_/a_93_21# _42_/a_209_311# 2.21e-19
C649 input5/a_664_47# _02_ 0.00187f
C650 _11_ _50_/a_223_47# 0.0329f
C651 output16/a_27_47# net5 4.08e-20
C652 _21_ _35_/a_226_47# 9.87e-19
C653 _36_/a_197_47# net5 0.00254f
C654 _53_/a_29_53# net6 2.11e-20
C655 _41_/a_59_75# _12_ 0.00101f
C656 _21_ _06_ 0.143f
C657 net11 _04_ 0.078f
C658 _16_ _42_/a_209_311# 0.00129f
C659 _00_ net8 3.23e-19
C660 _10_ net16 0.0338f
C661 _50_/a_27_47# p[12] 1.34e-19
C662 VPWR b[1] 0.396f
C663 _04_ _35_/a_226_47# 0.00551f
C664 _14_ _01_ 0.0193f
C665 _21_ _48_/a_27_47# 0.0121f
C666 _01_ _09_ 4.69e-21
C667 _04_ _06_ 0.0136f
C668 _42_/a_209_311# net15 0.0157f
C669 net11 _02_ 0.0327f
C670 net13 net15 8.84e-19
C671 _37_/a_197_47# net15 1.78e-19
C672 p[11] input14/a_27_47# 0.00118f
C673 _35_/a_226_47# _02_ 2.21e-19
C674 input5/a_62_47# _44_/a_93_21# 5.05e-20
C675 _52_/a_256_47# _06_ 0.00157f
C676 VPWR _40_/a_297_297# -5.42e-19
C677 _02_ _06_ 0.85f
C678 _03_ output17/a_27_47# 1.95e-19
C679 _49_/a_208_47# _09_ 5.43e-21
C680 _23_ _07_ 1.27e-19
C681 b[3] _22_ 1.28e-19
C682 _52_/a_93_21# _45_/a_193_297# 6.01e-19
C683 input13/a_27_47# p[5] 3.09e-19
C684 input7/a_27_47# input5/a_664_47# 1.08e-21
C685 net11 _33_/a_209_311# 2.49e-19
C686 p[10] _31_/a_35_297# 2.29e-19
C687 _33_/a_209_311# _35_/a_226_47# 1.31e-19
C688 _45_/a_27_47# _12_ 0.0866f
C689 _02_ _48_/a_27_47# 0.00435f
C690 _33_/a_209_311# _06_ 0.0187f
C691 input14/a_27_47# output19/a_27_47# 0.0101f
C692 input8/a_27_47# net8 0.0181f
C693 net1 net14 6.64e-20
C694 _55_/a_472_297# _01_ 6.28e-19
C695 _24_ _34_/a_47_47# 6.84e-21
C696 _40_/a_191_297# _20_ 2.07e-20
C697 net13 p[4] 2.34e-20
C698 _22_ _34_/a_47_47# 3.9e-21
C699 _55_/a_80_21# _28_/a_109_297# 2.05e-20
C700 _13_ _35_/a_76_199# 3.01e-21
C701 _45_/a_27_47# _09_ 0.00823f
C702 p[6] _34_/a_47_47# 4.28e-19
C703 _50_/a_515_93# _06_ 0.00244f
C704 _04_ net3 0.113f
C705 _11_ _28_/a_109_297# 6.29e-19
C706 _15_ _22_ 0.0236f
C707 _10_ _23_ 0.00192f
C708 input5/a_558_47# VPWR 0.0083f
C709 input14/a_27_47# net14 0.0232f
C710 net3 _02_ 9.52e-20
C711 _22_ _52_/a_584_47# 6.24e-19
C712 net8 _05_ 0.0146f
C713 _52_/a_250_297# _05_ 8.86e-22
C714 _52_/a_93_21# b[2] 1.63e-19
C715 _38_/a_197_47# _10_ 6.29e-19
C716 _39_/a_47_47# net16 7.7e-20
C717 net7 _21_ 3e-19
C718 net13 net12 0.363f
C719 net13 _50_/a_27_47# 7.27e-21
C720 _53_/a_29_53# net18 0.0118f
C721 net6 _24_ 0.00121f
C722 _50_/a_27_47# _38_/a_27_47# 2.37e-20
C723 net1 _27_/a_27_297# 6.05e-21
C724 net7 _04_ 0.0602f
C725 _33_/a_109_93# _05_ 0.0206f
C726 net10 _34_/a_129_47# 0.003f
C727 _32_/a_27_47# _06_ 0.00663f
C728 net19 net4 2.65e-20
C729 net5 net8 0.48f
C730 _22_ net6 0.163f
C731 VPWR _35_/a_76_199# -0.00947f
C732 _52_/a_250_297# net5 0.018f
C733 p[11] p[13] 0.00897f
C734 net4 _45_/a_193_297# 7.41e-19
C735 p[1] _19_ 2.82e-20
C736 net9 _30_/a_465_297# 0.00138f
C737 net13 _49_/a_75_199# 3.2e-19
C738 net7 _02_ 0.445f
C739 net9 net1 0.47f
C740 _38_/a_27_47# output18/a_27_47# 8.6e-19
C741 input2/a_27_47# net1 4.81e-19
C742 _36_/a_197_47# net6 6.94e-20
C743 output16/a_27_47# net6 1.5e-19
C744 net13 _29_/a_29_53# 0.00104f
C745 _39_/a_47_47# _23_ 5.24e-21
C746 _21_ _52_/a_93_21# 9.4e-19
C747 b[1] _05_ 5.29e-20
C748 net12 _30_/a_215_297# 0.00676f
C749 _44_/a_93_21# _44_/a_346_47# -5.12e-20
C750 input5/a_664_47# _06_ 3.21e-19
C751 _42_/a_368_53# net14 7.39e-19
C752 _54_/a_75_212# VPWR 0.0475f
C753 net14 p[13] 1.91e-19
C754 _04_ _52_/a_93_21# 2.35e-19
C755 _16_ _43_/a_27_47# 2.47e-19
C756 _53_/a_29_53# _10_ 0.00779f
C757 net2 VPWR 0.918f
C758 VPWR net19 0.181f
C759 net7 input7/a_27_47# 0.00318f
C760 _03_ _31_/a_35_297# 0.00749f
C761 _52_/a_93_21# _52_/a_256_47# -6.6e-20
C762 VPWR _45_/a_193_297# -0.00859f
C763 _52_/a_93_21# _02_ 0.0957f
C764 p[2] _31_/a_285_297# 0.00156f
C765 _01_ net17 0.0988f
C766 net11 _35_/a_226_47# 3.21e-19
C767 net11 _06_ 0.546f
C768 net7 _32_/a_27_47# 0.00559f
C769 _22_ _20_ 0.183f
C770 _35_/a_226_47# _06_ 0.00487f
C771 _37_/a_27_47# p[9] 0.0117f
C772 _29_/a_29_53# _30_/a_215_297# 1.72e-19
C773 VPWR _36_/a_303_47# -4.83e-19
C774 input5/a_664_47# net3 0.00215f
C775 _14_ _49_/a_201_297# 4.76e-21
C776 _25_ _54_/a_75_212# 0.0247f
C777 net11 _48_/a_27_47# 0.0179f
C778 _26_/a_111_297# _06_ 9e-19
C779 net18 _24_ 5.57e-21
C780 _49_/a_201_297# _09_ 1.74e-20
C781 _44_/a_93_21# _14_ 0.04f
C782 net18 _22_ 1.68e-19
C783 _15_ net8 1.79e-19
C784 _48_/a_27_47# _06_ 0.0251f
C785 _35_/a_489_413# _08_ 5.56e-19
C786 _54_/a_75_212# input10/a_27_47# 1.17e-22
C787 _21_ net4 0.00535f
C788 VPWR b[2] 0.262f
C789 net2 _00_ 0.00732f
C790 _47_/a_384_47# _12_ 9.51e-20
C791 input13/a_27_47# net1 1.9e-19
C792 _14_ _16_ 0.0584f
C793 _47_/a_81_21# _22_ 7.25e-19
C794 p[3] net8 0.0015f
C795 _19_ net8 0.0322f
C796 input5/a_558_47# net5 0.0597f
C797 _52_/a_346_47# _02_ 0.00526f
C798 _21_ _13_ 1.69e-19
C799 _22_ _18_ 0.0211f
C800 _00_ _45_/a_193_297# 4.38e-20
C801 net3 p[8] 2.53e-19
C802 net9 _23_ 1.21e-19
C803 _03_ _08_ 0.0144f
C804 net9 p[13] 1.72e-19
C805 _24_ _07_ 5.67e-19
C806 _25_ _36_/a_303_47# 2.03e-21
C807 net15 _12_ 8.14e-21
C808 _35_/a_76_199# _05_ 0.00238f
C809 p[10] _42_/a_109_93# 1.82e-21
C810 net7 input5/a_664_47# 0.00199f
C811 _14_ net15 0.0538f
C812 net3 _06_ 0.0072f
C813 _22_ _07_ 1.19e-20
C814 p[6] _07_ 1.26e-19
C815 b[3] b[1] 6.12e-20
C816 _13_ _04_ 1.17e-21
C817 input3/a_27_47# input14/a_27_47# 5.08e-20
C818 net6 _52_/a_250_297# 0.00133f
C819 net4 _02_ 0.00376f
C820 net1 input1/a_75_212# 0.00208f
C821 input5/a_62_47# output17/a_27_47# 1.02e-19
C822 _03_ _30_/a_109_53# 0.0189f
C823 net1 _49_/a_544_297# 0.00175f
C824 _50_/a_223_47# _03_ 1.41e-21
C825 _13_ _02_ 0.0676f
C826 _25_ b[2] 0.0015f
C827 _55_/a_472_297# _16_ 3.71e-19
C828 _35_/a_76_199# net5 3.38e-19
C829 input15/a_27_47# p[8] 7.57e-19
C830 net11 net7 1.77e-19
C831 _10_ _24_ 0.00484f
C832 net7 _35_/a_226_47# 2.93e-20
C833 _22_ _10_ 0.0904f
C834 input15/a_27_47# _06_ 4.73e-19
C835 net7 _06_ 0.00447f
C836 _21_ VPWR 0.871f
C837 input5/a_381_47# net14 0.00479f
C838 net2 _05_ 4.03e-20
C839 net12 _12_ 7.94e-21
C840 _50_/a_27_47# _12_ 0.00354f
C841 net12 _36_/a_27_47# 0.0185f
C842 _04_ VPWR 0.456f
C843 _50_/a_27_47# _36_/a_27_47# 6.08e-19
C844 _40_/a_191_297# _17_ 4.35e-19
C845 _45_/a_193_297# _05_ 4.84e-22
C846 net12 _09_ 0.0374f
C847 _14_ _43_/a_469_47# 0.00259f
C848 _50_/a_27_47# _09_ 1.3e-19
C849 _10_ _36_/a_197_47# 1.54e-19
C850 net2 p[14] 1.38e-19
C851 VPWR _52_/a_256_47# -9.47e-19
C852 net19 p[14] 0.101f
C853 _01_ _31_/a_285_47# 3.36e-19
C854 _03_ _29_/a_111_297# 7.48e-19
C855 VPWR _02_ 0.33f
C856 net10 p[4] 0.00268f
C857 net19 net5 0.00124f
C858 _25_ _21_ 0.00164f
C859 net2 net5 0.0616f
C860 net11 _52_/a_93_21# 2.8e-19
C861 p[11] _22_ 3.13e-20
C862 net3 input15/a_27_47# 8.74e-20
C863 net7 net3 7.45e-20
C864 input5/a_381_47# _27_/a_27_297# 1.47e-19
C865 _52_/a_93_21# _35_/a_226_47# 4.89e-20
C866 _20_ net8 5.07e-19
C867 _40_/a_297_297# net6 7.47e-22
C868 _45_/a_193_297# net5 0.00935f
C869 _33_/a_209_311# VPWR -0.0131f
C870 net12 _30_/a_392_297# 2.19e-20
C871 input3/a_27_47# p[13] 0.00499f
C872 _15_ input5/a_558_47# 0.00166f
C873 _21_ _00_ 9.26e-20
C874 _52_/a_93_21# _06_ 0.0574f
C875 _14_ _49_/a_75_199# 6.79e-20
C876 input12/a_27_47# _21_ 2.32e-19
C877 _49_/a_75_199# _09_ 2.93e-19
C878 _50_/a_515_93# VPWR -5.03e-19
C879 _39_/a_129_47# _12_ 0.00175f
C880 _50_/a_27_47# net10 3.78e-21
C881 net12 net10 0.539f
C882 _11_ _50_/a_343_93# 0.0384f
C883 _55_/a_80_21# _55_/a_217_297# 1.42e-32
C884 _36_/a_303_47# net5 0.00256f
C885 _36_/a_27_47# _29_/a_29_53# 6.92e-20
C886 net13 _31_/a_35_297# 1.86e-20
C887 net9 input5/a_381_47# 3.4e-19
C888 _04_ _00_ 1.98e-20
C889 _25_ _02_ 0.0156f
C890 _09_ _29_/a_29_53# 0.00488f
C891 input7/a_27_47# VPWR 0.0768f
C892 input1/a_75_212# p[13] 4.16e-19
C893 _47_/a_81_21# net8 2.08e-21
C894 _00_ _02_ 0.0269f
C895 _18_ net8 1.15e-21
C896 _22_ net14 2.23e-19
C897 input12/a_27_47# _02_ 1.88e-19
C898 _18_ _52_/a_250_297# 1.77e-19
C899 net5 b[2] 7.33e-20
C900 _11_ p[12] 3.51e-21
C901 VPWR _32_/a_27_47# 0.0395f
C902 _37_/a_303_47# net15 0.00118f
C903 _52_/a_346_47# _06_ 0.0031f
C904 input14/a_27_47# p[9] 8.53e-21
C905 input5/a_62_47# _44_/a_250_297# 2.45e-20
C906 b[3] net19 0.0439f
C907 b[3] net2 0.311f
C908 net10 _29_/a_29_53# 1.77e-19
C909 input8/a_27_47# _04_ 2.36e-22
C910 net15 net17 5.19e-19
C911 net6 _35_/a_76_199# 4.6e-21
C912 _45_/a_109_297# _12_ 0.00587f
C913 p[1] net14 0.0025f
C914 _21_ _05_ 0.0104f
C915 _33_/a_296_53# _06_ 1.11e-20
C916 _30_/a_215_297# _31_/a_35_297# 6.37e-19
C917 _33_/a_109_93# _07_ 3.2e-19
C918 net1 _01_ 0.0509f
C919 net11 _13_ 2.34e-19
C920 _27_/a_277_297# net15 1.93e-19
C921 net13 _08_ 1.82e-19
C922 _34_/a_285_47# _21_ 6.94e-20
C923 _13_ _35_/a_226_47# 5.62e-21
C924 _40_/a_297_297# _20_ 9.18e-21
C925 net4 _06_ 0.281f
C926 input8/a_27_47# _02_ 5.08e-20
C927 p[10] _03_ 8.74e-20
C928 _10_ net8 5.86e-19
C929 p[6] _34_/a_377_297# 5.39e-19
C930 _50_/a_615_93# _06_ 0.00264f
C931 _55_/a_300_47# _01_ 0.00113f
C932 _10_ _52_/a_250_297# 0.00368f
C933 _13_ _06_ 0.00188f
C934 _15_ net19 0.166f
C935 _15_ net2 9.8e-19
C936 _04_ _05_ 0.0352f
C937 input5/a_664_47# VPWR 0.00488f
C938 _22_ _17_ 0.00334f
C939 _21_ net5 0.00784f
C940 _37_/a_27_47# _44_/a_93_21# 3.19e-19
C941 net2 _19_ 0.101f
C942 net9 _22_ 0.0023f
C943 _32_/a_27_47# _00_ 0.00228f
C944 net13 _30_/a_109_53# 1.05e-19
C945 _55_/a_80_21# _42_/a_209_311# 0.0175f
C946 _02_ _05_ 0.00163f
C947 _34_/a_285_47# _02_ 7.14e-19
C948 _37_/a_27_47# _16_ 2.07e-19
C949 _04_ net5 0.00476f
C950 net4 net3 9.28e-21
C951 p[1] _27_/a_27_297# 2.27e-19
C952 net19 net6 0.00352f
C953 net2 net6 0.00139f
C954 _33_/a_209_311# _05_ 0.0311f
C955 net1 _32_/a_197_47# 0.00142f
C956 net11 VPWR 0.996f
C957 _26_/a_29_53# _24_ 2.11e-20
C958 _37_/a_27_47# net15 0.0541f
C959 VPWR p[8] 0.208f
C960 net12 net17 2.11e-21
C961 input8/a_27_47# input7/a_27_47# 3.2e-20
C962 VPWR _35_/a_226_47# 0.00159f
C963 _40_/a_109_297# net15 0.0016f
C964 _02_ net5 0.233f
C965 p[0] output17/a_27_47# 0.00805f
C966 _22_ _26_/a_29_53# 0.09f
C967 _11_ _38_/a_27_47# 0.071f
C968 net6 _45_/a_193_297# 9.84e-20
C969 VPWR _06_ 1.4f
C970 net10 output17/a_27_47# 1.31e-20
C971 _13_ _45_/a_205_47# 7.51e-20
C972 VPWR _26_/a_111_297# -5.92e-20
C973 p[5] p[4] 0.385f
C974 p[1] input2/a_27_47# 0.0119f
C975 _20_ _35_/a_76_199# 3.21e-20
C976 VPWR _48_/a_27_47# 0.0158f
C977 _36_/a_303_47# net6 1.25e-19
C978 _49_/a_75_199# net17 0.00127f
C979 _45_/a_27_47# net16 8.68e-19
C980 net11 _25_ 0.0262f
C981 net14 net8 0.0516f
C982 _32_/a_27_47# _05_ 2.2e-20
C983 _25_ _06_ 0.144f
C984 _01_ p[13] 2.02e-20
C985 net12 p[5] 0.00294f
C986 input6/a_27_47# p[12] 2.78e-19
C987 VPWR net3 0.351f
C988 input12/a_27_47# net11 0.00246f
C989 _43_/a_193_413# _12_ 7.94e-22
C990 net11 input10/a_27_47# 0.112f
C991 _03_ _31_/a_117_297# 5.32e-19
C992 _35_/a_489_413# _03_ 0.0205f
C993 _14_ _43_/a_193_413# 0.0297f
C994 p[11] b[1] 1.84e-20
C995 _52_/a_93_21# _52_/a_346_47# -5.12e-20
C996 _00_ _06_ 0.1f
C997 _21_ _34_/a_47_47# 8.93e-19
C998 _18_ _35_/a_76_199# 6.82e-21
C999 VPWR _45_/a_205_47# -1.62e-19
C1000 input12/a_27_47# _06_ 5.3e-22
C1001 _26_/a_111_297# _00_ 3.7e-19
C1002 _15_ _21_ 1.13e-21
C1003 _32_/a_27_47# net5 0.0961f
C1004 input13/a_27_47# p[6] 1.07e-19
C1005 _35_/a_76_199# _07_ 0.00226f
C1006 b[3] _02_ 1.07e-19
C1007 input3/a_27_47# _22_ 5.13e-20
C1008 net19 _20_ 1.29e-19
C1009 net2 _20_ 8.83e-19
C1010 _04_ _34_/a_47_47# 1.17e-20
C1011 net18 _54_/a_75_212# 0.0143f
C1012 _52_/a_93_21# net4 7.93e-20
C1013 VPWR input15/a_27_47# 0.0113f
C1014 p[3] _21_ 3.95e-21
C1015 net11 _48_/a_109_47# 1.74e-19
C1016 net7 VPWR 0.784f
C1017 _26_/a_183_297# _06_ 3.16e-19
C1018 _15_ _04_ 3.61e-20
C1019 _32_/a_109_47# net8 0.0011f
C1020 _44_/a_250_297# _14_ 4.82e-19
C1021 _13_ _52_/a_93_21# 1.31e-19
C1022 _45_/a_27_47# _23_ 1.74e-19
C1023 _27_/a_27_297# net8 0.0108f
C1024 _02_ _34_/a_47_47# 1.09e-19
C1025 _04_ _52_/a_584_47# 2.5e-19
C1026 _48_/a_109_47# _06_ 9.47e-19
C1027 _17_ net8 4.52e-20
C1028 _04_ _19_ 0.356f
C1029 _15_ _02_ 0.101f
C1030 _21_ net6 2.92e-20
C1031 _00_ net3 2.12e-19
C1032 p[3] _04_ 8.93e-22
C1033 _10_ _35_/a_76_199# 7.19e-20
C1034 net2 _47_/a_81_21# 4.95e-19
C1035 _33_/a_209_311# _34_/a_47_47# 0.017f
C1036 net19 _18_ 4.89e-20
C1037 net9 net8 0.0605f
C1038 input5/a_664_47# net5 0.0536f
C1039 _52_/a_584_47# _02_ 0.00389f
C1040 net2 _18_ 0.00181f
C1041 _19_ _02_ 0.213f
C1042 input2/a_27_47# net8 0.0207f
C1043 net11 _05_ 2.76e-19
C1044 output17/a_27_47# net17 0.0149f
C1045 p[10] _42_/a_209_311# 2.37e-20
C1046 net1 _49_/a_201_297# 0.00304f
C1047 _35_/a_226_47# _05_ 0.0134f
C1048 _04_ net6 2.61e-20
C1049 b[0] _12_ 2.61e-20
C1050 _55_/a_80_21# _43_/a_27_47# 1.56e-19
C1051 _50_/a_515_93# _15_ 0.00147f
C1052 _06_ _05_ 0.00724f
C1053 _11_ _43_/a_27_47# 4.27e-19
C1054 _34_/a_285_47# _06_ 0.00598f
C1055 p[14] p[8] 0.226f
C1056 net6 _02_ 0.00427f
C1057 p[1] input1/a_75_212# 0.00231f
C1058 net10 _31_/a_35_297# 3.95e-20
C1059 net9 _33_/a_109_93# 0.00211f
C1060 net7 _00_ 8.12e-21
C1061 VPWR _52_/a_93_21# -0.00838f
C1062 net18 b[2] 0.0131f
C1063 net11 net5 0.0129f
C1064 _03_ _30_/a_297_297# 0.00117f
C1065 p[14] _06_ 1.04e-19
C1066 _34_/a_285_47# _48_/a_27_47# 6.66e-20
C1067 net5 _06_ 0.41f
C1068 p[2] net1 0.0269f
C1069 net2 _10_ 2.65e-19
C1070 net19 _10_ 0.00224f
C1071 input9/a_75_212# _21_ 1.17e-21
C1072 net1 net15 7.44e-20
C1073 input5/a_558_47# net14 0.0325f
C1074 _08_ _09_ 0.103f
C1075 input7/a_27_47# _19_ 3.12e-21
C1076 _50_/a_515_93# net6 4.7e-19
C1077 _13_ net4 0.212f
C1078 _15_ _32_/a_27_47# 1.19e-19
C1079 _10_ _45_/a_193_297# 0.0047f
C1080 _55_/a_300_47# net15 1.09e-19
C1081 _50_/a_223_47# _12_ 0.00327f
C1082 input9/a_75_212# _04_ 7.69e-22
C1083 input2/a_27_47# b[1] 8.55e-19
C1084 _50_/a_223_47# _36_/a_27_47# 1.27e-20
C1085 _21_ _20_ 0.191f
C1086 _10_ _36_/a_303_47# 4.09e-19
C1087 _55_/a_80_21# _14_ 0.0175f
C1088 input8/a_27_47# net7 1.47e-19
C1089 p[14] net3 0.00446f
C1090 _11_ _12_ 0.195f
C1091 VPWR _52_/a_346_47# -0.00109f
C1092 _11_ _14_ 0.0415f
C1093 net3 net5 0.0365f
C1094 net10 _08_ 0.189f
C1095 p[11] net2 0.0204f
C1096 p[11] net19 0.00646f
C1097 net18 _21_ 0.00215f
C1098 _11_ _09_ 0.0665f
C1099 _04_ _20_ 0.0677f
C1100 net13 p[7] 0.00809f
C1101 _33_/a_296_53# VPWR -1.15e-19
C1102 input5/a_558_47# _27_/a_27_297# 1.57e-19
C1103 net7 _05_ 0.0129f
C1104 _45_/a_205_47# net5 8.28e-20
C1105 _15_ input5/a_664_47# 9.15e-22
C1106 net12 _30_/a_465_297# 8.01e-20
C1107 _20_ _02_ 0.1f
C1108 VPWR net4 1.07f
C1109 input5/a_558_47# _17_ 2.13e-21
C1110 b[3] p[8] 0.226f
C1111 _50_/a_615_93# VPWR -5.34e-19
C1112 net12 net1 1.17e-19
C1113 p[14] input15/a_27_47# 6.15e-19
C1114 _39_/a_285_47# _12_ 0.0221f
C1115 _13_ VPWR 0.0804f
C1116 net10 _30_/a_109_53# 5.6e-20
C1117 net19 output19/a_27_47# 0.0279f
C1118 net2 output19/a_27_47# 0.00168f
C1119 b[3] _06_ 9.96e-21
C1120 input5/a_664_47# _19_ 2.19e-21
C1121 input13/a_27_47# _33_/a_109_93# 0.00348f
C1122 net13 _35_/a_489_413# 7.36e-20
C1123 net9 input5/a_558_47# 4.42e-19
C1124 p[12] _41_/a_145_75# 0.00339f
C1125 net18 _02_ 6.8e-20
C1126 input5/a_558_47# input2/a_27_47# 2.04e-20
C1127 net11 _34_/a_47_47# 0.0309f
C1128 _21_ _07_ 0.133f
C1129 _09_ _29_/a_111_297# 5.79e-20
C1130 net7 net5 0.195f
C1131 _22_ _41_/a_59_75# 6.24e-22
C1132 _39_/a_47_47# _45_/a_193_297# 1.4e-20
C1133 _04_ _18_ 1.94e-21
C1134 _22_ _01_ 0.15f
C1135 _34_/a_47_47# _06_ 0.0391f
C1136 net19 net14 0.148f
C1137 net2 net14 0.151f
C1138 _14_ _28_/a_109_297# 5.66e-19
C1139 net13 _03_ 0.271f
C1140 _47_/a_81_21# _02_ 1.59e-20
C1141 net17 _31_/a_35_297# 0.0514f
C1142 net1 _49_/a_75_199# 0.00799f
C1143 _04_ _07_ 9.74e-20
C1144 _15_ _06_ 0.22f
C1145 net11 _19_ 6.27e-21
C1146 _18_ _02_ 2.96e-20
C1147 net15 p[13] 1.48e-19
C1148 _52_/a_93_21# _05_ 1.12e-20
C1149 _34_/a_47_47# _48_/a_27_47# 4.45e-21
C1150 _52_/a_584_47# _06_ 0.00218f
C1151 _21_ _10_ 0.00421f
C1152 net1 _29_/a_29_53# 9.76e-19
C1153 _02_ _07_ 0.0083f
C1154 input3/a_27_47# b[1] 1.31e-20
C1155 b[3] net3 0.0026f
C1156 _00_ net4 0.0166f
C1157 _50_/a_27_47# net16 2.35e-20
C1158 p[3] _06_ 1.59e-20
C1159 _37_/a_27_47# _43_/a_193_413# 0.0102f
C1160 _13_ _00_ 3.77e-20
C1161 net11 net6 1.08e-19
C1162 _14_ _42_/a_109_93# 0.00141f
C1163 net6 p[8] 5.98e-19
C1164 _04_ _10_ 9.24e-20
C1165 _27_/a_205_297# _03_ 1.46e-20
C1166 _32_/a_27_47# _20_ 0.0069f
C1167 _45_/a_27_47# _24_ 4.57e-19
C1168 _33_/a_209_311# _07_ 0.00859f
C1169 _02_ _48_/a_181_47# 3.9e-19
C1170 _33_/a_368_53# _06_ 1.7e-19
C1171 _45_/a_27_47# _22_ 0.0131f
C1172 _52_/a_93_21# net5 0.0124f
C1173 net6 _06_ 0.308f
C1174 output18/a_27_47# net16 3.45e-19
C1175 input1/a_75_212# b[1] 4.16e-19
C1176 net2 _27_/a_27_297# 0.0131f
C1177 net19 _27_/a_27_297# 1.98e-19
C1178 _26_/a_111_297# net6 1.12e-19
C1179 _10_ _02_ 0.0537f
C1180 _10_ _52_/a_256_47# 1.65e-19
C1181 _15_ net3 0.224f
C1182 net19 _17_ 0.0269f
C1183 net2 _17_ 0.181f
C1184 _03_ _30_/a_215_297# 0.0393f
C1185 b[3] input15/a_27_47# 1.77e-19
C1186 _38_/a_303_47# net4 5.95e-19
C1187 _19_ net3 0.0129f
C1188 _25_ VPWR 0.0829f
C1189 net9 net2 3.64e-20
C1190 net13 _30_/a_297_297# 3.27e-20
C1191 _47_/a_81_21# _32_/a_27_47# 5.06e-21
C1192 net12 _23_ 2.28e-21
C1193 net2 input2/a_27_47# 0.024f
C1194 input2/a_27_47# net19 2.9e-23
C1195 _32_/a_27_47# _18_ 1.18e-20
C1196 input6/a_27_47# _14_ 3.75e-21
C1197 _50_/a_515_93# _10_ 0.00129f
C1198 VPWR _00_ 0.416f
C1199 _15_ input15/a_27_47# 2.15e-20
C1200 net6 net3 0.00152f
C1201 input12/a_27_47# VPWR 0.0646f
C1202 input9/a_75_212# net11 1.1e-20
C1203 net1 _32_/a_303_47# 1.45e-19
C1204 _33_/a_296_53# _05_ 4.53e-19
C1205 VPWR input10/a_27_47# 0.00986f
C1206 net17 _30_/a_109_53# 4.18e-20
C1207 _15_ net7 8.4e-20
C1208 _52_/a_346_47# net5 7.03e-19
C1209 _40_/a_191_297# net15 8.41e-19
C1210 net1 output17/a_27_47# 8.12e-19
C1211 _13_ _05_ 2.57e-20
C1212 net6 _45_/a_205_47# 2.59e-20
C1213 net7 _19_ 0.0458f
C1214 VPWR _26_/a_183_297# -3.03e-19
C1215 _13_ _45_/a_465_47# 0.00134f
C1216 _21_ net14 7.17e-21
C1217 net11 _20_ 0.00128f
C1218 _20_ _35_/a_226_47# 5.19e-20
C1219 net4 net5 0.0447f
C1220 input5/a_664_47# _18_ 1.09e-20
C1221 _10_ _32_/a_27_47# 0.00217f
C1222 _38_/a_303_47# VPWR -4.83e-19
C1223 net6 input15/a_27_47# 0.146f
C1224 _20_ _06_ 0.133f
C1225 _39_/a_47_47# _02_ 0.0127f
C1226 p[10] p[0] 8.21e-20
C1227 input8/a_27_47# VPWR 0.0863f
C1228 _30_/a_215_297# _30_/a_297_297# -8.88e-34
C1229 _13_ net5 0.0352f
C1230 input5/a_381_47# net15 7.15e-19
C1231 _25_ input10/a_27_47# 2.03e-20
C1232 net11 net18 0.00221f
C1233 _45_/a_109_297# net16 5.1e-20
C1234 _04_ net14 0.0863f
C1235 _04_ _49_/a_315_47# 7.71e-19
C1236 _01_ net8 0.0802f
C1237 net18 _06_ 0.0211f
C1238 net14 _02_ 0.00952f
C1239 input12/a_27_47# input10/a_27_47# 0.0154f
C1240 VPWR _05_ 0.127f
C1241 _49_/a_208_47# net8 1.4e-19
C1242 _49_/a_315_47# _02_ 0.00134f
C1243 _03_ _31_/a_285_297# 0.00677f
C1244 _35_/a_226_297# _03_ 0.00101f
C1245 _21_ _34_/a_377_297# 2.37e-19
C1246 _34_/a_285_47# VPWR -0.00233f
C1247 VPWR _45_/a_465_47# -5.05e-19
C1248 _47_/a_81_21# _06_ 0.0388f
C1249 _26_/a_183_297# _00_ 4.53e-19
C1250 _11_ _37_/a_27_47# 0.0018f
C1251 net11 _07_ 0.0206f
C1252 input3/a_27_47# net2 0.0222f
C1253 input3/a_27_47# net19 0.00105f
C1254 VPWR p[14] 0.0416f
C1255 _11_ _40_/a_109_297# 0.00522f
C1256 _18_ _06_ 0.54f
C1257 _20_ net3 4.07e-19
C1258 _35_/a_226_47# _07_ 8.96e-19
C1259 p[7] _09_ 9.25e-21
C1260 _50_/a_515_93# net14 1.39e-20
C1261 _04_ _34_/a_377_297# 1.7e-20
C1262 _06_ _07_ 0.185f
C1263 VPWR net5 0.612f
C1264 _04_ _27_/a_27_297# 0.0526f
C1265 net9 _21_ 0.0282f
C1266 _22_ _49_/a_201_297# 2.45e-20
C1267 _52_/a_93_21# net6 2.33e-19
C1268 _32_/a_197_47# net8 3.39e-20
C1269 _44_/a_256_47# _14_ 0.00124f
C1270 _04_ _17_ 4.34e-19
C1271 input7/a_27_47# net14 3.48e-19
C1272 _27_/a_27_297# _02_ 0.00179f
C1273 _48_/a_27_47# _07_ 0.0524f
C1274 _35_/a_556_47# _08_ 7.71e-19
C1275 _48_/a_181_47# _06_ 6.4e-19
C1276 _35_/a_489_413# _09_ 0.0296f
C1277 _02_ _32_/a_109_47# 3.98e-19
C1278 _42_/a_109_93# net17 3.1e-21
C1279 net11 _10_ 0.0109f
C1280 net9 _04_ 0.0213f
C1281 _53_/a_29_53# output18/a_27_47# 9.46e-19
C1282 output17/a_27_47# p[13] 0.00118f
C1283 _12_ _03_ 2.76e-20
C1284 _10_ _35_/a_226_47# 1.25e-19
C1285 _47_/a_81_21# net3 6.66e-19
C1286 net2 _47_/a_299_297# 1.18e-19
C1287 _17_ _02_ 0.00482f
C1288 input2/a_27_47# _04_ 4.5e-21
C1289 _00_ _05_ 5.03e-22
C1290 _22_ _16_ 3.8e-19
C1291 net7 _20_ 0.0257f
C1292 _10_ _06_ 1.14f
C1293 p[7] net10 4.96e-19
C1294 net3 _18_ 7.34e-20
C1295 _25_ net5 6.42e-19
C1296 _10_ _26_/a_111_297# 7.13e-20
C1297 net9 _02_ 0.00611f
C1298 _03_ _09_ 0.326f
C1299 _22_ net15 2.74e-19
C1300 _15_ net4 0.00427f
C1301 _55_/a_217_297# _43_/a_27_47# 2.18e-19
C1302 _15_ _13_ 3.69e-20
C1303 _50_/a_615_93# _15_ 0.00183f
C1304 _10_ _48_/a_27_47# 4.55e-19
C1305 net1 _31_/a_35_297# 0.0111f
C1306 _37_/a_109_47# net19 1.16e-20
C1307 _04_ _26_/a_29_53# 2.3e-21
C1308 _00_ net5 0.00954f
C1309 net13 _30_/a_215_297# 0.0246f
C1310 net9 _33_/a_209_311# 4.33e-20
C1311 _43_/a_297_47# _06_ 4.81e-20
C1312 p[10] net17 0.18f
C1313 input7/a_27_47# _27_/a_27_297# 0.00119f
C1314 _03_ _30_/a_392_297# 6.33e-19
C1315 _26_/a_29_53# _02_ 0.0466f
C1316 _18_ input15/a_27_47# 8.27e-21
C1317 p[11] p[8] 0.0023f
C1318 net7 _18_ 2.58e-20
C1319 input14/a_27_47# _44_/a_250_297# 8.25e-21
C1320 input8/a_27_47# _05_ 1.58e-19
C1321 _37_/a_27_47# _42_/a_109_93# 2.55e-20
C1322 _10_ net3 3.89e-19
C1323 b[3] VPWR 0.367f
C1324 p[2] p[1] 0.178f
C1325 p[6] p[4] 0.0051f
C1326 p[1] net15 6.22e-20
C1327 net10 _03_ 0.32f
C1328 net4 net6 0.713f
C1329 input5/a_558_47# _01_ 3.97e-20
C1330 input5/a_664_47# net14 0.0179f
C1331 _50_/a_615_93# net6 1.43e-19
C1332 _37_/a_27_47# input5/a_841_47# 4.64e-20
C1333 _13_ net6 0.0106f
C1334 _10_ _45_/a_205_47# 6.19e-20
C1335 input7/a_27_47# input2/a_27_47# 1.62e-19
C1336 VPWR _34_/a_47_47# 0.0372f
C1337 output19/a_27_47# p[8] 0.0218f
C1338 _50_/a_343_93# _12_ 5.63e-20
C1339 _50_/a_343_93# _14_ 9.76e-19
C1340 net12 _22_ 5.73e-20
C1341 _50_/a_27_47# _22_ 0.0276f
C1342 net18 _52_/a_93_21# 8.21e-21
C1343 _53_/a_111_297# _09_ 3.4e-19
C1344 output19/a_27_47# _06_ 1.53e-19
C1345 _15_ VPWR 0.912f
C1346 _39_/a_47_47# _06_ 1.44e-19
C1347 net12 p[6] 0.0255f
C1348 _34_/a_285_47# _05_ 7.85e-21
C1349 _55_/a_217_297# _14_ 0.0116f
C1350 net9 _32_/a_27_47# 0.0136f
C1351 net11 net14 9.95e-19
C1352 VPWR _52_/a_584_47# -9.47e-19
C1353 _10_ input15/a_27_47# 4.5e-19
C1354 VPWR _19_ 0.0335f
C1355 net7 _10_ 6.22e-20
C1356 net14 p[8] 0.00868f
C1357 p[3] VPWR 0.0874f
C1358 _01_ _35_/a_76_199# 3.08e-21
C1359 input6/a_27_47# _37_/a_27_47# 9.35e-19
C1360 input3/a_27_47# _04_ 3.55e-19
C1361 p[11] net3 0.00406f
C1362 net14 _06_ 1.94e-19
C1363 net2 p[9] 0.00112f
C1364 b[3] _00_ 1.04e-19
C1365 _52_/a_93_21# _18_ 1.97e-19
C1366 net19 p[9] 0.0729f
C1367 p[12] _12_ 2.08e-20
C1368 _22_ output18/a_27_47# 7.51e-19
C1369 _33_/a_368_53# VPWR -4.26e-19
C1370 input5/a_664_47# _27_/a_27_297# 0.0116f
C1371 net12 _36_/a_197_47# 4.67e-20
C1372 _25_ _34_/a_47_47# 1.08e-19
C1373 _22_ _49_/a_75_199# 9.85e-21
C1374 VPWR net6 0.999f
C1375 input5/a_381_47# output17/a_27_47# 6.6e-20
C1376 _49_/a_201_297# net8 7.3e-19
C1377 net1 _30_/a_109_53# 0.0297f
C1378 b[0] net16 0.0306f
C1379 output19/a_27_47# net3 0.00348f
C1380 _39_/a_47_47# net3 1.66e-20
C1381 net10 _30_/a_297_297# 1.68e-19
C1382 _55_/a_80_21# net1 1.8e-19
C1383 input13/a_27_47# _33_/a_209_311# 5.85e-20
C1384 net13 _35_/a_226_297# 6.88e-19
C1385 _22_ _29_/a_29_53# 2.24e-21
C1386 net13 _31_/a_285_297# 3.85e-20
C1387 net9 input5/a_664_47# 5.29e-19
C1388 input12/a_27_47# _34_/a_47_47# 2.17e-19
C1389 _04_ _49_/a_544_297# 0.00204f
C1390 _44_/a_250_297# p[13] 4.09e-20
C1391 net19 _41_/a_59_75# 3.1e-20
C1392 _15_ _00_ 0.207f
C1393 input5/a_664_47# input2/a_27_47# 4.47e-21
C1394 _45_/a_27_47# _35_/a_76_199# 2.04e-21
C1395 _20_ net4 3.01e-20
C1396 output18/a_27_47# output16/a_27_47# 7.85e-19
C1397 net11 _27_/a_27_297# 1.58e-20
C1398 _13_ _20_ 7.38e-21
C1399 _16_ net8 0.00624f
C1400 _34_/a_377_297# _06_ 0.00427f
C1401 _50_/a_615_93# _20_ 8.8e-19
C1402 _10_ _52_/a_93_21# 0.00534f
C1403 net3 net14 0.689f
C1404 net2 _01_ 2.72e-19
C1405 net19 _01_ 4.9e-19
C1406 net17 _31_/a_117_297# 0.00149f
C1407 input14/a_27_47# _11_ 1.42e-19
C1408 p[2] net8 0.00956f
C1409 net15 net8 0.2f
C1410 net9 net11 0.136f
C1411 _17_ _06_ 0.0341f
C1412 _15_ _26_/a_183_297# 4.63e-36
C1413 net9 _35_/a_226_47# 1.22e-20
C1414 _50_/a_223_47# net16 4.77e-21
C1415 _00_ net6 0.00178f
C1416 input9/a_75_212# VPWR 0.0641f
C1417 _03_ net17 5.1e-19
C1418 net9 _06_ 0.0505f
C1419 p[7] p[5] 6.77e-20
C1420 net13 _12_ 0.00632f
C1421 net4 _18_ 0.023f
C1422 _27_/a_277_297# _03_ 2.1e-20
C1423 _14_ _42_/a_209_311# 0.00142f
C1424 _11_ net16 0.172f
C1425 net11 input11/a_27_47# 0.00318f
C1426 net7 net14 2.23e-19
C1427 _13_ _18_ 0.019f
C1428 net13 _36_/a_27_47# 0.0488f
C1429 net11 _26_/a_29_53# 1.08e-20
C1430 _45_/a_109_297# _22_ 0.0425f
C1431 input7/a_27_47# input1/a_75_212# 3.2e-20
C1432 net13 _09_ 0.0379f
C1433 _38_/a_27_47# _12_ 0.0527f
C1434 b[3] p[14] 0.0645f
C1435 input8/a_27_47# p[3] 0.0023f
C1436 net7 _49_/a_315_47# 0.00706f
C1437 _34_/a_47_47# _05_ 1.26e-20
C1438 _13_ _07_ 3.22e-23
C1439 net3 _27_/a_27_297# 0.0166f
C1440 VPWR _20_ 0.342f
C1441 _08_ _23_ 1.81e-19
C1442 _26_/a_29_53# _06_ 0.0135f
C1443 _38_/a_27_47# _09_ 0.00195f
C1444 _17_ net3 0.0698f
C1445 net18 VPWR 0.104f
C1446 net9 net3 5.09e-20
C1447 _39_/a_285_47# net16 1.29e-19
C1448 _39_/a_47_47# _52_/a_93_21# 1.44e-20
C1449 net13 _30_/a_392_297# 6.64e-20
C1450 net12 net8 0.00458f
C1451 _15_ p[14] 5.32e-19
C1452 p[3] _05_ 5.83e-21
C1453 _10_ net4 0.183f
C1454 _50_/a_615_93# _10_ 8.82e-19
C1455 net13 net10 0.375f
C1456 net1 input5/a_841_47# 1.33e-19
C1457 _13_ _10_ 0.0621f
C1458 _47_/a_81_21# VPWR 0.00889f
C1459 _15_ net5 0.0352f
C1460 _11_ _23_ 2e-20
C1461 net7 _27_/a_27_297# 1.22e-19
C1462 _33_/a_368_53# _05_ 9.2e-19
C1463 _17_ input15/a_27_47# 6.14e-19
C1464 VPWR _18_ 0.0721f
C1465 _36_/a_27_47# _30_/a_215_297# 7.13e-20
C1466 _29_/a_183_297# _04_ 0.0015f
C1467 _52_/a_584_47# net5 0.0022f
C1468 _40_/a_297_297# net15 4.08e-19
C1469 _19_ net5 6.41e-21
C1470 net12 _33_/a_109_93# 0.0435f
C1471 _26_/a_29_53# net3 2.83e-21
C1472 net6 _45_/a_465_47# 6.06e-20
C1473 VPWR _07_ 0.0728f
C1474 input5/a_558_47# _44_/a_93_21# 2.71e-19
C1475 _20_ _00_ 0.271f
C1476 _25_ net18 0.0594f
C1477 _49_/a_75_199# net8 0.00214f
C1478 net9 net7 0.00233f
C1479 p[14] net6 0.00237f
C1480 input13/a_27_47# _35_/a_226_47# 3.94e-20
C1481 _21_ _01_ 7.94e-19
C1482 input3/a_27_47# p[8] 6.2e-19
C1483 input5/a_62_47# p[0] 1.39e-19
C1484 net7 input2/a_27_47# 0.00213f
C1485 net6 net5 0.722f
C1486 input13/a_27_47# _06_ 7.75e-19
C1487 VPWR _48_/a_181_47# -3.35e-19
C1488 input8/a_27_47# input9/a_75_212# 3.09e-20
C1489 p[10] net1 1.22e-19
C1490 _39_/a_285_47# _23_ 1.9e-20
C1491 net18 input10/a_27_47# 4.16e-20
C1492 input5/a_558_47# net15 0.00672f
C1493 _04_ _01_ 0.119f
C1494 VPWR _10_ 0.577f
C1495 net10 _30_/a_215_297# 0.0512f
C1496 _47_/a_81_21# _00_ 0.0258f
C1497 _39_/a_47_47# net4 0.0202f
C1498 _01_ _02_ 0.106f
C1499 _00_ _18_ 0.157f
C1500 input9/a_75_212# _05_ 1.24e-21
C1501 _21_ _45_/a_27_47# 1.18e-20
C1502 _39_/a_47_47# _13_ 0.00117f
C1503 _03_ _31_/a_285_47# 8.54e-19
C1504 b[3] _15_ 0.00162f
C1505 _22_ _43_/a_193_413# 0.00133f
C1506 _47_/a_299_297# _06_ 0.0174f
C1507 _02_ _49_/a_208_47# 0.00193f
C1508 _11_ _40_/a_191_297# 0.00207f
C1509 input3/a_27_47# net3 0.03f
C1510 VPWR _43_/a_297_47# -2.11e-19
C1511 net4 net14 2.21e-21
C1512 _25_ _10_ 0.0109f
C1513 _50_/a_615_93# net14 1.69e-20
C1514 _20_ _05_ 6.79e-19
C1515 p[11] VPWR 0.247f
C1516 _43_/a_27_47# _12_ 2.33e-21
C1517 _14_ _43_/a_27_47# 0.00938f
C1518 _53_/a_29_53# _11_ 2.33e-20
C1519 input5/a_841_47# p[13] 1.73e-19
C1520 _44_/a_346_47# _14_ 3.76e-19
C1521 _35_/a_226_297# _12_ 3.35e-20
C1522 _45_/a_27_47# _02_ 0.00449f
C1523 _44_/a_93_21# net19 0.0074f
C1524 net2 _44_/a_93_21# 0.0273f
C1525 _10_ _00_ 0.301f
C1526 _32_/a_303_47# net8 2.22e-34
C1527 b[3] net6 7.68e-19
C1528 _48_/a_109_47# _07_ 3.01e-19
C1529 _02_ _32_/a_197_47# 3.78e-19
C1530 _42_/a_209_311# net17 1.04e-21
C1531 net13 net17 5.21e-20
C1532 _35_/a_226_297# _09_ 4.98e-19
C1533 _15_ _19_ 1.46e-20
C1534 _20_ net5 0.0651f
C1535 output17/a_27_47# net8 0.0043f
C1536 _47_/a_299_297# net3 2.55e-19
C1537 VPWR output19/a_27_47# 0.0229f
C1538 _39_/a_47_47# VPWR 0.0668f
C1539 p[7] net1 7.5e-20
C1540 net19 _16_ 0.206f
C1541 net2 _16_ 0.00654f
C1542 _32_/a_27_47# _01_ 0.0266f
C1543 _10_ _26_/a_183_297# 5.74e-19
C1544 _43_/a_297_47# _00_ 1.26e-19
C1545 net2 net15 0.324f
C1546 net19 net15 0.0501f
C1547 _15_ net6 0.17f
C1548 _17_ net4 7.52e-21
C1549 p[10] p[13] 0.124f
C1550 _07_ _05_ 1.21e-19
C1551 net12 _35_/a_76_199# 0.0132f
C1552 _37_/a_109_47# net3 0.00212f
C1553 _38_/a_303_47# _10_ 7.36e-19
C1554 VPWR net14 0.182f
C1555 net7 input1/a_75_212# 3.77e-19
C1556 _35_/a_226_297# net10 2.48e-19
C1557 _34_/a_285_47# _07_ 0.00975f
C1558 _47_/a_81_21# net5 4.59e-19
C1559 net7 _49_/a_544_297# 2.72e-19
C1560 VPWR _49_/a_315_47# 6.26e-19
C1561 net10 _31_/a_285_297# 1.68e-19
C1562 net9 net4 1.99e-22
C1563 _12_ _36_/a_27_47# 0.00178f
C1564 _03_ _30_/a_465_297# 7.72e-19
C1565 _43_/a_369_47# _06_ -2.02e-19
C1566 _18_ net5 0.0426f
C1567 _14_ _12_ 1.98e-20
C1568 net13 p[5] 1.05e-19
C1569 _12_ _09_ 0.00509f
C1570 p[9] p[8] 0.0518f
C1571 net11 _29_/a_183_297# 3.64e-19
C1572 net1 _03_ 0.298f
C1573 _37_/a_27_47# _42_/a_209_311# 1.59e-20
C1574 p[6] _08_ 1.55e-19
C1575 net17 _30_/a_215_297# 4.69e-20
C1576 _39_/a_47_47# _00_ 1.85e-20
C1577 input4/a_75_212# _06_ 0.00205f
C1578 p[9] _06_ 0.00205f
C1579 b[0] output16/a_27_47# 0.014f
C1580 _10_ _05_ 9.25e-21
C1581 b[1] output17/a_27_47# 0.00945f
C1582 _26_/a_29_53# net4 0.00412f
C1583 _10_ _45_/a_465_47# 3.32e-19
C1584 VPWR _34_/a_377_297# -0.00192f
C1585 b[3] _20_ 1.37e-19
C1586 VPWR _27_/a_27_297# 0.0329f
C1587 VPWR _32_/a_109_47# 0.00124f
C1588 _53_/a_183_297# _09_ 4.18e-19
C1589 p[14] _10_ 1.53e-19
C1590 _22_ _30_/a_109_53# 3.67e-21
C1591 _35_/a_76_199# _29_/a_29_53# 9.88e-19
C1592 _00_ net14 4.11e-20
C1593 _50_/a_223_47# _22_ 0.031f
C1594 _39_/a_377_297# _06_ 8.76e-20
C1595 VPWR _17_ 0.306f
C1596 _10_ net5 0.199f
C1597 _55_/a_472_297# _14_ 0.00192f
C1598 _55_/a_80_21# _22_ 0.00926f
C1599 net10 _12_ 7.82e-20
C1600 _11_ _24_ 7.29e-20
C1601 net11 _01_ 3.82e-20
C1602 net10 _36_/a_27_47# 0.0366f
C1603 _11_ _22_ 0.15f
C1604 _41_/a_59_75# _06_ 0.0429f
C1605 p[3] input9/a_75_212# 0.0157f
C1606 input5/a_381_47# _42_/a_109_93# 0.00763f
C1607 _43_/a_193_413# net8 1.62e-20
C1608 net10 _09_ 0.037f
C1609 net9 VPWR 0.5f
C1610 _54_/a_75_212# output18/a_27_47# 2.28e-19
C1611 input2/a_27_47# VPWR 0.00872f
C1612 _15_ _20_ 0.691f
C1613 _01_ _06_ 0.00157f
C1614 net3 p[9] 1.63e-19
C1615 _29_/a_183_297# net3 7.38e-21
C1616 net12 _36_/a_303_47# 1.37e-19
C1617 _04_ _49_/a_201_297# 0.0253f
C1618 _19_ _20_ 0.00734f
C1619 p[11] p[14] 3.13e-20
C1620 _44_/a_93_21# _04_ 4.47e-21
C1621 net1 _30_/a_297_297# 7.34e-20
C1622 VPWR input11/a_27_47# 0.0375f
C1623 net10 _30_/a_392_297# 3.4e-19
C1624 VPWR _26_/a_29_53# 0.0356f
C1625 net8 _31_/a_35_297# 0.0408f
C1626 net11 _45_/a_27_47# 3.64e-20
C1627 _45_/a_27_47# _35_/a_226_47# 5.71e-21
C1628 net11 _34_/a_129_47# 0.00242f
C1629 input15/a_27_47# p[9] 0.0196f
C1630 input4/a_75_212# input15/a_27_47# 1.1e-21
C1631 _17_ _00_ 0.0851f
C1632 _20_ net6 9.69e-20
C1633 _15_ _47_/a_81_21# 0.00332f
C1634 net2 _27_/a_109_297# 7.24e-20
C1635 _15_ _18_ 0.042f
C1636 _45_/a_27_47# _06_ 0.0021f
C1637 output19/a_27_47# p[14] 0.0932f
C1638 p[2] _04_ 1.83e-20
C1639 net3 _01_ 1.16e-19
C1640 _34_/a_47_47# _07_ 0.011f
C1641 _34_/a_129_47# _06_ 5.3e-19
C1642 _04_ net15 0.0569f
C1643 _16_ _02_ 0.00564f
C1644 net9 _00_ 0.00501f
C1645 _39_/a_47_47# net5 0.0352f
C1646 _03_ _23_ 0.0564f
C1647 b[3] _10_ 3.27e-20
C1648 p[2] _02_ 7.08e-19
C1649 output18/a_27_47# b[2] 0.0141f
C1650 net15 _02_ 0.0806f
C1651 p[14] net14 6.11e-20
C1652 _41_/a_59_75# input15/a_27_47# 3.96e-20
C1653 _47_/a_81_21# net6 2.14e-19
C1654 _47_/a_299_297# net4 3.28e-19
C1655 net14 net5 0.0263f
C1656 _26_/a_29_53# _00_ 0.0466f
C1657 net6 _18_ 0.166f
C1658 net13 _36_/a_109_47# 0.00126f
C1659 _22_ _42_/a_109_93# 1.21e-19
C1660 input10/a_27_47# input11/a_27_47# 5.3e-19
C1661 net7 _01_ 0.233f
C1662 _15_ _10_ 0.479f
C1663 input13/a_27_47# VPWR 0.0696f
C1664 net12 _21_ 0.23f
C1665 _50_/a_27_47# _21_ 3.38e-21
C1666 b[1] _31_/a_35_297# 3.21e-19
C1667 input3/a_27_47# VPWR 0.0687f
C1668 _38_/a_109_47# _12_ 0.00179f
C1669 input8/a_27_47# net9 3.71e-20
C1670 net7 _49_/a_208_47# 0.00312f
C1671 net2 output17/a_27_47# 0.0285f
C1672 p[11] b[3] 0.243f
C1673 p[3] _10_ 1.37e-20
C1674 p[2] input7/a_27_47# 0.0023f
C1675 _14_ net17 2.4e-20
C1676 _50_/a_27_47# _04_ 2.07e-21
C1677 input7/a_27_47# net15 1.88e-19
C1678 net12 _04_ 0.267f
C1679 _21_ output18/a_27_47# 0.00103f
C1680 net8 _30_/a_109_53# 1.76e-20
C1681 net13 _30_/a_465_297# 6.36e-20
C1682 _10_ net6 0.0965f
C1683 input1/a_75_212# VPWR 0.0786f
C1684 _55_/a_80_21# net8 1.84e-21
C1685 net13 net1 3.51e-19
C1686 net9 _05_ 0.124f
C1687 net12 _02_ 2.28e-19
C1688 _50_/a_27_47# _02_ 2.09e-19
C1689 p[14] _17_ 5.46e-21
C1690 _27_/a_27_297# net5 3.48e-19
C1691 _21_ _49_/a_75_199# 6.64e-19
C1692 VPWR _49_/a_544_297# 0.00569f
C1693 input2/a_27_47# _05_ 1.83e-19
C1694 _32_/a_109_47# net5 5.69e-21
C1695 b[3] output19/a_27_47# 0.00809f
C1696 _11_ net8 1.81e-20
C1697 p[11] _15_ 2.93e-19
C1698 _47_/a_299_297# VPWR 0.0643f
C1699 _17_ net5 0.00408f
C1700 _21_ _29_/a_29_53# 0.0775f
C1701 net12 _33_/a_209_311# 0.0769f
C1702 _04_ _49_/a_75_199# 0.0782f
C1703 input5/a_664_47# _44_/a_93_21# 1.88e-20
C1704 net9 net5 0.0368f
C1705 output18/a_27_47# _02_ 3.6e-19
C1706 b[3] net14 0.0172f
C1707 net10 net17 8.67e-21
C1708 _43_/a_297_47# net6 8.23e-22
C1709 _37_/a_109_47# VPWR -4.38e-19
C1710 _47_/a_81_21# _20_ 0.0457f
C1711 _20_ _18_ 0.0151f
C1712 _49_/a_75_199# _02_ 0.0354f
C1713 _04_ _29_/a_29_53# 0.0408f
C1714 input5/a_62_47# net1 7.59e-20
C1715 _37_/a_27_47# _14_ 0.00137f
C1716 p[1] p[10] 9.52e-20
C1717 _04_ _27_/a_109_297# 7.2e-20
C1718 _40_/a_109_297# _14_ -1.78e-33
C1719 input4/a_75_212# net4 0.0189f
C1720 net11 _49_/a_201_297# 1.42e-19
C1721 _20_ _07_ 1.28e-21
C1722 _02_ _29_/a_29_53# 6.76e-21
C1723 _49_/a_201_297# _35_/a_226_47# 1.66e-20
C1724 _26_/a_29_53# net5 0.0237f
C1725 input5/a_664_47# net15 0.0216f
C1726 _15_ net14 0.225f
C1727 input9/a_75_212# _10_ 5.49e-21
C1728 _45_/a_27_47# _52_/a_93_21# 1.18e-19
C1729 net1 _30_/a_215_297# 0.00375f
C1730 _47_/a_299_297# _00_ 7.59e-21
C1731 _38_/a_27_47# net16 0.114f
C1732 output19/a_27_47# net6 0.00112f
C1733 _39_/a_47_47# net6 0.0249f
C1734 _39_/a_377_297# net4 8.88e-19
C1735 _19_ net14 0.0512f
C1736 net12 _32_/a_27_47# 1.52e-19
C1737 _47_/a_81_21# _18_ 7.96e-20
C1738 p[5] net10 0.00544f
C1739 net19 _43_/a_193_413# 3.31e-19
C1740 _10_ _20_ 0.179f
C1741 net2 _43_/a_193_413# 1.52e-19
C1742 _41_/a_59_75# net4 1.76e-19
C1743 _19_ _49_/a_315_47# 1.33e-19
C1744 _16_ _06_ 0.00162f
C1745 b[3] _17_ 0.00637f
C1746 net6 net14 2.82e-21
C1747 VPWR _43_/a_369_47# -3.75e-19
C1748 net15 p[8] 3.39e-19
C1749 _11_ _40_/a_297_297# 9.94e-19
C1750 p[7] p[6] 0.217f
C1751 input13/a_27_47# _05_ 3.93e-19
C1752 net15 _06_ 0.033f
C1753 _15_ _27_/a_27_297# 9.85e-20
C1754 VPWR p[9] 0.374f
C1755 input4/a_75_212# VPWR 0.06f
C1756 input5/a_841_47# net8 0.025f
C1757 net13 _23_ 4.11e-19
C1758 _29_/a_183_297# VPWR -8.13e-19
C1759 net2 _44_/a_250_297# 0.0169f
C1760 _45_/a_109_297# _02_ 8.44e-19
C1761 _44_/a_93_21# net3 0.0102f
C1762 _44_/a_250_297# net19 0.00592f
C1763 _15_ _17_ 0.0752f
C1764 net2 _31_/a_35_297# 0.0635f
C1765 _04_ output17/a_27_47# 0.027f
C1766 _47_/a_81_21# _10_ 0.0061f
C1767 net11 p[4] 0.0557f
C1768 _19_ _27_/a_27_297# 0.082f
C1769 net9 _34_/a_47_47# 1.41e-20
C1770 _48_/a_181_47# _07_ 5.93e-19
C1771 _35_/a_556_47# _09_ 3.74e-19
C1772 _02_ _32_/a_303_47# 1.15e-20
C1773 _35_/a_76_199# _08_ 0.0061f
C1774 _10_ _18_ 0.133f
C1775 _16_ net3 1.77e-19
C1776 _17_ _19_ 8.82e-21
C1777 _15_ net9 0.00113f
C1778 _15_ input2/a_27_47# 3.18e-20
C1779 _24_ _03_ 9.46e-20
C1780 _45_/a_27_47# net4 0.024f
C1781 _22_ _03_ 2.55e-20
C1782 _10_ _07_ 2.19e-19
C1783 _13_ _45_/a_27_47# 0.0703f
C1784 VPWR _41_/a_59_75# 0.0179f
C1785 net7 _49_/a_201_297# 0.00419f
C1786 net15 net3 0.394f
C1787 input2/a_27_47# _19_ 5.26e-20
C1788 p[3] net9 0.0376f
C1789 net12 net11 0.358f
C1790 input5/a_62_47# p[13] 0.0202f
C1791 net11 _50_/a_27_47# 6.05e-21
C1792 p[10] net8 0.0097f
C1793 _39_/a_47_47# _20_ 2.3e-20
C1794 VPWR _01_ 0.521f
C1795 _17_ net6 3.12e-19
C1796 net12 _35_/a_226_47# 8.29e-19
C1797 _15_ _26_/a_29_53# 0.00192f
C1798 net1 _31_/a_285_297# 5.85e-19
C1799 net12 _06_ 0.284f
C1800 _47_/a_299_297# net5 0.00198f
C1801 _50_/a_27_47# _06_ 0.00972f
C1802 _11_ _35_/a_76_199# 6.99e-22
C1803 _26_/a_29_53# _52_/a_584_47# 7.45e-20
C1804 _16_ input15/a_27_47# 7.13e-19
C1805 VPWR _49_/a_208_47# -5.93e-19
C1806 net7 _16_ 7.5e-20
C1807 net11 output18/a_27_47# 6.84e-20
C1808 _20_ net14 8.01e-20
C1809 net12 _48_/a_27_47# 0.0126f
C1810 p[2] net7 0.00156f
C1811 net15 input15/a_27_47# 0.00325f
C1812 net7 net15 2.91e-19
C1813 net11 _49_/a_75_199# 4.49e-19
C1814 output18/a_27_47# _06_ 0.0114f
C1815 _49_/a_75_199# _35_/a_226_47# 8.73e-20
C1816 _39_/a_47_47# _18_ 1.23e-19
C1817 _26_/a_29_53# net6 0.0032f
C1818 _45_/a_27_47# VPWR -0.00418f
C1819 _53_/a_111_297# _24_ 9.08e-21
C1820 _41_/a_59_75# _00_ 2.43e-20
C1821 VPWR _34_/a_129_47# -9.47e-19
C1822 _53_/a_111_297# _22_ 4.7e-20
C1823 net11 _29_/a_29_53# 0.00514f
C1824 input3/a_27_47# b[3] 0.012f
C1825 _10_ _43_/a_297_47# 0.00118f
C1826 _35_/a_226_47# _29_/a_29_53# 2.64e-19
C1827 VPWR _32_/a_197_47# 0.00146f
C1828 _00_ _01_ 0.00124f
C1829 _50_/a_343_93# _22_ 0.0597f
C1830 p[10] b[1] 0.286f
C1831 _29_/a_29_53# _06_ 0.00111f
C1832 _55_/a_80_21# net19 0.00423f
C1833 net1 _36_/a_27_47# 6.99e-20
C1834 _11_ _54_/a_75_212# 3.22e-20
C1835 b[0] b[2] 0.183f
C1836 _04_ _43_/a_193_413# 5.67e-21
C1837 net1 _09_ 5.26e-20
C1838 input5/a_381_47# _42_/a_209_311# 3.88e-19
C1839 input5/a_558_47# _42_/a_109_93# 1.75e-19
C1840 net14 _18_ 0.0147f
C1841 _53_/a_29_53# _38_/a_27_47# 1.29e-19
C1842 _11_ net19 2.19e-19
C1843 _11_ net2 0.234f
C1844 net9 input9/a_75_212# 0.0247f
C1845 _55_/a_300_47# _14_ 8.09e-19
C1846 _20_ _27_/a_27_297# 3.14e-20
C1847 input3/a_27_47# _15_ 7.53e-19
C1848 _43_/a_193_413# _02_ 9.4e-21
C1849 input5/a_558_47# input5/a_841_47# -4.44e-34
C1850 _11_ _45_/a_193_297# 0.0292f
C1851 _17_ _20_ 0.102f
C1852 output19/a_27_47# _10_ 3.23e-20
C1853 p[12] _22_ 2.13e-21
C1854 _39_/a_47_47# _10_ 0.00824f
C1855 input13/a_27_47# p[3] 0.00101f
C1856 _49_/a_75_199# net3 2.01e-19
C1857 _44_/a_250_297# _04_ 5.57e-21
C1858 net12 net7 1.57e-19
C1859 net9 _20_ 0.328f
C1860 _04_ _31_/a_35_297# 1.89e-20
C1861 _45_/a_27_47# _00_ 4.84e-20
C1862 p[14] p[9] 0.4f
C1863 p[0] net1 0.00473f
C1864 net10 _30_/a_465_297# 0.00106f
C1865 net3 _29_/a_29_53# 1.68e-20
C1866 input8/a_27_47# _01_ 1.43e-19
C1867 p[7] _33_/a_109_93# 1.15e-19
C1868 net16 _12_ 0.131f
C1869 net8 _31_/a_117_297# 5.91e-19
C1870 net1 net10 0.00388f
C1871 net11 _45_/a_109_297# 7.46e-20
C1872 _10_ net14 2.4e-19
C1873 input4/a_75_212# net5 0.0104f
C1874 _02_ _31_/a_35_297# 0.00316f
C1875 _45_/a_109_297# _35_/a_226_47# 1.59e-21
C1876 _27_/a_109_297# net3 5.45e-19
C1877 _15_ _47_/a_299_297# 0.0103f
C1878 net16 _09_ 0.00707f
C1879 _47_/a_81_21# _17_ 0.0456f
C1880 input5/a_558_47# p[10] 1.09e-19
C1881 _45_/a_109_297# _06_ 0.0023f
C1882 _34_/a_377_297# _07_ 5.8e-19
C1883 _26_/a_29_53# _20_ 0.00447f
C1884 _17_ _18_ 0.271f
C1885 _03_ net8 0.0287f
C1886 net7 _49_/a_75_199# 0.09f
C1887 _01_ _05_ 5.03e-19
C1888 net17 _31_/a_285_47# 0.00134f
C1889 p[14] _41_/a_59_75# 5.13e-20
C1890 _39_/a_377_297# net5 0.00234f
C1891 net9 _47_/a_81_21# 3.49e-19
C1892 net9 _18_ 1.51e-19
C1893 net18 _26_/a_29_53# 2.57e-21
C1894 _41_/a_59_75# net5 2.41e-19
C1895 _21_ _08_ 0.00139f
C1896 _43_/a_297_47# net14 1.09e-21
C1897 net7 _29_/a_29_53# 6.01e-19
C1898 _33_/a_109_93# _03_ 2.78e-19
C1899 net9 _07_ 1.39e-20
C1900 _16_ net4 2.73e-20
C1901 _47_/a_299_297# net6 3.63e-19
C1902 _01_ net5 0.0779f
C1903 p[11] net14 0.00182f
C1904 net2 _42_/a_109_93# 0.00507f
C1905 _22_ _42_/a_209_311# 1.72e-19
C1906 net19 _42_/a_109_93# 0.0448f
C1907 _04_ _08_ 5.99e-19
C1908 net15 net4 8.68e-19
C1909 net13 _22_ 4.63e-20
C1910 input13/a_27_47# input9/a_75_212# 0.00732f
C1911 _26_/a_29_53# _18_ 5.26e-20
C1912 _12_ _23_ 0.00743f
C1913 b[1] _31_/a_117_297# 2.34e-19
C1914 _45_/a_27_47# _05_ 9.34e-23
C1915 _21_ _30_/a_109_53# 3.31e-20
C1916 _50_/a_223_47# _21_ 2.91e-21
C1917 _36_/a_27_47# _23_ 0.00118f
C1918 _10_ _17_ 0.0233f
C1919 _02_ _08_ 2.26e-20
C1920 _09_ _23_ 0.207f
C1921 _38_/a_27_47# _22_ 2.86e-19
C1922 _32_/a_27_47# _31_/a_35_297# 9.17e-20
C1923 net9 _10_ 0.0438f
C1924 _38_/a_197_47# _12_ 0.00173f
C1925 _11_ _21_ 9.98e-20
C1926 output19/a_27_47# net14 0.00142f
C1927 VPWR _49_/a_201_297# 0.0185f
C1928 net3 output17/a_27_47# 0.00248f
C1929 b[3] p[9] 0.0898f
C1930 _04_ _30_/a_109_53# 9.19e-21
C1931 b[1] _03_ 0.00143f
C1932 _50_/a_223_47# _04_ 7.89e-22
C1933 _44_/a_93_21# VPWR 0.005f
C1934 net8 _30_/a_297_297# 2.42e-21
C1935 net13 _36_/a_197_47# 1.06e-19
C1936 _33_/a_209_311# _08_ 0.0122f
C1937 _50_/a_343_93# net8 7.25e-19
C1938 _45_/a_27_47# net5 0.0288f
C1939 _17_ _43_/a_297_47# 5.72e-20
C1940 _02_ _30_/a_109_53# 5.03e-22
C1941 _32_/a_197_47# net5 5.61e-21
C1942 _50_/a_223_47# _02_ 2.51e-20
C1943 input6/a_27_47# net19 0.00586f
C1944 input6/a_27_47# net2 0.0047f
C1945 p[0] p[13] 1.88e-19
C1946 _38_/a_27_47# output16/a_27_47# 9.02e-19
C1947 _47_/a_384_47# VPWR -1.45e-19
C1948 p[10] net2 0.0632f
C1949 p[10] net19 1.26e-21
C1950 VPWR _16_ 0.126f
C1951 _55_/a_80_21# _02_ 0.164f
C1952 _10_ _26_/a_29_53# 0.0265f
C1953 _15_ p[9] 2.06e-19
C1954 p[11] _17_ 1.93e-19
C1955 _11_ _02_ 0.0621f
C1956 _22_ _30_/a_215_297# 2.46e-21
C1957 net10 _23_ 7.53e-19
C1958 p[2] VPWR 0.103f
C1959 net7 output17/a_27_47# 0.00185f
C1960 net12 _33_/a_296_53# 1.23e-20
C1961 VPWR net15 0.61f
C1962 net1 net17 2.89e-19
C1963 net12 net4 2.57e-20
C1964 _50_/a_27_47# net4 0.0239f
C1965 b[3] _01_ 9.26e-20
C1966 _47_/a_299_297# _20_ 0.002f
C1967 p[12] _52_/a_250_297# 1.84e-20
C1968 _50_/a_27_47# _13_ 0.00169f
C1969 _43_/a_193_413# _06_ 0.0138f
C1970 _43_/a_369_47# net6 3.62e-21
C1971 _39_/a_47_47# _17_ 1.47e-20
C1972 output19/a_27_47# _17_ 0.00122f
C1973 _04_ _29_/a_111_297# 9.25e-19
C1974 _40_/a_191_297# _14_ 2.4e-19
C1975 _15_ _41_/a_59_75# 0.0139f
C1976 _44_/a_93_21# _00_ 4.54e-20
C1977 _39_/a_285_47# _02_ 0.0019f
C1978 input4/a_75_212# net6 0.0273f
C1979 net6 p[9] 0.14f
C1980 VPWR p[4] 0.112f
C1981 net14 _27_/a_27_297# 0.0118f
C1982 _15_ _01_ 0.007f
C1983 _53_/a_29_53# _12_ 3.46e-20
C1984 _16_ _00_ 0.00613f
C1985 _17_ net14 0.104f
C1986 _47_/a_384_47# _00_ 5.15e-20
C1987 _38_/a_109_47# net16 4.17e-19
C1988 _32_/a_27_47# _30_/a_109_53# 1.51e-19
C1989 _53_/a_29_53# _09_ 0.00642f
C1990 _39_/a_377_297# net6 0.00143f
C1991 net9 net14 7.12e-20
C1992 _19_ _01_ 0.031f
C1993 net15 _00_ 0.00147f
C1994 _43_/a_193_413# net3 5.65e-20
C1995 input2/a_27_47# net14 0.0102f
C1996 _21_ input5/a_841_47# 1.59e-21
C1997 _41_/a_59_75# net6 0.0373f
C1998 input8/a_27_47# _49_/a_201_297# 2.46e-21
C1999 _35_/a_76_199# _03_ 0.0733f
C2000 input5/a_381_47# _14_ 5.68e-20
C2001 _11_ _32_/a_27_47# 1.65e-20
C2002 net12 VPWR 0.817f
C2003 _50_/a_27_47# VPWR -0.00335f
C2004 _19_ _49_/a_208_47# 7.12e-20
C2005 VPWR _43_/a_469_47# -2.75e-19
C2006 _04_ _42_/a_109_93# 5.77e-22
C2007 _42_/a_209_311# net8 7.7e-21
C2008 net13 net8 7.51e-20
C2009 _26_/a_29_53# net14 1.33e-20
C2010 _17_ _27_/a_27_297# 6.78e-22
C2011 _44_/a_250_297# net3 0.0088f
C2012 _22_ _43_/a_27_47# 0.091f
C2013 _53_/a_29_53# net10 7.88e-22
C2014 VPWR output18/a_27_47# 0.0689f
C2015 _02_ input5/a_841_47# 0.00591f
C2016 _43_/a_193_413# input15/a_27_47# 1.62e-20
C2017 _47_/a_299_297# _10_ 0.0134f
C2018 input12/a_27_47# p[4] 8.26e-19
C2019 net7 _43_/a_193_413# 3.49e-19
C2020 VPWR _49_/a_75_199# 0.0177f
C2021 input8/a_27_47# p[2] 0.0159f
C2022 input10/a_27_47# p[4] 0.0215f
C2023 net11 _08_ 8.83e-19
C2024 net9 _32_/a_109_47# 6.44e-19
C2025 net12 _25_ 4.46e-20
C2026 net13 _33_/a_109_93# 0.0254f
C2027 _54_/a_75_212# _03_ 5.45e-21
C2028 _35_/a_226_47# _08_ 0.00117f
C2029 input3/a_27_47# p[11] 0.0157f
C2030 input2/a_27_47# _27_/a_27_297# 1.16e-19
C2031 _39_/a_129_47# VPWR -9.47e-19
C2032 VPWR _29_/a_29_53# 0.0299f
C2033 _08_ _06_ 0.0343f
C2034 _45_/a_109_297# net4 6.43e-20
C2035 _44_/a_93_21# p[14] 2.82e-20
C2036 net9 _17_ 2.89e-23
C2037 _45_/a_27_47# net6 0.021f
C2038 net2 _03_ 1.89e-19
C2039 _50_/a_27_47# _00_ 0.00197f
C2040 p[10] _04_ 0.00306f
C2041 VPWR _27_/a_109_297# -2.45e-19
C2042 net12 input12/a_27_47# 0.0295f
C2043 input5/a_62_47# net8 2.05e-19
C2044 _44_/a_93_21# net5 3.61e-20
C2045 p[2] _05_ 3.69e-19
C2046 net12 input10/a_27_47# 0.00115f
C2047 _03_ _45_/a_193_297# 2.57e-20
C2048 _25_ output18/a_27_47# 0.072f
C2049 input3/a_27_47# output19/a_27_47# 4.77e-21
C2050 _08_ _48_/a_27_47# 2.58e-19
C2051 p[10] _02_ 2.17e-19
C2052 net7 _31_/a_35_297# 0.0384f
C2053 _43_/a_369_47# _18_ 1.49e-19
C2054 _30_/a_215_297# net8 8.14e-21
C2055 _06_ _30_/a_109_53# 1.96e-19
C2056 _16_ net5 1.99e-20
C2057 _50_/a_223_47# _06_ 0.0481f
C2058 _47_/a_384_47# net5 0.00129f
C2059 _12_ _24_ 1.67e-19
C2060 _11_ p[8] 7.7e-20
C2061 _20_ _41_/a_59_75# 1.78e-20
C2062 _55_/a_80_21# _06_ 5.15e-19
C2063 p[14] net15 0.00132f
C2064 _22_ _12_ 0.196f
C2065 _14_ _22_ 0.00449f
C2066 _22_ _36_/a_27_47# 2.82e-20
C2067 input4/a_75_212# _18_ 4.36e-19
C2068 _11_ _06_ 0.493f
C2069 input3/a_27_47# net14 3.47e-19
C2070 _20_ _01_ 0.161f
C2071 net9 _26_/a_29_53# 0.00343f
C2072 _24_ _09_ 0.0202f
C2073 net15 net5 0.0226f
C2074 _22_ _09_ 0.0279f
C2075 _39_/a_129_47# _00_ 1.63e-20
C2076 _33_/a_109_93# _30_/a_215_297# 0.00104f
C2077 p[11] _37_/a_109_47# 2.84e-20
C2078 _45_/a_109_297# VPWR -0.011f
C2079 _53_/a_183_297# _22_ 3.71e-20
C2080 _47_/a_81_21# _41_/a_59_75# 1.5e-19
C2081 net11 _29_/a_111_297# 8.27e-19
C2082 _10_ _43_/a_369_47# 0.00199f
C2083 VPWR _32_/a_303_47# 6.03e-19
C2084 _50_/a_343_93# net2 1.25e-20
C2085 _39_/a_285_47# _06_ 1.23e-20
C2086 VPWR output17/a_27_47# 0.0263f
C2087 _29_/a_111_297# _06_ 6.74e-20
C2088 net12 _05_ 0.0414f
C2089 _55_/a_80_21# net3 2.35e-19
C2090 _47_/a_81_21# _01_ 6.05e-21
C2091 _01_ _18_ 6.1e-20
C2092 net7 _08_ 9.54e-25
C2093 _34_/a_285_47# net12 8.07e-20
C2094 _10_ p[9] 0.00225f
C2095 _11_ net3 0.165f
C2096 input4/a_75_212# _10_ 0.00372f
C2097 input8/a_27_47# _49_/a_75_199# 1.99e-20
C2098 input5/a_558_47# _42_/a_209_311# 7.85e-20
C2099 b[3] _44_/a_93_21# 0.00491f
C2100 _29_/a_183_297# _10_ 6.24e-20
C2101 p[7] _04_ 0.00142f
C2102 net10 p[6] 0.0023f
C2103 _35_/a_489_413# _21_ 0.0448f
C2104 b[3] _16_ 2.9e-19
C2105 _50_/a_27_47# net5 0.0169f
C2106 net12 net5 0.0674f
C2107 _37_/a_109_47# net14 1.71e-19
C2108 _39_/a_377_297# _10_ 7.42e-19
C2109 p[12] net19 6.8e-20
C2110 input13/a_27_47# net9 2.42e-19
C2111 input5/a_381_47# net17 1.37e-20
C2112 _15_ _44_/a_93_21# 0.0168f
C2113 _45_/a_109_297# _00_ 4.86e-20
C2114 _10_ _41_/a_59_75# 0.0172f
C2115 p[1] p[0] 0.161f
C2116 net7 _55_/a_80_21# 0.00163f
C2117 _21_ _03_ 0.0818f
C2118 b[3] net15 0.00408f
C2119 _11_ input15/a_27_47# 4.4e-19
C2120 p[7] _33_/a_209_311# 1.34e-19
C2121 net8 _31_/a_285_297# 0.0215f
C2122 _13_ _43_/a_193_413# 5.58e-21
C2123 _45_/a_27_47# _18_ 0.00347f
C2124 p[11] p[9] 0.114f
C2125 net13 _35_/a_76_199# 0.0337f
C2126 _10_ _01_ 2.22e-19
C2127 _42_/a_109_93# _06_ 5.53e-20
C2128 _29_/a_29_53# _05_ 3.79e-20
C2129 _35_/a_489_413# _02_ 3.86e-19
C2130 _15_ _16_ 0.0607f
C2131 _15_ _47_/a_384_47# 0.00112f
C2132 _04_ _03_ 0.586f
C2133 _45_/a_27_47# _07_ 1.02e-20
C2134 input5/a_841_47# _06_ 1.66e-19
C2135 _39_/a_129_47# net5 0.00344f
C2136 _15_ net15 0.156f
C2137 _35_/a_489_413# _33_/a_209_311# 2.77e-20
C2138 _44_/a_93_21# net6 1.08e-20
C2139 _02_ _03_ 0.00474f
C2140 output19/a_27_47# p[9] 0.0852f
C2141 _29_/a_29_53# net5 8.1e-20
C2142 _39_/a_47_47# input4/a_75_212# 3.1e-19
C2143 p[3] p[2] 0.164f
C2144 _37_/a_109_47# _17_ 8.86e-21
C2145 net15 _19_ 0.00628f
C2146 _43_/a_369_47# net14 6.79e-21
C2147 input6/a_27_47# p[8] 0.00139f
C2148 _33_/a_209_311# _03_ 8.38e-19
C2149 _16_ net6 1.62e-20
C2150 _45_/a_27_47# _10_ 0.0143f
C2151 _42_/a_109_93# net3 0.0435f
C2152 input6/a_27_47# _06_ 2.85e-19
C2153 net19 _42_/a_209_311# 0.0766f
C2154 _53_/a_111_297# _21_ 4.38e-19
C2155 _52_/a_250_297# _12_ 0.0139f
C2156 VPWR _43_/a_193_413# 0.0063f
C2157 net14 p[9] 1.05e-19
C2158 net2 _42_/a_209_311# 5.1e-19
C2159 _36_/a_27_47# net8 1.52e-19
C2160 _14_ net8 4.23e-19
C2161 net15 net6 0.0664f
C2162 _37_/a_197_47# net2 4.74e-20
C2163 _54_/a_75_212# _38_/a_27_47# 2.67e-19
C2164 b[1] _31_/a_285_297# 1.12e-19
C2165 _45_/a_109_297# _05_ 2.79e-22
C2166 _52_/a_250_297# _09_ 1.97e-20
C2167 _36_/a_109_47# _23_ 3.44e-19
C2168 b[0] net4 0.0024f
C2169 net12 _34_/a_47_47# 0.0385f
C2170 _33_/a_109_93# _12_ 9.75e-20
C2171 _13_ b[0] 0.00299f
C2172 output17/a_27_47# _05_ 1.12e-19
C2173 _15_ _50_/a_27_47# 5.65e-19
C2174 _33_/a_109_93# _09_ 7.36e-20
C2175 _44_/a_250_297# VPWR 0.0231f
C2176 net13 _36_/a_303_47# 5.5e-20
C2177 _53_/a_111_297# _02_ 9.57e-20
C2178 VPWR _31_/a_35_297# 0.0333f
C2179 _45_/a_109_297# net5 0.0184f
C2180 _32_/a_27_47# _03_ 1.9e-19
C2181 _17_ _43_/a_369_47# 5.87e-19
C2182 input5/a_62_47# net2 0.0197f
C2183 _50_/a_343_93# _02_ 6.94e-19
C2184 input6/a_27_47# net3 2.52e-19
C2185 net14 _01_ 8.29e-19
C2186 _32_/a_303_47# net5 7.18e-21
C2187 net10 net8 2.05e-21
C2188 p[10] net3 7.98e-19
C2189 net1 p[13] 2.13e-19
C2190 _49_/a_201_297# _20_ 5.24e-21
C2191 net7 input5/a_841_47# 0.00193f
C2192 _55_/a_217_297# _02_ 6.01e-19
C2193 net10 _52_/a_250_297# 2.86e-21
C2194 _43_/a_193_413# _00_ 0.00721f
C2195 _49_/a_315_47# _01_ 1.82e-19
C2196 net5 output17/a_27_47# 5.01e-20
C2197 _17_ p[9] 1.03e-20
C2198 input9/a_75_212# p[2] 5.13e-20
C2199 p[1] net17 6.65e-20
C2200 net12 _33_/a_368_53# 2.63e-19
C2201 _50_/a_223_47# net4 0.0107f
C2202 net12 net6 0.00643f
C2203 _50_/a_27_47# net6 0.0428f
C2204 _39_/a_47_47# _45_/a_27_47# 1.31e-19
C2205 input14/a_27_47# p[13] 1.37e-19
C2206 _16_ _20_ 0.00271f
C2207 _55_/a_80_21# net4 1.06e-19
C2208 _50_/a_223_47# _13_ 8.2e-20
C2209 _47_/a_384_47# _20_ 1.72e-19
C2210 _33_/a_109_93# net10 0.0336f
C2211 net9 _29_/a_183_297# 3.51e-19
C2212 _43_/a_469_47# net6 4.85e-21
C2213 VPWR b[0] 0.142f
C2214 p[5] p[6] 0.198f
C2215 _19_ _49_/a_75_199# 0.0206f
C2216 p[7] _35_/a_226_47# 2.82e-19
C2217 _11_ net4 0.0858f
C2218 input6/a_27_47# input15/a_27_47# 5.3e-19
C2219 p[7] _06_ 0.00864f
C2220 _40_/a_297_297# _14_ 1.58e-19
C2221 _44_/a_250_297# _00_ 6.39e-20
C2222 _11_ _13_ 0.164f
C2223 net15 _20_ 0.0021f
C2224 net7 p[10] 0.00481f
C2225 _17_ _41_/a_59_75# 0.00149f
C2226 _01_ _32_/a_109_47# 0.00129f
C2227 _01_ _27_/a_27_297# 8.04e-19
C2228 p[3] _29_/a_29_53# 2.07e-19
C2229 VPWR _08_ -0.0171f
C2230 _44_/a_93_21# _18_ 0.00485f
C2231 _17_ _01_ 1.46e-20
C2232 _27_/a_109_297# _19_ 7.54e-21
C2233 p[0] b[1] 0.00123f
C2234 _39_/a_129_47# net6 6.91e-19
C2235 _39_/a_285_47# net4 9.71e-19
C2236 _35_/a_489_413# _06_ 9.22e-19
C2237 _50_/a_343_93# _32_/a_27_47# 6.48e-20
C2238 net13 _21_ 0.13f
C2239 net6 _29_/a_29_53# 1.4e-20
C2240 _16_ _18_ 0.144f
C2241 net9 _01_ 0.157f
C2242 _38_/a_197_47# net16 5.89e-19
C2243 net11 _03_ 0.0952f
C2244 _39_/a_285_47# _13_ 0.00451f
C2245 VPWR _30_/a_109_53# 0.0012f
C2246 _35_/a_226_47# _03_ 0.028f
C2247 _47_/a_81_21# net15 0.00106f
C2248 _50_/a_223_47# VPWR -0.00601f
C2249 net15 _18_ 0.0382f
C2250 b[3] output17/a_27_47# 4.01e-20
C2251 _04_ _42_/a_209_311# 9.84e-22
C2252 _55_/a_80_21# VPWR 0.0289f
C2253 _38_/a_27_47# _21_ 3.87e-19
C2254 _03_ _06_ 0.00635f
C2255 net13 _04_ 0.569f
C2256 input8/a_27_47# _31_/a_35_297# 0.00955f
C2257 _11_ VPWR 0.352f
C2258 _45_/a_27_47# _17_ 1.16e-20
C2259 _44_/a_93_21# _10_ 2.48e-19
C2260 _42_/a_209_311# _02_ 9.92e-19
C2261 net12 _20_ 0.00437f
C2262 _43_/a_193_413# net5 1.39e-20
C2263 net13 _02_ 0.00154f
C2264 net2 _43_/a_27_47# 0.01f
C2265 net2 _44_/a_346_47# 1.64e-19
C2266 _44_/a_256_47# net3 0.00101f
C2267 _35_/a_76_199# _12_ 6.84e-20
C2268 _44_/a_346_47# net19 0.00124f
C2269 _35_/a_76_199# _36_/a_27_47# 3.22e-19
C2270 _10_ _16_ 0.00486f
C2271 _47_/a_384_47# _10_ 3.53e-19
C2272 _05_ _31_/a_35_297# 0.00649f
C2273 input5/a_381_47# net1 1.27e-19
C2274 net9 _32_/a_197_47# 6.06e-19
C2275 _38_/a_27_47# _02_ 0.00103f
C2276 net17 net8 0.18f
C2277 _04_ _27_/a_205_297# 6.42e-19
C2278 net13 _33_/a_209_311# 0.0227f
C2279 _35_/a_76_199# _09_ 0.0374f
C2280 _39_/a_285_47# VPWR -9.53e-19
C2281 _19_ output17/a_27_47# 7.69e-19
C2282 _21_ _30_/a_215_297# 1.48e-19
C2283 _10_ net15 0.0101f
C2284 input5/a_62_47# _04_ 0.00345f
C2285 _27_/a_277_297# net8 7.99e-20
C2286 input9/a_75_212# _29_/a_29_53# 9.7e-21
C2287 VPWR _29_/a_111_297# -5.85e-19
C2288 net3 _03_ 4.27e-20
C2289 _11_ _25_ 7.05e-19
C2290 _45_/a_109_297# net6 7.82e-19
C2291 _00_ _30_/a_109_53# 3.67e-20
C2292 _50_/a_223_47# _00_ 0.00738f
C2293 _49_/a_75_199# _20_ 0.0233f
C2294 _44_/a_250_297# net5 3.11e-20
C2295 net5 _31_/a_35_297# 2.04e-21
C2296 _55_/a_80_21# _00_ 5.5e-19
C2297 _04_ _30_/a_215_297# 0.00225f
C2298 _50_/a_27_47# _18_ 0.0665f
C2299 _39_/a_129_47# _20_ 1.71e-20
C2300 net12 _18_ 2.25e-21
C2301 net18 output18/a_27_47# 0.0106f
C2302 _53_/a_111_297# _06_ 3.82e-19
C2303 _11_ _00_ 0.238f
C2304 _53_/a_29_53# net16 2.04e-20
C2305 net7 _31_/a_117_297# 0.00472f
C2306 _20_ _29_/a_29_53# 0.0111f
C2307 _43_/a_469_47# _18_ 1.59e-19
C2308 VPWR _28_/a_109_297# -1.71e-19
C2309 net12 _07_ 0.18f
C2310 _50_/a_343_93# _06_ 0.0376f
C2311 _02_ _30_/a_215_297# 3.58e-21
C2312 net10 _35_/a_76_199# 0.0146f
C2313 _55_/a_217_297# _06_ 3.46e-19
C2314 p[11] _16_ 2.17e-20
C2315 net2 _12_ 1.02e-20
C2316 _44_/a_93_21# output19/a_27_47# 7.25e-20
C2317 _14_ net19 0.00714f
C2318 net2 _14_ 0.0104f
C2319 net7 _03_ 0.078f
C2320 p[11] net15 3.83e-19
C2321 _12_ _45_/a_193_297# 0.0103f
C2322 p[12] p[8] 0.0153f
C2323 _08_ _05_ 0.00897f
C2324 _33_/a_209_311# _30_/a_215_297# 1.56e-19
C2325 _39_/a_285_47# _00_ 1.47e-21
C2326 _37_/a_27_47# net8 6.66e-21
C2327 b[0] net5 2.76e-19
C2328 b[1] net17 0.00766f
C2329 _49_/a_201_297# net14 1.52e-19
C2330 VPWR _42_/a_109_93# -0.00118f
C2331 _34_/a_285_47# _08_ 0.00414f
C2332 net12 _10_ 0.00257f
C2333 _09_ _45_/a_193_297# 0.00961f
C2334 _50_/a_27_47# _10_ 0.0154f
C2335 p[12] _06_ 0.0535f
C2336 _49_/a_75_199# _07_ 4.05e-21
C2337 VPWR input5/a_841_47# 0.0775f
C2338 _44_/a_93_21# net14 0.0646f
C2339 _10_ _43_/a_469_47# 0.00124f
C2340 _47_/a_299_297# _41_/a_59_75# 0.00146f
C2341 _39_/a_47_47# net15 9.44e-22
C2342 output19/a_27_47# net15 6.88e-19
C2343 _49_/a_544_297# _01_ 0.00109f
C2344 _30_/a_109_53# _05_ 0.033f
C2345 _29_/a_29_53# _07_ 1.19e-20
C2346 _54_/a_75_212# net10 6.24e-19
C2347 _16_ net14 0.00266f
C2348 _55_/a_217_297# net3 5.78e-20
C2349 _15_ _43_/a_193_413# 4.86e-19
C2350 net1 _22_ 0.0129f
C2351 net1 p[6] 3.12e-20
C2352 net2 net10 2.05e-20
C2353 b[3] _44_/a_250_297# 0.0112f
C2354 input5/a_664_47# _42_/a_209_311# 0.0124f
C2355 _12_ b[2] 3.89e-20
C2356 _55_/a_300_47# _22_ 2.08e-19
C2357 _20_ _32_/a_303_47# 1.54e-19
C2358 net15 net14 1.07f
C2359 input5/a_381_47# p[13] 0.00153f
C2360 _43_/a_193_413# _19_ 4.85e-21
C2361 _52_/a_93_21# _03_ 0.00985f
C2362 input6/a_27_47# VPWR 0.00162f
C2363 _09_ b[2] 4.28e-20
C2364 p[2] _49_/a_315_47# 6.65e-20
C2365 p[10] VPWR 0.177f
C2366 net5 _30_/a_109_53# 5.84e-22
C2367 _50_/a_223_47# net5 0.00202f
C2368 _39_/a_129_47# _10_ 2.51e-19
C2369 _55_/a_80_21# net5 2.78e-19
C2370 _10_ _29_/a_29_53# 5.17e-19
C2371 input5/a_558_47# net17 2.88e-21
C2372 _35_/a_226_297# _04_ 4.51e-19
C2373 _15_ _44_/a_250_297# 0.00517f
C2374 _11_ net5 0.207f
C2375 p[1] net1 0.0291f
C2376 net7 _55_/a_217_297# 1.04e-19
C2377 _44_/a_93_21# _17_ 0.0646f
C2378 _43_/a_193_413# net6 2.41e-20
C2379 _43_/a_27_47# _02_ 1.88e-21
C2380 net13 net11 0.093f
C2381 net8 _31_/a_285_47# 0.00129f
C2382 net13 _35_/a_226_47# 0.00709f
C2383 net16 _24_ 6.93e-19
C2384 _02_ _31_/a_285_297# 5.86e-20
C2385 _16_ _27_/a_27_297# 3.74e-22
C2386 _42_/a_209_311# _06_ 1.66e-19
C2387 _22_ net16 0.00606f
C2388 _19_ _31_/a_35_297# 1.47e-19
C2389 _47_/a_384_47# _17_ 1.1e-20
C2390 net13 _06_ 0.0766f
C2391 net11 _38_/a_27_47# 1.68e-20
C2392 _16_ _17_ 0.242f
C2393 p[12] input15/a_27_47# 5.48e-19
C2394 net15 _27_/a_27_297# 0.00888f
C2395 _38_/a_27_47# _06_ 0.0172f
C2396 _21_ _12_ 7.99e-20
C2397 _17_ net15 0.195f
C2398 _39_/a_285_47# net5 0.0405f
C2399 _21_ _36_/a_27_47# 0.0276f
C2400 net9 p[2] 1.4e-20
C2401 _21_ _09_ 0.263f
C2402 output16/a_27_47# net16 0.0101f
C2403 net9 net15 8.49e-20
C2404 _43_/a_469_47# net14 1.44e-20
C2405 input5/a_62_47# p[8] 1.15e-19
C2406 _41_/a_59_75# p[9] 1.02e-19
C2407 input4/a_75_212# _41_/a_59_75# 0.00153f
C2408 _04_ _12_ 1.42e-19
C2409 input2/a_27_47# net15 1.61e-19
C2410 _04_ _36_/a_27_47# 0.00169f
C2411 _08_ _34_/a_47_47# 0.00123f
C2412 _04_ _14_ 2.04e-21
C2413 _45_/a_109_297# _10_ 0.00202f
C2414 _42_/a_209_311# net3 0.029f
C2415 net13 net3 3.25e-21
C2416 net11 _30_/a_215_297# 1.04e-19
C2417 _04_ _09_ 0.0904f
C2418 net19 _42_/a_296_53# 2.71e-19
C2419 _13_ _03_ 1.74e-20
C2420 _37_/a_197_47# net3 0.0028f
C2421 _24_ _23_ 0.012f
C2422 _12_ _02_ 0.265f
C2423 p[7] VPWR 0.0184f
C2424 _37_/a_303_47# net2 4.41e-19
C2425 b[3] _55_/a_80_21# 3.55e-19
C2426 _02_ _36_/a_27_47# 9.37e-20
C2427 _14_ _02_ 0.0316f
C2428 b[3] _11_ 2.37e-20
C2429 _49_/a_75_199# net14 3.67e-19
C2430 _30_/a_215_297# _06_ 2.03e-20
C2431 _26_/a_29_53# net15 9.06e-21
C2432 _22_ _23_ 0.0186f
C2433 b[0] net6 2.52e-19
C2434 _43_/a_27_47# _32_/a_27_47# 2.01e-20
C2435 _02_ _09_ 0.297f
C2436 net12 _34_/a_377_297# 0.00251f
C2437 _21_ net10 0.0254f
C2438 _43_/a_193_413# _20_ 0.00161f
C2439 _49_/a_315_47# _49_/a_75_199# 1.78e-33
C2440 net2 net17 0.261f
C2441 _33_/a_209_311# _12_ 2.88e-20
C2442 net19 net17 8.84e-23
C2443 net14 _29_/a_29_53# 1.61e-20
C2444 net2 _44_/a_584_47# 0.0053f
C2445 _42_/a_109_93# net5 0.00109f
C2446 _15_ _50_/a_223_47# 0.00698f
C2447 _50_/a_27_47# _17_ 3.93e-20
C2448 _44_/a_256_47# VPWR -7.56e-19
C2449 _27_/a_109_297# net14 1.32e-19
C2450 _27_/a_205_297# net3 4.37e-19
C2451 VPWR _31_/a_117_297# 8.41e-19
C2452 _35_/a_489_413# VPWR -0.00725f
C2453 _33_/a_209_311# _09_ 3.79e-20
C2454 _33_/a_368_53# _08_ 5.04e-19
C2455 _15_ _55_/a_80_21# 0.107f
C2456 _53_/a_183_297# _02_ 4.14e-19
C2457 net5 input5/a_841_47# 0.0221f
C2458 input4/a_75_212# _45_/a_27_47# 2.18e-20
C2459 _04_ net10 0.121f
C2460 net13 net7 1.72e-19
C2461 _17_ _43_/a_469_47# 0.00177f
C2462 input5/a_62_47# net3 0.00164f
C2463 net1 net8 0.381f
C2464 _11_ _15_ 0.113f
C2465 input11/a_27_47# p[4] 0.0646f
C2466 p[3] _30_/a_109_53# 3.23e-20
C2467 net12 net9 0.0596f
C2468 _55_/a_472_297# _02_ 1.25e-19
C2469 p[10] _05_ 6e-20
C2470 net10 _52_/a_256_47# 8.13e-20
C2471 VPWR _03_ 0.845f
C2472 net10 _02_ 3.52e-19
C2473 _20_ _31_/a_35_297# 1.69e-19
C2474 _53_/a_111_297# net4 2.09e-19
C2475 _49_/a_75_199# _27_/a_27_297# 0.011f
C2476 _01_ _49_/a_208_47# 2.13e-19
C2477 _43_/a_193_413# _18_ 0.0413f
C2478 _50_/a_343_93# net4 0.00124f
C2479 _50_/a_223_47# net6 0.0194f
C2480 input6/a_27_47# p[14] 0.0155f
C2481 p[7] input12/a_27_47# 3.2e-20
C2482 _33_/a_209_311# net10 0.0419f
C2483 _55_/a_217_297# net4 1.13e-19
C2484 _50_/a_343_93# _13_ 5.63e-20
C2485 b[3] _28_/a_109_297# 7.49e-20
C2486 net12 _26_/a_29_53# 6.55e-19
C2487 _50_/a_27_47# _26_/a_29_53# 5.56e-19
C2488 _32_/a_27_47# _36_/a_27_47# 0.011f
C2489 _11_ net6 0.0257f
C2490 p[10] net5 5.12e-21
C2491 net7 input5/a_62_47# 2.04e-19
C2492 _39_/a_129_47# _17_ 1.38e-20
C2493 _27_/a_109_297# _27_/a_27_297# -3.68e-20
C2494 net9 _49_/a_75_199# 0.00382f
C2495 input3/a_27_47# net15 6.19e-20
C2496 net2 _40_/a_109_297# 0.0011f
C2497 _37_/a_27_47# net2 0.0692f
C2498 _37_/a_27_47# net19 0.0105f
C2499 net13 _52_/a_93_21# 7.21e-19
C2500 _01_ _32_/a_197_47# 0.00156f
C2501 _25_ _03_ 0.00422f
C2502 p[12] net4 0.00758f
C2503 input7/a_27_47# p[0] 5.13e-20
C2504 net9 _29_/a_29_53# 0.0205f
C2505 _53_/a_29_53# _24_ 0.0835f
C2506 b[3] _42_/a_109_93# 3.29e-19
C2507 _15_ _28_/a_109_297# 0.00346f
C2508 _43_/a_27_47# _06_ 0.0329f
C2509 net1 b[1] 1.78e-20
C2510 _10_ _43_/a_193_413# 0.0174f
C2511 _53_/a_29_53# _22_ 0.00749f
C2512 _06_ _31_/a_285_297# 1.01e-20
C2513 _35_/a_226_297# _06_ 1.28e-19
C2514 _00_ _03_ 2.31e-20
C2515 _39_/a_285_47# net6 1.53e-19
C2516 VPWR _41_/a_145_75# -2.46e-19
C2517 input13/a_27_47# p[4] 7.37e-20
C2518 _53_/a_111_297# VPWR 1.11e-34
C2519 _47_/a_299_297# net15 1.44e-20
C2520 net10 _32_/a_27_47# 2.76e-20
C2521 VPWR _30_/a_297_297# -4.57e-19
C2522 _26_/a_29_53# _29_/a_29_53# 0.00121f
C2523 _50_/a_343_93# VPWR -0.0126f
C2524 _15_ _42_/a_109_93# 0.00367f
C2525 _55_/a_217_297# VPWR -0.00133f
C2526 net12 input13/a_27_47# 0.0163f
C2527 _45_/a_109_297# _17_ 4.29e-22
C2528 _42_/a_109_93# _19_ 1.14e-21
C2529 _50_/a_223_47# _20_ 1.71e-19
C2530 _20_ _30_/a_109_53# 8.12e-19
C2531 input6/a_27_47# b[3] 4.02e-19
C2532 p[13] net8 0.00345f
C2533 net11 _12_ 0.00799f
C2534 b[3] p[10] 3.13e-20
C2535 _44_/a_346_47# net3 8.04e-19
C2536 _35_/a_226_47# _12_ 8.38e-20
C2537 net11 _36_/a_27_47# 0.0717f
C2538 _55_/a_80_21# _20_ 0.0291f
C2539 _52_/a_250_297# _23_ 3.17e-19
C2540 p[12] VPWR 0.0378f
C2541 _04_ net17 0.0218f
C2542 _11_ _20_ 0.268f
C2543 net11 _09_ 0.0262f
C2544 _38_/a_109_47# _02_ 1.63e-19
C2545 _12_ _06_ 0.136f
C2546 _35_/a_226_47# _09_ 0.058f
C2547 input5/a_558_47# net1 1.1e-19
C2548 net9 _32_/a_303_47# 0.00218f
C2549 _36_/a_27_47# _06_ 0.0501f
C2550 _14_ _06_ 0.0556f
C2551 _04_ _27_/a_277_297# 0.00113f
C2552 net13 _33_/a_296_53# 3.71e-20
C2553 net13 net4 2.48e-19
C2554 _02_ net17 0.0608f
C2555 _08_ _07_ 0.348f
C2556 _09_ _06_ 0.0965f
C2557 input6/a_27_47# _15_ 5.75e-19
C2558 _50_/a_343_93# _00_ 0.102f
C2559 input2/a_27_47# output17/a_27_47# 0.107f
C2560 _03_ _05_ 0.135f
C2561 net13 _13_ 4e-21
C2562 _38_/a_27_47# net4 0.0119f
C2563 p[11] _44_/a_250_297# 1.13e-19
C2564 net7 _43_/a_27_47# 6.31e-19
C2565 _50_/a_223_47# _18_ 0.0367f
C2566 _33_/a_209_311# net17 7.03e-21
C2567 _09_ _48_/a_27_47# 0.00541f
C2568 _38_/a_27_47# _13_ 4.58e-19
C2569 _53_/a_183_297# _06_ 0.00146f
C2570 p[10] _19_ 0.00226f
C2571 net7 _31_/a_285_297# 0.00227f
C2572 _55_/a_80_21# _18_ 1.44e-20
C2573 _11_ _47_/a_81_21# 0.0454f
C2574 net11 net10 0.592f
C2575 _50_/a_429_93# _06_ 0.00169f
C2576 _43_/a_193_413# net14 1.11e-19
C2577 _11_ _18_ 0.484f
C2578 net10 _35_/a_226_47# 0.0159f
C2579 _03_ net5 1.04e-19
C2580 _10_ _08_ 1.51e-19
C2581 _22_ _24_ 0.0846f
C2582 net3 _12_ 3.09e-20
C2583 b[1] p[13] 0.00115f
C2584 net10 _06_ 0.184f
C2585 _14_ net3 0.0295f
C2586 _44_/a_250_297# output19/a_27_47# 6.42e-20
C2587 input6/a_27_47# net6 0.00208f
C2588 _12_ _45_/a_205_47# 7.46e-19
C2589 input7/a_27_47# net17 4.99e-20
C2590 _20_ _28_/a_109_297# 0.00221f
C2591 net15 p[9] 0.00306f
C2592 _49_/a_201_297# _01_ 0.0105f
C2593 VPWR _42_/a_209_311# -0.00753f
C2594 net13 VPWR 0.599f
C2595 net10 _48_/a_27_47# 8.4e-21
C2596 _44_/a_250_297# net14 4.24e-20
C2597 _50_/a_223_47# _10_ 0.0295f
C2598 _37_/a_197_47# VPWR -3.27e-19
C2599 _55_/a_80_21# _10_ 5.49e-19
C2600 _38_/a_27_47# VPWR -0.0142f
C2601 _11_ _10_ 0.176f
C2602 _14_ input15/a_27_47# 9.48e-21
C2603 net2 net1 1.64e-19
C2604 net7 _14_ 0.00251f
C2605 _16_ _01_ 3.24e-19
C2606 _39_/a_47_47# b[0] 2.04e-19
C2607 net15 _41_/a_59_75# 1.16e-20
C2608 net7 _09_ 0.00258f
C2609 _17_ _43_/a_193_413# 0.0503f
C2610 VPWR _27_/a_205_297# 1.05e-19
C2611 p[2] _01_ 0.00164f
C2612 input5/a_381_47# net8 7.48e-19
C2613 net15 _01_ 0.0314f
C2614 _35_/a_556_47# _21_ 2.69e-19
C2615 input5/a_558_47# p[13] 0.00158f
C2616 input5/a_62_47# VPWR 0.0601f
C2617 net13 _25_ 0.00297f
C2618 input3/a_27_47# output17/a_27_47# 3.15e-19
C2619 input14/a_27_47# net2 0.0176f
C2620 input14/a_27_47# net19 1.44e-19
C2621 _50_/a_343_93# net5 0.00124f
C2622 _39_/a_285_47# _10_ 0.00289f
C2623 p[7] p[3] 0.169f
C2624 _55_/a_217_297# net5 8.84e-20
C2625 _25_ _38_/a_27_47# 5.76e-19
C2626 VPWR _30_/a_215_297# -0.00472f
C2627 net7 p[0] 1.36e-19
C2628 _54_/a_75_212# net16 1.69e-21
C2629 p[11] _11_ 4.18e-20
C2630 _44_/a_250_297# _17_ 0.0336f
C2631 p[12] p[14] 0.00425f
C2632 _03_ _34_/a_47_47# 4.5e-20
C2633 _52_/a_93_21# _12_ 0.0157f
C2634 input1/a_75_212# output17/a_27_47# 0.0101f
C2635 _15_ _03_ 7.39e-20
C2636 _10_ _28_/a_109_297# 4.34e-19
C2637 p[12] net5 4.79e-20
C2638 _50_/a_27_47# _41_/a_59_75# 9.59e-22
C2639 _52_/a_93_21# _09_ 0.0227f
C2640 net16 _45_/a_193_297# 0.00187f
C2641 input2/a_27_47# _31_/a_35_297# 0.00136f
C2642 _11_ _39_/a_47_47# 3.9e-19
C2643 net11 net17 3.19e-20
C2644 _19_ _03_ 0.0019f
C2645 net12 _01_ 1.67e-21
C2646 p[3] _03_ 0.00348f
C2647 _50_/a_223_47# net14 5.89e-21
C2648 _13_ _43_/a_27_47# 1.66e-20
C2649 _55_/a_80_21# net14 4.7e-19
C2650 _11_ net14 5e-19
C2651 _04_ _36_/a_109_47# 2.39e-19
C2652 net6 _03_ 2.9e-20
C2653 net19 _42_/a_368_53# 5.12e-19
C2654 _42_/a_296_53# net3 1.81e-19
C2655 _52_/a_93_21# net10 7.84e-20
C2656 _52_/a_346_47# _12_ 3.8e-19
C2657 _22_ net8 3.3e-20
C2658 _52_/a_250_297# _24_ 3.03e-19
C2659 p[7] input9/a_75_212# 0.00102f
C2660 net13 _05_ 0.192f
C2661 net2 p[13] 0.0247f
C2662 b[3] _55_/a_217_297# 3.41e-19
C2663 _37_/a_303_47# net3 0.00133f
C2664 _22_ _52_/a_250_297# 0.099f
C2665 _49_/a_75_199# _01_ 0.009f
C2666 net13 _34_/a_285_47# 4.11e-20
C2667 p[5] net11 0.0598f
C2668 net1 _21_ 0.0252f
C2669 _50_/a_27_47# _45_/a_27_47# 0.109f
C2670 net9 _08_ 7.71e-21
C2671 _45_/a_193_297# _23_ 4.13e-19
C2672 p[14] _42_/a_209_311# 3.45e-22
C2673 net3 net17 3.72e-19
C2674 net4 _12_ 0.105f
C2675 _01_ _29_/a_29_53# 8.33e-20
C2676 _33_/a_109_93# _22_ 1.34e-22
C2677 _42_/a_209_311# net5 3.27e-21
C2678 net4 _36_/a_27_47# 0.0103f
C2679 _15_ _50_/a_343_93# 0.0098f
C2680 _37_/a_27_47# p[8] 9.82e-21
C2681 input6/a_27_47# _10_ 4.57e-20
C2682 VPWR _43_/a_27_47# 0.0186f
C2683 p[11] _42_/a_109_93# 4.55e-21
C2684 _44_/a_346_47# VPWR -8.74e-19
C2685 _50_/a_223_47# _17_ 5.24e-20
C2686 _14_ net4 1.54e-20
C2687 b[3] p[12] 7.54e-20
C2688 net13 net5 0.127f
C2689 _13_ _12_ 0.462f
C2690 _27_/a_277_297# net3 2.71e-19
C2691 VPWR _31_/a_285_297# 0.0174f
C2692 _35_/a_226_297# VPWR -8.54e-19
C2693 net1 _04_ 0.018f
C2694 _15_ _55_/a_217_297# 0.0474f
C2695 net4 _09_ 0.00262f
C2696 _37_/a_27_47# _06_ 2.5e-20
C2697 _13_ _14_ 1.47e-20
C2698 _55_/a_80_21# _17_ 7.64e-21
C2699 _40_/a_109_297# _06_ 0.00175f
C2700 _03_ VGND 0.481f
C2701 net10 VGND 0.909f
C2702 _30_/a_465_297# VGND 0.00105f
C2703 _30_/a_392_297# VGND 7.67e-19
C2704 _30_/a_297_297# VGND -4.43e-19
C2705 _30_/a_109_53# VGND 0.152f
C2706 _30_/a_215_297# VGND 0.158f
C2707 _05_ VGND 0.906f
C2708 net8 VGND 0.791f
C2709 _31_/a_285_297# VGND 1.12e-20
C2710 _31_/a_117_297# VGND -0.00177f
C2711 _31_/a_35_297# VGND 0.246f
C2712 _32_/a_303_47# VGND -4.83e-19
C2713 _32_/a_197_47# VGND 8.12e-20
C2714 _32_/a_109_47# VGND 1.05e-19
C2715 _32_/a_27_47# VGND 0.198f
C2716 _50_/a_615_93# VGND -5.19e-19
C2717 _50_/a_515_93# VGND -4.75e-19
C2718 _50_/a_429_93# VGND 4.71e-19
C2719 _50_/a_343_93# VGND 0.171f
C2720 _50_/a_223_47# VGND 0.157f
C2721 _50_/a_27_47# VGND 0.255f
C2722 _07_ VGND 0.483f
C2723 _06_ VGND 1.91f
C2724 net13 VGND 0.524f
C2725 _33_/a_368_53# VGND 2.38e-19
C2726 _33_/a_296_53# VGND -1.43e-19
C2727 _33_/a_209_311# VGND 0.136f
C2728 _33_/a_109_93# VGND 0.145f
C2729 net12 VGND 0.874f
C2730 _34_/a_285_47# VGND 0.0144f
C2731 _34_/a_129_47# VGND -8.76e-20
C2732 _34_/a_377_297# VGND -9.51e-19
C2733 _34_/a_47_47# VGND 0.289f
C2734 _23_ VGND 0.266f
C2735 p[9] VGND 0.51f
C2736 input15/a_27_47# VGND 0.223f
C2737 _09_ VGND 0.544f
C2738 _08_ VGND 0.293f
C2739 _35_/a_556_47# VGND 1.95e-19
C2740 _35_/a_226_297# VGND -4.55e-19
C2741 _35_/a_489_413# VGND 0.0246f
C2742 _35_/a_226_47# VGND 0.151f
C2743 _35_/a_76_199# VGND 0.137f
C2744 _24_ VGND 0.127f
C2745 _12_ VGND 1.2f
C2746 _52_/a_584_47# VGND -0.00112f
C2747 _52_/a_346_47# VGND -0.00175f
C2748 _52_/a_256_47# VGND -0.00161f
C2749 _52_/a_250_297# VGND 0.0246f
C2750 _52_/a_93_21# VGND 0.133f
C2751 _10_ VGND 1.75f
C2752 _36_/a_303_47# VGND 8.14e-19
C2753 _36_/a_197_47# VGND -3.75e-19
C2754 _36_/a_109_47# VGND 3.56e-19
C2755 _36_/a_27_47# VGND 0.196f
C2756 p[8] VGND 1.25f
C2757 input14/a_27_47# VGND 0.247f
C2758 _53_/a_183_297# VGND -4.34e-19
C2759 _53_/a_111_297# VGND -2.89e-19
C2760 _53_/a_29_53# VGND 0.163f
C2761 _11_ VGND 0.358f
C2762 _37_/a_303_47# VGND -1.63e-19
C2763 _37_/a_197_47# VGND -4.58e-19
C2764 _37_/a_109_47# VGND -7.9e-19
C2765 _37_/a_27_47# VGND 0.16f
C2766 p[7] VGND 0.887f
C2767 input13/a_27_47# VGND 0.255f
C2768 net18 VGND 0.463f
C2769 _25_ VGND 0.39f
C2770 _54_/a_75_212# VGND 0.263f
C2771 _38_/a_303_47# VGND 1.78e-19
C2772 _38_/a_197_47# VGND 2.29e-19
C2773 _38_/a_109_47# VGND 2.3e-19
C2774 _38_/a_27_47# VGND 0.183f
C2775 net19 VGND 0.31f
C2776 _22_ VGND 0.256f
C2777 _14_ VGND 0.454f
C2778 _15_ VGND 0.487f
C2779 _55_/a_300_47# VGND -0.00109f
C2780 _55_/a_472_297# VGND -0.00188f
C2781 _55_/a_217_297# VGND -0.00225f
C2782 _55_/a_80_21# VGND 0.213f
C2783 p[6] VGND 0.742f
C2784 input12/a_27_47# VGND 0.248f
C2785 net9 VGND 0.685f
C2786 p[3] VGND 0.853f
C2787 input9/a_75_212# VGND 0.276f
C2788 _39_/a_285_47# VGND 0.0128f
C2789 _39_/a_129_47# VGND -0.00126f
C2790 _39_/a_377_297# VGND -6.28e-19
C2791 _39_/a_47_47# VGND 0.266f
C2792 net11 VGND 1.25f
C2793 p[5] VGND 0.76f
C2794 input11/a_27_47# VGND 0.235f
C2795 p[2] VGND 0.997f
C2796 input8/a_27_47# VGND 0.265f
C2797 p[4] VGND 1.25f
C2798 input10/a_27_47# VGND 0.211f
C2799 net7 VGND 0.881f
C2800 p[1] VGND 0.914f
C2801 input7/a_27_47# VGND 0.265f
C2802 p[14] VGND 0.985f
C2803 input6/a_27_47# VGND 0.205f
C2804 net5 VGND 2.04f
C2805 p[13] VGND 0.557f
C2806 input5/a_841_47# VGND 0.187f
C2807 input5/a_664_47# VGND 0.144f
C2808 input5/a_558_47# VGND 0.163f
C2809 input5/a_381_47# VGND 0.107f
C2810 input5/a_62_47# VGND 0.218f
C2811 p[12] VGND 1.93f
C2812 input4/a_75_212# VGND 0.263f
C2813 p[11] VGND 0.865f
C2814 input3/a_27_47# VGND 0.249f
C2815 net2 VGND 1.5f
C2816 p[10] VGND 0.79f
C2817 input2/a_27_47# VGND 0.194f
C2818 net1 VGND 0.855f
C2819 p[0] VGND 1.04f
C2820 input1/a_75_212# VGND 0.268f
C2821 b[3] VGND 0.546f
C2822 output19/a_27_47# VGND 0.534f
C2823 b[2] VGND 0.593f
C2824 output18/a_27_47# VGND 0.601f
C2825 _40_/a_297_297# VGND -5.1e-19
C2826 _40_/a_191_297# VGND -9.29e-19
C2827 _40_/a_109_297# VGND -0.00181f
C2828 b[1] VGND 0.526f
C2829 net17 VGND 0.385f
C2830 output17/a_27_47# VGND 0.545f
C2831 _41_/a_145_75# VGND 3.75e-19
C2832 _41_/a_59_75# VGND 0.191f
C2833 b[0] VGND 0.708f
C2834 output16/a_27_47# VGND 0.616f
C2835 _16_ VGND 0.119f
C2836 _42_/a_368_53# VGND -4.05e-19
C2837 _42_/a_209_311# VGND 0.135f
C2838 _42_/a_109_93# VGND 0.153f
C2839 _17_ VGND 0.563f
C2840 _00_ VGND 0.516f
C2841 _43_/a_369_47# VGND -8.43e-19
C2842 _43_/a_297_47# VGND -1.33e-19
C2843 _43_/a_193_413# VGND 0.122f
C2844 _43_/a_27_47# VGND 0.209f
C2845 net6 VGND 1f
C2846 net4 VGND 0.888f
C2847 _26_/a_183_297# VGND 2.42e-19
C2848 _26_/a_111_297# VGND -2.75e-19
C2849 _26_/a_29_53# VGND 0.218f
C2850 _01_ VGND 0.244f
C2851 net14 VGND 0.958f
C2852 net3 VGND 0.786f
C2853 net15 VGND 0.673f
C2854 _27_/a_277_297# VGND -4.65e-19
C2855 _27_/a_205_297# VGND -3.36e-19
C2856 _27_/a_109_297# VGND -6.15e-19
C2857 _27_/a_27_297# VGND 0.147f
C2858 _18_ VGND 0.159f
C2859 _44_/a_584_47# VGND -0.00145f
C2860 _44_/a_346_47# VGND -0.00198f
C2861 _44_/a_256_47# VGND -0.00184f
C2862 _44_/a_250_297# VGND 0.0219f
C2863 _44_/a_93_21# VGND 0.128f
C2864 net16 VGND 0.375f
C2865 _13_ VGND 0.496f
C2866 _45_/a_465_47# VGND -8.14e-19
C2867 _45_/a_205_47# VGND -2.47e-19
C2868 _45_/a_193_297# VGND -0.00131f
C2869 _45_/a_109_297# VGND -0.00108f
C2870 _45_/a_27_47# VGND 0.187f
C2871 _28_/a_109_297# VGND -9.87e-19
C2872 _29_/a_183_297# VGND 4.41e-19
C2873 _29_/a_111_297# VGND -1.9e-19
C2874 _29_/a_29_53# VGND 0.234f
C2875 _19_ VGND 0.497f
C2876 _04_ VGND 0.478f
C2877 _47_/a_384_47# VGND -2.05e-19
C2878 _47_/a_299_297# VGND 0.0344f
C2879 _47_/a_81_21# VGND 0.136f
C2880 VPWR VGND 40.2f
C2881 _48_/a_181_47# VGND 3.03e-19
C2882 _48_/a_109_47# VGND 9.44e-19
C2883 _48_/a_27_47# VGND 0.232f
C2884 _21_ VGND 0.586f
C2885 _20_ VGND 0.709f
C2886 _02_ VGND 2.08f
C2887 _49_/a_315_47# VGND -0.0034f
C2888 _49_/a_208_47# VGND -0.00164f
C2889 _49_/a_544_297# VGND -0.00256f
C2890 _49_/a_201_297# VGND -5.82e-19
C2891 _49_/a_75_199# VGND 0.205f
.ends

.subckt sky130_fd_pr__pfet_01v8_MYW2PY a_n73_n48# a_n33_n145# a_15_n48# w_n211_n267#
+ VSUBS
X0 a_15_n48# a_n33_n145# a_n73_n48# w_n211_n267# sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.54 as=0.139 ps=1.54 w=0.48 l=0.15
C0 a_n73_n48# a_n33_n145# 0.0197f
C1 w_n211_n267# a_n33_n145# 0.237f
C2 a_n33_n145# a_15_n48# 0.0197f
C3 a_n73_n48# w_n211_n267# 0.05f
C4 a_n73_n48# a_15_n48# 0.0795f
C5 w_n211_n267# a_15_n48# 0.05f
C6 a_15_n48# VSUBS 0.0287f
C7 a_n73_n48# VSUBS 0.0287f
C8 a_n33_n145# VSUBS 0.115f
C9 w_n211_n267# VSUBS 1.05f
.ends

.subckt sky130_fd_pr__nfet_01v8_JRGCPP a_n1108_n42# a_1050_n42# a_n1210_n216# a_n1050_n130#
X0 a_1050_n42# a_n1050_n130# a_n1108_n42# a_n1210_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=10.5
C0 a_n1050_n130# a_n1108_n42# 0.0251f
C1 a_1050_n42# a_n1050_n130# 0.0251f
C2 a_1050_n42# a_n1210_n216# 0.0931f
C3 a_n1108_n42# a_n1210_n216# 0.0931f
C4 a_n1050_n130# a_n1210_n216# 5.94f
.ends

.subckt sky130_fd_pr__pfet_01v8_XJ78MR a_n73_n1050# w_n211_n1269# a_15_n1050# a_n33_n1147#
+ VSUBS
X0 a_15_n1050# a_n33_n1147# a_n73_n1050# w_n211_n1269# sky130_fd_pr__pfet_01v8 ad=3.05 pd=21.6 as=3.05 ps=21.6 w=10.5 l=0.15
C0 a_n73_n1050# a_n33_n1147# 0.065f
C1 w_n211_n1269# a_n33_n1147# 0.242f
C2 a_n33_n1147# a_15_n1050# 0.065f
C3 a_n73_n1050# w_n211_n1269# 0.661f
C4 a_n73_n1050# a_15_n1050# 1.67f
C5 w_n211_n1269# a_15_n1050# 0.661f
C6 a_15_n1050# VSUBS 0.434f
C7 a_n73_n1050# VSUBS 0.434f
C8 a_n33_n1147# VSUBS 0.129f
C9 w_n211_n1269# VSUBS 4.56f
.ends

.subckt sky130_fd_pr__pfet_01v8_6M437L a_n1108_n42# a_1050_n42# a_n1050_n139# w_n1246_n261#
+ VSUBS
X0 a_1050_n42# a_n1050_n139# a_n1108_n42# w_n1246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=10.5
C0 a_n1108_n42# a_n1050_n139# 0.0251f
C1 w_n1246_n261# a_n1050_n139# 3.36f
C2 a_n1050_n139# a_1050_n42# 0.0251f
C3 a_n1108_n42# w_n1246_n261# 0.0498f
C4 w_n1246_n261# a_1050_n42# 0.0498f
C5 a_1050_n42# VSUBS 0.0428f
C6 a_n1108_n42# VSUBS 0.0428f
C7 a_n1050_n139# VSUBS 2.7f
C8 w_n1246_n261# VSUBS 5.27f
.ends

.subckt sky130_fd_pr__nfet_01v8_A5ES5P a_n73_n1000# a_15_n1000# a_n33_n1088# a_n175_n1174#
X0 a_15_n1000# a_n33_n1088# a_n73_n1000# a_n175_n1174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.6 as=2.9 ps=20.6 w=10 l=0.15
C0 a_15_n1000# a_n73_n1000# 1.59f
C1 a_n33_n1088# a_n73_n1000# 0.0649f
C2 a_15_n1000# a_n33_n1088# 0.0649f
C3 a_15_n1000# a_n175_n1174# 1.04f
C4 a_n73_n1000# a_n175_n1174# 1.04f
C5 a_n33_n1088# a_n175_n1174# 0.359f
.ends

.subckt th15 Vout Vin m1_1074_6# m1_915_n714# Vp m1_4024_602# Vn m1_1076_814#
XXM0 m1_915_n714# Vn Vn Vp Vn sky130_fd_pr__pfet_01v8_MYW2PY
XXM1 m1_1074_6# m1_915_n714# Vn Vin sky130_fd_pr__nfet_01v8_JRGCPP
XXM2 m1_1076_814# m1_1074_6# Vn Vin sky130_fd_pr__nfet_01v8_JRGCPP
XXM3 m1_1076_814# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_XJ78MR
XXM4 Vp m1_4024_602# m1_1076_814# Vp Vn sky130_fd_pr__pfet_01v8_6M437L
XXM5 Vn Vout m1_1076_814# Vn sky130_fd_pr__nfet_01v8_A5ES5P
XXM7 m1_4024_602# Vout m1_1076_814# Vp Vn sky130_fd_pr__pfet_01v8_6M437L
C0 Vin m1_1076_814# 0.6f
C1 m1_915_n714# m1_1074_6# 0.0137f
C2 m1_4024_602# Vp 0.404f
C3 Vout m1_4024_602# 0.00816f
C4 m1_915_n714# m1_1076_814# 3.02e-20
C5 Vout Vp 0.129f
C6 Vp m1_1074_6# 0.0774f
C7 m1_4024_602# m1_1076_814# 0.999f
C8 Vp m1_1076_814# 1.22f
C9 Vout m1_1076_814# 0.214f
C10 Vin m1_915_n714# 0.378f
C11 m1_1074_6# m1_1076_814# 0.0103f
C12 m1_4024_602# Vin 1.79e-19
C13 Vin Vp 0.222f
C14 Vin m1_1074_6# 1.03f
C15 m1_915_n714# Vp 0.596f
C16 Vin Vn 11.5f
C17 Vout Vn 1.46f
C18 m1_4024_602# Vn 0.411f
C19 Vp Vn 18.4f
C20 m1_1076_814# Vn 6.13f
C21 m1_915_n714# Vn 1.17f
C22 m1_1074_6# Vn 0.844f
.ends

.subckt sky130_fd_pr__nfet_01v8_42G4RD a_n80_n42# a_n33_n130# a_n182_n216# a_22_n42#
X0 a_22_n42# a_n33_n130# a_n80_n42# a_n182_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_n33_n130# a_n80_n42# 0.00866f
C1 a_22_n42# a_n33_n130# 0.00866f
C2 a_22_n42# a_n80_n42# 0.0604f
C3 a_22_n42# a_n182_n216# 0.0785f
C4 a_n80_n42# a_n182_n216# 0.0785f
C5 a_n33_n130# a_n182_n216# 0.341f
.ends

.subckt sky130_fd_pr__pfet_01v8_DDPLQ8 a_n77_n42# w_n215_n261# a_n33_n139# a_19_n42#
+ VSUBS
X0 a_19_n42# a_n33_n139# a_n77_n42# w_n215_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_19_n42# a_n33_n139# 0.0127f
C1 w_n215_n261# a_n33_n139# 0.234f
C2 a_19_n42# a_n77_n42# 0.0641f
C3 a_n77_n42# w_n215_n261# 0.0484f
C4 a_n77_n42# a_n33_n139# 0.0127f
C5 a_19_n42# w_n215_n261# 0.0484f
C6 a_19_n42# VSUBS 0.0275f
C7 a_n77_n42# VSUBS 0.0275f
C8 a_n33_n139# VSUBS 0.119f
C9 w_n215_n261# VSUBS 1.04f
.ends

.subckt sky130_fd_pr__nfet_01v8_VWP3K3 a_n33_n130# a_15_n42# a_n175_n216# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
C0 a_n33_n130# a_n73_n42# 0.0209f
C1 a_15_n42# a_n33_n130# 0.0209f
C2 a_15_n42# a_n73_n42# 0.0699f
C3 a_15_n42# a_n175_n216# 0.0729f
C4 a_n73_n42# a_n175_n216# 0.0729f
C5 a_n33_n130# a_n175_n216# 0.338f
.ends

.subckt sky130_fd_pr__pfet_01v8_LZD9A4 a_n80_n42# a_22_n42# a_n33_n139# w_n218_n261#
+ VSUBS
X0 a_22_n42# a_n33_n139# a_n80_n42# w_n218_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.22
C0 a_22_n42# a_n33_n139# 0.0084f
C1 w_n218_n261# a_n33_n139# 0.233f
C2 a_22_n42# a_n80_n42# 0.0604f
C3 a_n80_n42# w_n218_n261# 0.0496f
C4 a_n80_n42# a_n33_n139# 0.0084f
C5 a_22_n42# w_n218_n261# 0.0496f
C6 a_22_n42# VSUBS 0.0285f
C7 a_n80_n42# VSUBS 0.0285f
C8 a_n33_n139# VSUBS 0.122f
C9 w_n218_n261# VSUBS 1.06f
.ends

.subckt sky130_fd_pr__nfet_01v8_VRD6K3 a_n77_n42# a_n33_n130# a_19_n42# a_n179_n216#
X0 a_19_n42# a_n33_n130# a_n77_n42# a_n179_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.19
C0 a_n33_n130# a_n77_n42# 0.0136f
C1 a_19_n42# a_n33_n130# 0.0136f
C2 a_19_n42# a_n77_n42# 0.0641f
C3 a_19_n42# a_n179_n216# 0.0763f
C4 a_n77_n42# a_n179_n216# 0.0763f
C5 a_n33_n130# a_n179_n216# 0.339f
.ends

.subckt th04 Vp V04 Vin Vn m1_397_n357# m1_960_n972#
XXM0 m1_960_n972# Vin Vn Vn sky130_fd_pr__nfet_01v8_42G4RD
XXM1 m1_397_n357# Vp Vin m1_960_n972# Vn sky130_fd_pr__pfet_01v8_DDPLQ8
XXM2 Vp m1_397_n357# Vn Vp sky130_fd_pr__nfet_01v8_VWP3K3
XXM3 Vp V04 m1_960_n972# Vp Vn sky130_fd_pr__pfet_01v8_LZD9A4
XXM4 V04 m1_960_n972# Vn Vn sky130_fd_pr__nfet_01v8_VRD6K3
C0 Vp Vn 0.228f
C1 V04 Vin 5.12e-19
C2 V04 Vn 0.181f
C3 Vn Vin 0.0911f
C4 m1_960_n972# m1_397_n357# 0.027f
C5 Vp m1_397_n357# 0.401f
C6 m1_960_n972# Vp 0.257f
C7 m1_397_n357# V04 0.0695f
C8 m1_960_n972# V04 0.39f
C9 m1_397_n357# Vin 0.109f
C10 m1_960_n972# Vin 0.395f
C11 Vp V04 0.173f
C12 m1_397_n357# Vn 0.0588f
C13 m1_960_n972# Vn 0.346f
C14 Vp Vin 0.103f
C15 Vin 0 0.599f
C16 Vn 0 0.213f
C17 V04 0 0.324f
C18 m1_960_n972# 0 0.53f
C19 Vp 0 2.61f
C20 m1_397_n357# 0 0.189f
.ends

.subckt sky130_fd_pr__pfet_01v8_PZD9SE a_n112_n139# w_n308_n261# a_112_n42# a_n170_n42#
+ VSUBS
X0 a_112_n42# a_n112_n139# a_n170_n42# w_n308_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.12
C0 a_n112_n139# a_n170_n42# 0.0153f
C1 w_n308_n261# a_n112_n139# 0.472f
C2 w_n308_n261# a_n170_n42# 0.0499f
C3 a_112_n42# a_n112_n139# 0.0153f
C4 a_112_n42# a_n170_n42# 0.0219f
C5 a_112_n42# w_n308_n261# 0.0499f
C6 a_112_n42# VSUBS 0.0318f
C7 a_n170_n42# VSUBS 0.0318f
C8 a_n112_n139# VSUBS 0.332f
C9 w_n308_n261# VSUBS 1.43f
.ends

.subckt sky130_fd_pr__nfet_01v8_UNLS3X a_n33_n200# a_n175_n286# a_n73_n112# a_15_n112#
X0 a_15_n112# a_n33_n200# a_n73_n112# a_n175_n286# sky130_fd_pr__nfet_01v8 ad=0.325 pd=2.82 as=0.325 ps=2.82 w=1.12 l=0.15
C0 a_n73_n112# a_15_n112# 0.181f
C1 a_n33_n200# a_n73_n112# 0.0262f
C2 a_n33_n200# a_15_n112# 0.0262f
C3 a_15_n112# a_n175_n286# 0.144f
C4 a_n73_n112# a_n175_n286# 0.144f
C5 a_n33_n200# a_n175_n286# 0.344f
.ends

.subckt th05 Vp V05 Vin m1_836_n724# Vn
XXM0 m1_836_n724# Vn Vn Vin sky130_fd_pr__nfet_01v8_ATLS57
XXM1 m1_836_n724# Vp Vin Vp Vn sky130_fd_pr__pfet_01v8_VZ9GC6
XXM2 m1_836_n724# Vp V05 Vp Vn sky130_fd_pr__pfet_01v8_PZD9SE
XXM3 m1_836_n724# Vn Vn V05 sky130_fd_pr__nfet_01v8_UNLS3X
C0 V05 Vp 0.103f
C1 Vin Vp 0.324f
C2 V05 m1_836_n724# 0.122f
C3 Vin m1_836_n724# 0.185f
C4 Vp m1_836_n724# 0.372f
C5 Vin V05 5.09e-20
C6 m1_836_n724# Vn 1.23f
C7 V05 Vn 0.48f
C8 Vin Vn 1.06f
C9 Vp Vn 3.53f
.ends

.subckt analog_therm
Xth09_0 th09_0/V09 x30/Vin th09_0/m1_891_n977# x31/Vp th09_0/m1_1725_85# VSUBS th09
Xx30 x31/Vp x30/Vin VSUBS VSUBS preamp
Xx31 x31/Vp VSUBS x31/Vout x31/m1_931_n929# VSUBS th01
Xx20 x31/Vp x30/Vin x20/V06 x20/m1_528_n874# VSUBS th06
Xx21 x30/Vin x21/V07 x31/Vp x21/m1_400_n1066# VSUBS th07
Xx22 x22/V08 x30/Vin x22/m1_451_n1105# x31/Vp VSUBS th08
Xx24 x24/V10 x30/Vin x24/m1_718_n418# x31/Vp VSUBS x24/m1_878_n414# th10
Xx25 x25/V11 x30/Vin x31/Vp x25/m1_717_301# x25/m1_509_303# VSUBS th11
Xx26 x26/Vout x30/Vin x26/m1_532_n361# x31/Vp x26/m1_773_n853# VSUBS th12
Xx27 x27/Vout x30/Vin x27/m1_724_n958# x27/m1_546_n454# x31/Vp VSUBS th13
Xx16 x16/Vout VSUBS x31/Vp x16/m1_4146_502# x30/Vin x16/m1_1199_9# th02
Xx28 x30/Vin x28/m1_1594_n962# x28/Vout x31/Vp x28/m1_710_n388# x28/m1_2498_n384#
+ VSUBS th14
Xx17 x31/Vp x17/Vout x30/Vin x17/m1_782_n682# VSUBS x17/li_1010_10# x17/m1_522_n210#
+ th03
Xtherm_0 therm_0/b[0] therm_0/b[1] therm_0/b[2] therm_0/b[3] x31/Vout x25/V11 x26/Vout
+ x27/Vout x28/Vout x29/Vout x16/Vout x17/Vout x18/V04 x19/V05 x20/V06 x21/V07 x22/V08
+ th09_0/V09 therm_0/net7 therm_0/_04_ therm_0/net19 therm_0/net15 therm_0/net14 therm_0/_31_/a_35_297#
+ therm_0/input7/a_27_47# therm_0/_27_/a_27_297# therm_0/input1/a_75_212# therm_0/input5/a_62_47#
+ therm_0/net2 therm_0/input5/a_841_47# therm_0/_19_ therm_0/net8 therm_0/_17_ therm_0/_01_
+ therm_0/_44_/a_250_297# x24/V10 therm_0/input15/a_27_47# therm_0/_20_ therm_0/_14_
+ therm_0/net1 therm_0/_16_ therm_0/net9 x31/Vp therm_0/net5 VSUBS therm_0/_29_/a_29_53#
+ therm
Xx29 x29/Vout x30/Vin x29/m1_1074_6# x29/m1_915_n714# x31/Vp x29/m1_4024_602# VSUBS
+ x29/m1_1076_814# th15
Xx18 x31/Vp x18/V04 x30/Vin VSUBS x18/m1_397_n357# x18/m1_960_n972# th04
Xx19 x31/Vp x19/V05 x30/Vin x19/m1_836_n724# VSUBS th05
C0 x18/m1_960_n972# x25/V11 0.00234f
C1 x27/m1_546_n454# x29/Vout 0.0022f
C2 x16/m1_4146_502# x24/V10 1.32e-19
C3 x25/V11 therm_0/_19_ 4.44e-34
C4 x29/Vout x26/Vout 2.47e-19
C5 x19/V05 x30/Vin 0.0106f
C6 x18/m1_397_n357# x18/V04 0.00319f
C7 x28/m1_710_n388# x26/m1_532_n361# 1.3e-19
C8 x21/V07 x30/Vin 0.0713f
C9 x21/V07 x25/V11 0.0109f
C10 x31/Vp x25/m1_717_301# 5.4e-19
C11 x29/m1_1076_814# x30/Vin 0.282f
C12 x31/Vp th09_0/m1_891_n977# 0.0806f
C13 therm_0/b[3] x28/m1_710_n388# 2.33e-20
C14 x24/V10 x30/Vin 0.245f
C15 x24/V10 x25/V11 2.43f
C16 x22/V08 x20/V06 4.14f
C17 x29/Vout x24/m1_718_n418# 1.86e-20
C18 x17/m1_782_n682# x18/V04 0.0273f
C19 x17/m1_522_n210# x18/V04 0.0112f
C20 x21/m1_400_n1066# x30/Vin 0.0261f
C21 x31/Vp x18/m1_397_n357# 0.0139f
C22 x28/m1_710_n388# x27/Vout 9.44e-20
C23 x22/m1_451_n1105# x17/Vout 0.00533f
C24 x17/m1_782_n682# x17/Vout 0.0227f
C25 x17/Vout x17/m1_522_n210# 0.00497f
C26 x21/m1_400_n1066# x25/V11 0.0121f
C27 x27/m1_724_n958# x31/Vp 5.68e-32
C28 x29/m1_1076_814# th09_0/V09 1.54e-19
C29 x31/Vp x29/m1_915_n714# 0.0064f
C30 x31/m1_931_n929# x18/V04 0.0419f
C31 x19/V05 x22/V08 9.26e-19
C32 x31/Vp therm_0/net7 0.00165f
C33 x28/m1_710_n388# x28/Vout 0.00283f
C34 x31/m1_931_n929# x16/Vout 0.0294f
C35 x31/m1_931_n929# x17/Vout 0.00136f
C36 x29/m1_4024_602# x30/Vin 0.0183f
C37 x21/V07 x22/V08 1.75f
C38 x27/m1_724_n958# th09_0/m1_891_n977# 0.00391f
C39 x31/Vout x20/V06 4.62e-19
C40 x17/li_1010_10# x30/Vin 0.0107f
C41 x31/Vp x26/m1_773_n853# 0.00752f
C42 x28/m1_2498_n384# x28/Vout 0.0172f
C43 x31/Vp x26/m1_532_n361# 0.0972f
C44 x22/m1_451_n1105# x31/Vp 0.0149f
C45 x20/m1_528_n874# x19/m1_836_n724# 0.00244f
C46 x17/m1_782_n682# x31/Vp 0.0227f
C47 x16/m1_4146_502# x28/m1_710_n388# 0.00123f
C48 x17/m1_522_n210# x31/Vp 0.0183f
C49 x31/Vp x16/m1_1199_9# 0.0353f
C50 therm_0/net14 x26/Vout 5.54e-21
C51 x31/Vp therm_0/b[3] 9.65e-20
C52 therm_0/_04_ x25/V11 4.44e-34
C53 x24/V10 x26/Vout 2.44f
C54 x16/m1_4146_502# x28/m1_2498_n384# 1.09e-21
C55 x31/m1_931_n929# x31/Vp 0.00892f
C56 x31/Vout x19/V05 3.47e-19
C57 x20/m1_528_n874# x20/V06 0.0131f
C58 x25/m1_509_303# x30/Vin 0.0113f
C59 x19/m1_836_n724# x20/V06 4.12e-19
C60 x31/Vout x21/V07 0.015f
C61 x28/m1_710_n388# x30/Vin 0.00118f
C62 x16/m1_4146_502# x18/V04 0.0381f
C63 x25/m1_509_303# x25/V11 0.00588f
C64 x31/Vp x27/Vout 0.0629f
C65 x16/Vout x16/m1_4146_502# 0.103f
C66 x28/m1_710_n388# x25/V11 0.00354f
C67 th09_0/m1_1725_85# x30/Vin 0.054f
C68 x17/Vout x16/m1_4146_502# 3.37e-19
C69 x18/m1_397_n357# x26/m1_532_n361# 6.58e-20
C70 x29/m1_1076_814# x29/Vout 0.00808f
C71 x18/m1_397_n357# x16/m1_1199_9# 0.0133f
C72 x24/m1_878_n414# x29/m1_1076_814# 2e-20
C73 x24/V10 x24/m1_718_n418# 0.00674f
C74 therm_0/net2 x28/Vout -3.55e-33
C75 x20/m1_528_n874# x19/V05 0.0275f
C76 x28/m1_2498_n384# x25/V11 2.83e-19
C77 x17/li_1010_10# x22/V08 0.00638f
C78 x24/V10 x29/Vout 0.0827f
C79 x31/Vp x28/Vout 0.0137f
C80 x19/m1_836_n724# x19/V05 0.00448f
C81 th09_0/m1_891_n977# x27/Vout 2.75e-20
C82 x30/Vin x18/V04 0.377f
C83 x20/m1_528_n874# x21/V07 3.47e-19
C84 x17/Vout x30/Vin 0.00929f
C85 x25/V11 x18/V04 0.0147f
C86 th09_0/V09 x28/m1_710_n388# 0.00165f
C87 x21/m1_400_n1066# x24/m1_718_n418# 1.03e-19
C88 x16/Vout x25/V11 0.00589f
C89 x31/Vp x16/m1_4146_502# 0.0101f
C90 x19/V05 x20/V06 6.37f
C91 therm_0/net15 x25/V11 1.78e-33
C92 x17/m1_782_n682# x22/m1_451_n1105# 0.00574f
C93 x21/V07 x20/V06 0.504f
C94 therm_0/b[1] x31/Vp 0.126f
C95 x19/m1_836_n724# x21/m1_400_n1066# 2.51e-19
C96 x29/m1_4024_602# x29/Vout 1.91e-20
C97 x27/m1_546_n454# x28/m1_710_n388# 0.00137f
C98 therm_0/_01_ x25/V11 -1.39e-35
C99 x31/Vp x30/Vin 3.85f
C100 x21/V07 x18/m1_960_n972# 0.00331f
C101 x26/Vout x28/m1_710_n388# 0.18f
C102 x27/m1_546_n454# th09_0/m1_1725_85# 2.12e-19
C103 x31/Vp x25/V11 0.826f
C104 x21/V07 x19/V05 0.119f
C105 x24/V10 x18/m1_960_n972# 4.66e-20
C106 x26/Vout x28/m1_2498_n384# 0.0316f
C107 x22/V08 x18/V04 0.0619f
C108 x25/m1_717_301# x30/Vin 0.031f
C109 th09_0/m1_891_n977# x30/Vin 0.055f
C110 x16/Vout x22/V08 0.00194f
C111 x17/Vout x22/V08 4.2f
C112 x18/m1_960_n972# x21/m1_400_n1066# 0.00136f
C113 x25/m1_509_303# x24/m1_718_n418# 1.64e-19
C114 therm_0/input5/a_62_47# therm_0/net2 7.11e-33
C115 x21/V07 x24/V10 6.04e-19
C116 x31/Vp th09_0/V09 0.0955f
C117 x25/m1_509_303# x24/m1_878_n414# 6.26e-20
C118 x29/Vout x28/m1_710_n388# 0.0466f
C119 therm_0/net15 x26/Vout -5.55e-35
C120 x18/m1_397_n357# x30/Vin 0.00521f
C121 th09_0/m1_1725_85# x29/Vout 5.9e-19
C122 therm_0/b[3] x28/Vout 0.00935f
C123 x31/Vp therm_0/input7/a_27_47# 1.23e-19
C124 x17/li_1010_10# x20/V06 7.81e-19
C125 x18/m1_397_n357# x25/V11 0.00418f
C126 x27/m1_724_n958# x30/Vin 1.49e-19
C127 x21/V07 x21/m1_400_n1066# 0.00822f
C128 x29/Vout x28/m1_2498_n384# 0.00317f
C129 x31/Vp x28/m1_1594_n962# -1.14e-31
C130 th09_0/V09 th09_0/m1_891_n977# 0.00797f
C131 x29/m1_915_n714# x30/Vin 0.0157f
C132 x31/Vout x18/V04 0.192f
C133 x31/Vp x22/V08 0.156f
C134 x25/m1_509_303# x19/m1_836_n724# 7.72e-20
C135 x16/Vout x31/Vout 0.324f
C136 x17/li_1010_10# x18/m1_960_n972# 5.11e-19
C137 x31/Vout x17/Vout 0.0189f
C138 x24/V10 x21/m1_400_n1066# 5.83e-19
C139 x27/m1_546_n454# x31/Vp 0.00653f
C140 therm_0/net2 x26/Vout 3.36e-20
C141 x27/Vout x28/Vout 3.68e-20
C142 x31/Vp x26/Vout 0.58f
C143 x31/m1_931_n929# x16/m1_4146_502# 0.00436f
C144 th09_0/m1_891_n977# x28/m1_1594_n962# 1.28e-19
C145 x26/m1_773_n853# x30/Vin 0.00934f
C146 x17/li_1010_10# x19/V05 5.78e-19
C147 x26/m1_532_n361# x30/Vin 0.0277f
C148 x17/m1_782_n682# x30/Vin 0.00792f
C149 x22/m1_451_n1105# x30/Vin 0.00108f
C150 x17/m1_522_n210# x30/Vin 0.0401f
C151 x17/li_1010_10# x21/V07 0.0726f
C152 x30/Vin x16/m1_1199_9# 0.016f
C153 x26/m1_532_n361# x25/V11 3.91e-19
C154 x27/m1_546_n454# th09_0/m1_891_n977# 0.00251f
C155 therm_0/input15/a_27_47# x24/V10 -5.55e-35
C156 x27/m1_724_n958# th09_0/V09 0.0274f
C157 x25/V11 x16/m1_1199_9# 0.00558f
C158 x31/Vout x31/Vp 2.9e-19
C159 x31/m1_931_n929# x30/Vin 1.36e-19
C160 x31/Vp x24/m1_718_n418# 0.0302f
C161 x31/Vp x29/Vout 0.149f
C162 therm_0/net7 therm_0/input7/a_27_47# -1.42e-32
C163 x31/Vp therm_0/_31_/a_35_297# -1.42e-32
C164 x24/m1_878_n414# x31/Vp 0.00965f
C165 x20/V06 x18/V04 0.00318f
C166 x27/Vout x30/Vin 0.003f
C167 x17/Vout x20/V06 5.65e-20
C168 x27/m1_546_n454# x27/m1_724_n958# -3.55e-33
C169 therm_0/b[1] x28/Vout -1.39e-35
C170 x29/Vout th09_0/m1_891_n977# 0.0143f
C171 x20/m1_528_n874# x31/Vp 0.0171f
C172 x18/m1_960_n972# x18/V04 0.0335f
C173 x24/m1_878_n414# x25/m1_717_301# 0.00464f
C174 x25/m1_509_303# x24/V10 5.66e-20
C175 x31/Vp x19/m1_836_n724# 0.0398f
C176 x28/Vout x30/Vin 3.57e-21
C177 x24/V10 x28/m1_710_n388# 0.00796f
C178 th09_0/m1_1725_85# x29/m1_1076_814# 2.08e-20
C179 x17/m1_782_n682# x22/V08 0.00308f
C180 x25/V11 x28/Vout 0.0212f
C181 x22/m1_451_n1105# x22/V08 0.0109f
C182 x17/m1_522_n210# x22/V08 2.24e-20
C183 x19/V05 x18/V04 0.00182f
C184 therm_0/b[1] x16/m1_4146_502# 2.77e-19
C185 x17/Vout x19/V05 4.32e-20
C186 x24/V10 x28/m1_2498_n384# 0.00279f
C187 x21/V07 x18/V04 0.862f
C188 x26/Vout x26/m1_532_n361# 0.0135f
C189 x16/m1_4146_502# x30/Vin 0.0896f
C190 th09_0/V09 x27/Vout 0.283f
C191 x31/Vp x20/V06 0.336f
C192 x16/Vout x21/V07 0.00662f
C193 x17/Vout x21/V07 1.53f
C194 x26/Vout x16/m1_1199_9# 2.37e-19
C195 x31/m1_931_n929# x22/V08 0.00102f
C196 x16/m1_4146_502# x25/V11 0.0133f
C197 x24/V10 x18/V04 5.08e-19
C198 therm_0/b[3] x26/Vout 2.96e-20
C199 x31/Vp x18/m1_960_n972# 0.00326f
C200 th09_0/V09 x28/Vout 6.29e-19
C201 x26/m1_773_n853# x24/m1_718_n418# 3.69e-21
C202 x21/m1_400_n1066# x18/V04 0.00623f
C203 x31/Vp x19/V05 0.507f
C204 x27/m1_546_n454# x27/Vout 0.11f
C205 x26/m1_532_n361# x24/m1_718_n418# 3.04e-19
C206 x25/V11 x30/Vin 0.666f
C207 x17/Vout x21/m1_400_n1066# 3.02e-21
C208 x31/Vp x21/V07 0.28f
C209 therm_0/input5/a_841_47# x28/Vout -2.78e-35
C210 x31/m1_931_n929# x31/Vout 0.0105f
C211 x31/Vp therm_0/_29_/a_29_53# -1.42e-32
C212 x31/Vp x29/m1_1076_814# 0.666f
C213 therm_0/_44_/a_250_297# x26/Vout 1.9e-20
C214 x27/m1_546_n454# x28/Vout 2.24e-19
C215 x31/Vp x24/V10 0.66f
C216 x26/Vout x28/Vout 0.194f
C217 x17/li_1010_10# x18/V04 0.0485f
C218 x29/m1_1076_814# th09_0/m1_891_n977# 0.00205f
C219 th09_0/V09 x30/Vin 0.111f
C220 x17/li_1010_10# x17/Vout 0.0881f
C221 x31/Vp x21/m1_400_n1066# 0.0116f
C222 x29/Vout x27/Vout 0.00204f
C223 x16/m1_4146_502# x26/Vout 1.07e-19
C224 x21/V07 x18/m1_397_n357# 0.0021f
C225 x28/m1_1594_n962# x30/Vin 0.00819f
C226 x17/m1_782_n682# x20/V06 9.22e-20
C227 x22/m1_451_n1105# x20/V06 0.00567f
C228 x22/V08 x30/Vin 0.00289f
C229 x29/Vout x28/Vout 0.0211f
C230 x31/Vp x29/m1_4024_602# 0.0611f
C231 x27/m1_546_n454# x30/Vin 0.00347f
C232 x18/m1_960_n972# x26/m1_532_n361# 1.89e-20
C233 x31/Vout x16/m1_4146_502# 4.17e-20
C234 x17/m1_782_n682# x18/m1_960_n972# 1.3e-19
C235 therm_0/net5 therm_0/net2 -7.11e-33
C236 x26/Vout x30/Vin 0.377f
C237 x31/m1_931_n929# x20/V06 7.88e-19
C238 x17/li_1010_10# x31/Vp 0.0865f
C239 x16/Vout x28/m1_710_n388# 1.55e-19
C240 x18/m1_960_n972# x16/m1_1199_9# 0.0015f
C241 x26/Vout x25/V11 0.00131f
C242 x17/m1_782_n682# x19/V05 7.06e-20
C243 x22/m1_451_n1105# x19/V05 3.42e-19
C244 x18/m1_397_n357# x21/m1_400_n1066# 7.85e-19
C245 x29/m1_4024_602# th09_0/m1_891_n977# 5.01e-20
C246 th09_0/V09 x28/m1_1594_n962# 1.16e-19
C247 x22/m1_451_n1105# x21/V07 0.013f
C248 x17/m1_782_n682# x21/V07 0.0449f
C249 x29/m1_1076_814# x26/m1_773_n853# 1.86e-20
C250 x17/m1_522_n210# x21/V07 0.00528f
C251 therm_0/net1 x31/Vp 2.5e-19
C252 x29/m1_1076_814# x26/m1_532_n361# 0.00108f
C253 x24/V10 x26/m1_773_n853# 0.00125f
C254 x29/m1_1074_6# x30/Vin 0.00242f
C255 x31/m1_931_n929# x19/V05 6.06e-19
C256 x16/Vout x18/V04 0.0705f
C257 x24/V10 x26/m1_532_n361# 0.0267f
C258 x17/Vout x18/V04 3.29f
C259 x27/m1_546_n454# th09_0/V09 0.0457f
C260 x24/m1_718_n418# x30/Vin 0.0179f
C261 x25/m1_509_303# x31/Vp 0.0212f
C262 x29/Vout x30/Vin 0.388f
C263 x16/Vout x17/Vout 0.0964f
C264 x24/V10 x16/m1_1199_9# 3.37e-19
C265 x31/Vp x28/m1_710_n388# 0.317f
C266 x31/m1_931_n929# x21/V07 0.0217f
C267 x24/m1_878_n414# x30/Vin 0.0194f
C268 x25/V11 x24/m1_718_n418# 0.0105f
C269 therm_0/b[3] x24/V10 0.016f
C270 x31/Vp th09_0/m1_1725_85# 0.0294f
C271 x24/m1_878_n414# x25/V11 5.31e-19
C272 x22/m1_451_n1105# x21/m1_400_n1066# 1.15e-21
C273 x31/Vp x28/m1_2498_n384# 0.00561f
C274 x26/Vout x28/m1_1594_n962# 0.00132f
C275 x20/m1_528_n874# x30/Vin 0.00779f
C276 therm_0/_27_/a_27_297# x25/V11 -1.11e-34
C277 x19/m1_836_n724# x30/Vin 0.0152f
C278 therm_0/input1/a_75_212# x31/Vp 6.38e-19
C279 x31/Vp x18/V04 0.464f
C280 x19/m1_836_n724# x25/V11 2.28e-20
C281 x31/Vp therm_0/net8 2.87e-21
C282 x16/Vout x31/Vp 0.109f
C283 x17/Vout x31/Vp 0.263f
C284 x29/Vout th09_0/V09 1.53f
C285 x20/V06 x30/Vin 0.00618f
C286 x17/m1_782_n682# x17/li_1010_10# 2.84e-32
C287 x22/m1_451_n1105# x17/li_1010_10# 0.00327f
C288 x31/Vout x22/V08 6.17e-19
C289 therm_0/net9 x31/Vp 2.84e-32
C290 x24/V10 x28/Vout 0.102f
C291 x25/m1_509_303# x29/m1_915_n714# 7.46e-21
C292 x27/m1_724_n958# x28/m1_710_n388# 5.19e-20
C293 x21/V07 x16/m1_4146_502# 4.29e-19
C294 x29/Vout x28/m1_1594_n962# 0.0144f
C295 x18/m1_960_n972# x30/Vin 0.00703f
C296 x31/Vp therm_0/_01_ -1.14e-31
C297 x19/m1_836_n724# VSUBS 1.03f
C298 x19/V05 VSUBS 6.75f
C299 x18/V04 VSUBS 4.74f
C300 x18/m1_960_n972# VSUBS 0.548f
C301 x18/m1_397_n357# VSUBS 0.204f
C302 x29/Vout VSUBS 3.92f
C303 x29/m1_4024_602# VSUBS 0.411f
C304 x29/m1_1076_814# VSUBS 6.09f
C305 x29/m1_915_n714# VSUBS 1.1f
C306 x29/m1_1074_6# VSUBS 0.644f
C307 therm_0/_03_ VSUBS 0.36f
C308 therm_0/net10 VSUBS 0.458f
C309 therm_0/_30_/a_109_53# VSUBS 0.159f
C310 therm_0/_30_/a_215_297# VSUBS 0.142f
C311 therm_0/_05_ VSUBS 0.152f
C312 therm_0/net8 VSUBS 0.386f
C313 therm_0/_31_/a_285_297# VSUBS 0.00137f
C314 therm_0/_31_/a_35_297# VSUBS 0.255f
C315 therm_0/_32_/a_27_47# VSUBS 0.175f
C316 therm_0/_50_/a_343_93# VSUBS 0.172f
C317 therm_0/_50_/a_223_47# VSUBS 0.141f
C318 therm_0/_50_/a_27_47# VSUBS 0.259f
C319 therm_0/_07_ VSUBS 0.288f
C320 therm_0/_06_ VSUBS 0.819f
C321 therm_0/net13 VSUBS 0.379f
C322 therm_0/_33_/a_209_311# VSUBS 0.143f
C323 therm_0/_33_/a_109_93# VSUBS 0.158f
C324 therm_0/net12 VSUBS 0.529f
C325 therm_0/_34_/a_285_47# VSUBS 0.0174f
C326 therm_0/_34_/a_47_47# VSUBS 0.199f
C327 therm_0/_23_ VSUBS 0.106f
C328 therm_0/input15/a_27_47# VSUBS 0.208f
C329 therm_0/_09_ VSUBS 0.149f
C330 therm_0/_08_ VSUBS 0.131f
C331 therm_0/_35_/a_489_413# VSUBS 0.0254f
C332 therm_0/_35_/a_226_47# VSUBS 0.162f
C333 therm_0/_35_/a_76_199# VSUBS 0.141f
C334 therm_0/_24_ VSUBS 0.135f
C335 therm_0/_12_ VSUBS 0.387f
C336 therm_0/_52_/a_250_297# VSUBS 0.0278f
C337 therm_0/_52_/a_93_21# VSUBS 0.151f
C338 therm_0/_10_ VSUBS 0.643f
C339 therm_0/_36_/a_27_47# VSUBS 0.175f
C340 therm_0/input14/a_27_47# VSUBS 0.208f
C341 therm_0/_53_/a_29_53# VSUBS 0.18f
C342 therm_0/_11_ VSUBS 0.267f
C343 therm_0/_37_/a_27_47# VSUBS 0.175f
C344 therm_0/input13/a_27_47# VSUBS 0.208f
C345 therm_0/net18 VSUBS 0.207f
C346 therm_0/_25_ VSUBS 0.191f
C347 therm_0/_54_/a_75_212# VSUBS 0.21f
C348 therm_0/_38_/a_27_47# VSUBS 0.175f
C349 therm_0/net19 VSUBS 0.177f
C350 therm_0/_22_ VSUBS 0.216f
C351 therm_0/_14_ VSUBS 0.228f
C352 therm_0/_15_ VSUBS 0.338f
C353 therm_0/_55_/a_217_297# VSUBS 0.00117f
C354 therm_0/_55_/a_80_21# VSUBS 0.21f
C355 therm_0/input12/a_27_47# VSUBS 0.208f
C356 therm_0/net9 VSUBS 0.306f
C357 therm_0/input9/a_75_212# VSUBS 0.21f
C358 therm_0/_39_/a_285_47# VSUBS 0.0174f
C359 therm_0/_39_/a_47_47# VSUBS 0.199f
C360 therm_0/net11 VSUBS 0.771f
C361 therm_0/input11/a_27_47# VSUBS 0.208f
C362 therm_0/input8/a_27_47# VSUBS 0.208f
C363 therm_0/input10/a_27_47# VSUBS 0.208f
C364 therm_0/net7 VSUBS 0.462f
C365 therm_0/input7/a_27_47# VSUBS 0.208f
C366 therm_0/input6/a_27_47# VSUBS 0.208f
C367 therm_0/net5 VSUBS 0.842f
C368 therm_0/input5/a_841_47# VSUBS 0.0929f
C369 therm_0/input5/a_664_47# VSUBS 0.13f
C370 therm_0/input5/a_558_47# VSUBS 0.164f
C371 therm_0/input5/a_381_47# VSUBS 0.11f
C372 therm_0/input5/a_62_47# VSUBS 0.169f
C373 therm_0/input4/a_75_212# VSUBS 0.21f
C374 therm_0/input3/a_27_47# VSUBS 0.208f
C375 therm_0/net2 VSUBS 0.668f
C376 therm_0/input2/a_27_47# VSUBS 0.208f
C377 therm_0/net1 VSUBS 0.342f
C378 therm_0/input1/a_75_212# VSUBS 0.21f
C379 therm_0/b[3] VSUBS 0.408f
C380 therm_0/output19/a_27_47# VSUBS 0.543f
C381 therm_0/b[2] VSUBS 0.515f
C382 therm_0/output18/a_27_47# VSUBS 0.543f
C383 therm_0/b[1] VSUBS 0.529f
C384 therm_0/net17 VSUBS 0.173f
C385 therm_0/output17/a_27_47# VSUBS 0.543f
C386 therm_0/_41_/a_59_75# VSUBS 0.177f
C387 therm_0/b[0] VSUBS 0.528f
C388 therm_0/output16/a_27_47# VSUBS 0.543f
C389 therm_0/_16_ VSUBS 0.125f
C390 therm_0/_42_/a_209_311# VSUBS 0.143f
C391 therm_0/_42_/a_109_93# VSUBS 0.158f
C392 therm_0/_17_ VSUBS 0.251f
C393 therm_0/_00_ VSUBS 0.377f
C394 therm_0/_43_/a_193_413# VSUBS 0.136f
C395 therm_0/_43_/a_27_47# VSUBS 0.224f
C396 therm_0/net6 VSUBS 0.532f
C397 therm_0/net4 VSUBS 0.324f
C398 therm_0/_26_/a_29_53# VSUBS 0.18f
C399 therm_0/_01_ VSUBS 0.15f
C400 therm_0/net14 VSUBS 0.516f
C401 therm_0/net3 VSUBS 0.464f
C402 therm_0/net15 VSUBS 0.452f
C403 therm_0/_27_/a_27_297# VSUBS 0.163f
C404 therm_0/_18_ VSUBS 0.143f
C405 therm_0/_44_/a_250_297# VSUBS 0.0278f
C406 therm_0/_44_/a_93_21# VSUBS 0.151f
C407 therm_0/net16 VSUBS 0.231f
C408 therm_0/_13_ VSUBS 0.133f
C409 therm_0/_45_/a_193_297# VSUBS 0.0011f
C410 therm_0/_45_/a_109_297# VSUBS 7.11e-19
C411 therm_0/_45_/a_27_47# VSUBS 0.216f
C412 therm_0/_29_/a_29_53# VSUBS 0.18f
C413 therm_0/_19_ VSUBS 0.118f
C414 therm_0/_04_ VSUBS 0.339f
C415 therm_0/_47_/a_299_297# VSUBS 0.0348f
C416 therm_0/_47_/a_81_21# VSUBS 0.147f
C417 x31/Vp VSUBS 0.134p
C418 therm_0/_48_/a_27_47# VSUBS 0.177f
C419 therm_0/_21_ VSUBS 0.29f
C420 therm_0/_20_ VSUBS 0.238f
C421 therm_0/_02_ VSUBS 0.453f
C422 therm_0/_49_/a_201_297# VSUBS 0.00345f
C423 therm_0/_49_/a_75_199# VSUBS 0.205f
C424 x17/Vout VSUBS 1.97f
C425 x17/m1_782_n682# VSUBS 1.43f
C426 x17/li_1010_10# VSUBS 2.83f
C427 x17/m1_522_n210# VSUBS 0.241f
C428 x28/Vout VSUBS 2.26f
C429 x28/m1_710_n388# VSUBS 3.53f
C430 x28/m1_2498_n384# VSUBS 0.297f
C431 x28/m1_1594_n962# VSUBS 0.299f
C432 x16/Vout VSUBS 2.48f
C433 x16/m1_4146_502# VSUBS 8.47f
C434 x16/m1_1199_9# VSUBS 0.388f
C435 x27/Vout VSUBS 3.02f
C436 x27/m1_546_n454# VSUBS 1.54f
C437 x27/m1_724_n958# VSUBS 0.188f
C438 x26/m1_532_n361# VSUBS 0.851f
C439 x26/Vout VSUBS 2.5f
C440 x26/m1_773_n853# VSUBS 0.198f
C441 x25/m1_509_303# VSUBS 0.633f
C442 x25/V11 VSUBS 2.68f
C443 x25/m1_717_301# VSUBS 0.238f
C444 x24/m1_718_n418# VSUBS 0.584f
C445 x24/V10 VSUBS 1.91f
C446 x24/m1_878_n414# VSUBS 0.172f
C447 x22/m1_451_n1105# VSUBS 0.669f
C448 x30/Vin VSUBS 38.9f
C449 x22/V08 VSUBS 2.01f
C450 x21/m1_400_n1066# VSUBS 0.769f
C451 x21/V07 VSUBS 6.52f
C452 x20/V06 VSUBS 2.53f
C453 x20/m1_528_n874# VSUBS 0.727f
C454 x31/m1_931_n929# VSUBS 2.22f
C455 x31/Vout VSUBS 2.02f
C456 th09_0/m1_891_n977# VSUBS 1.15f
C457 th09_0/V09 VSUBS 2.96f
C458 th09_0/m1_1725_85# VSUBS 0.13f
.ends

