* NGSPICE file created from th11.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_XGAKDL a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
+ VSUBS
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_15_n200# a_n73_n200# 0.321f
C1 w_n211_n419# a_n33_n297# 0.191f
C2 a_15_n200# a_n33_n297# 0.0293f
C3 a_15_n200# w_n211_n419# 0.0336f
C4 a_n73_n200# a_n33_n297# 0.0293f
C5 a_n73_n200# w_n211_n419# 0.0336f
C6 a_15_n200# VSUBS 0.164f
C7 a_n73_n200# VSUBS 0.164f
C8 a_n33_n297# VSUBS 0.147f
C9 w_n211_n419# VSUBS 1.14f
.ends

.subckt sky130_fd_pr__nfet_01v8_4X3CDA a_n306_n216# a_n180_n130# a_n238_n42# a_180_n42#
X0 a_180_n42# a_n180_n130# a_n238_n42# a_n306_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=1.8
C0 a_n180_n130# a_n238_n42# 0.0189f
C1 a_180_n42# a_n238_n42# 0.0147f
C2 a_180_n42# a_n180_n130# 0.0189f
C3 a_180_n42# a_n306_n216# 0.075f
C4 a_n238_n42# a_n306_n216# 0.075f
C5 a_n180_n130# a_n306_n216# 1.1f
.ends

.subckt sky130_fd_pr__pfet_01v8_MWB9BZ a_15_n43# w_n211_n262# a_n73_n43# a_n33_n140#
+ VSUBS
X0 a_15_n43# a_n33_n140# a_n73_n43# w_n211_n262# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1.44 as=0.125 ps=1.44 w=0.43 l=0.15
C0 a_n33_n140# a_15_n43# 0.0193f
C1 w_n211_n262# a_n73_n43# 0.0198f
C2 a_n73_n43# a_15_n43# 0.0715f
C3 w_n211_n262# a_15_n43# 0.0198f
C4 a_n33_n140# a_n73_n43# 0.0193f
C5 a_n33_n140# w_n211_n262# 0.187f
C6 a_15_n43# VSUBS 0.0453f
C7 a_n73_n43# VSUBS 0.0453f
C8 a_n33_n140# VSUBS 0.143f
C9 w_n211_n262# VSUBS 0.752f
.ends

.subckt sky130_fd_pr__pfet_01v8_JM8GTH a_50_n42# w_n246_n261# a_n50_n139# a_n108_n42#
+ VSUBS
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n246_n261# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 a_n50_n139# a_n108_n42# 0.00909f
C1 w_n246_n261# a_50_n42# 0.0224f
C2 a_50_n42# a_n108_n42# 0.0391f
C3 w_n246_n261# a_n108_n42# 0.0224f
C4 a_n50_n139# a_50_n42# 0.00909f
C5 a_n50_n139# w_n246_n261# 0.223f
C6 a_50_n42# VSUBS 0.0488f
C7 a_n108_n42# VSUBS 0.0488f
C8 a_n50_n139# VSUBS 0.209f
C9 w_n246_n261# VSUBS 0.88f
.ends

.subckt sky130_fd_pr__nfet_01v8_L9ESAD a_n175_n190# a_n73_n50# a_n33_n138# a_15_n50#
X0 a_15_n50# a_n33_n138# a_n73_n50# a_n175_n190# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
C0 a_n73_n50# a_15_n50# 0.0826f
C1 a_n33_n138# a_15_n50# 0.0216f
C2 a_n73_n50# a_n33_n138# 0.0216f
C3 a_15_n50# a_n175_n190# 0.0704f
C4 a_n73_n50# a_n175_n190# 0.0797f
C5 a_n33_n138# a_n175_n190# 0.315f
.ends

.subckt th11 Vp V11 Vin Vn
XXM0 Vn Vp Vn m1_577_n654# Vn sky130_fd_pr__pfet_01v8_XGAKDL
XXM1 Vn Vin m1_577_n654# m1_705_187# sky130_fd_pr__nfet_01v8_4X3CDA
XXM2 m1_705_187# Vp Vp Vin Vn sky130_fd_pr__pfet_01v8_MWB9BZ
XXM3 V11 Vp m1_705_187# Vp Vn sky130_fd_pr__pfet_01v8_JM8GTH
XXM4 Vn Vn m1_705_187# V11 sky130_fd_pr__nfet_01v8_L9ESAD
C0 Vin Vn 0.135f
C1 m1_577_n654# Vin 0.213f
C2 V11 Vn 0.00327f
C3 V11 m1_577_n654# 6.11e-19
C4 Vp Vn 0.0775f
C5 Vp m1_577_n654# 0.0405f
C6 m1_705_187# Vin 0.0649f
C7 V11 m1_705_187# 0.376f
C8 Vp m1_705_187# 0.286f
C9 m1_577_n654# Vn 0.0457f
C10 V11 Vin 2.69e-19
C11 Vp Vin 0.285f
C12 m1_705_187# Vn 0.463f
C13 m1_705_187# m1_577_n654# 0.0258f
C14 Vp V11 0.026f
C15 Vp 0 2.61f
C16 Vn 0 0.355f
C17 V11 0 0.404f
C18 m1_705_187# 0 0.602f
C19 m1_577_n654# 0 0.286f
C20 Vin 0 1.27f
.ends

