magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 214 29 220
rect -29 180 -17 214
rect -29 174 29 180
rect -29 -180 29 -174
rect -29 -214 -17 -180
rect -29 -220 29 -214
<< pwell >>
rect -211 -352 211 352
<< nmos >>
rect -15 -142 15 142
<< ndiff >>
rect -73 130 -15 142
rect -73 -130 -61 130
rect -27 -130 -15 130
rect -73 -142 -15 -130
rect 15 130 73 142
rect 15 -130 27 130
rect 61 -130 73 130
rect 15 -142 73 -130
<< ndiffc >>
rect -61 -130 -27 130
rect 27 -130 61 130
<< psubdiff >>
rect -175 282 -79 316
rect 79 282 175 316
rect -175 220 -141 282
rect 141 220 175 282
rect -175 -282 -141 -220
rect 141 -282 175 -220
rect -175 -316 -79 -282
rect 79 -316 175 -282
<< psubdiffcont >>
rect -79 282 79 316
rect -175 -220 -141 220
rect 141 -220 175 220
rect -79 -316 79 -282
<< poly >>
rect -33 214 33 230
rect -33 180 -17 214
rect 17 180 33 214
rect -33 164 33 180
rect -15 142 15 164
rect -15 -164 15 -142
rect -33 -180 33 -164
rect -33 -214 -17 -180
rect 17 -214 33 -180
rect -33 -230 33 -214
<< polycont >>
rect -17 180 17 214
rect -17 -214 17 -180
<< locali >>
rect -175 282 -79 316
rect 79 282 175 316
rect -175 220 -141 282
rect 141 220 175 282
rect -33 180 -17 214
rect 17 180 33 214
rect -61 130 -27 146
rect -61 -146 -27 -130
rect 27 130 61 146
rect 27 -146 61 -130
rect -33 -214 -17 -180
rect 17 -214 33 -180
rect -175 -282 -141 -220
rect 141 -282 175 -220
rect -175 -316 -79 -282
rect 79 -316 175 -282
<< viali >>
rect -17 180 17 214
rect -61 -130 -27 130
rect 27 -130 61 130
rect -17 -214 17 -180
<< metal1 >>
rect -29 214 29 220
rect -29 180 -17 214
rect 17 180 29 214
rect -29 174 29 180
rect -67 130 -21 142
rect -67 -130 -61 130
rect -27 -130 -21 130
rect -67 -142 -21 -130
rect 21 130 67 142
rect 21 -130 27 130
rect 61 -130 67 130
rect 21 -142 67 -130
rect -29 -180 29 -174
rect -29 -214 -17 -180
rect 17 -214 29 -180
rect -29 -220 29 -214
<< properties >>
string FIXED_BBOX -158 -299 158 299
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.42 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
