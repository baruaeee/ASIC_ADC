magic
tech sky130A
magscale 1 2
timestamp 1704404416
<< error_p >>
rect -29 114 29 120
rect -29 80 -17 114
rect -29 74 29 80
rect -29 -80 29 -74
rect -29 -114 -17 -80
rect -29 -120 29 -114
<< pwell >>
rect -215 -252 215 252
<< nmos >>
rect -19 -42 19 42
<< ndiff >>
rect -77 30 -19 42
rect -77 -30 -65 30
rect -31 -30 -19 30
rect -77 -42 -19 -30
rect 19 30 77 42
rect 19 -30 31 30
rect 65 -30 77 30
rect 19 -42 77 -30
<< ndiffc >>
rect -65 -30 -31 30
rect 31 -30 65 30
<< psubdiff >>
rect -179 182 -83 216
rect 83 182 179 216
rect -179 120 -145 182
rect 145 120 179 182
rect -179 -182 -145 -120
rect 145 -182 179 -120
rect -179 -216 -83 -182
rect 83 -216 179 -182
<< psubdiffcont >>
rect -83 182 83 216
rect -179 -120 -145 120
rect 145 -120 179 120
rect -83 -216 83 -182
<< poly >>
rect -33 114 33 130
rect -33 80 -17 114
rect 17 80 33 114
rect -33 64 33 80
rect -19 42 19 64
rect -19 -64 19 -42
rect -33 -80 33 -64
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -33 -130 33 -114
<< polycont >>
rect -17 80 17 114
rect -17 -114 17 -80
<< locali >>
rect -179 182 -83 216
rect 83 182 179 216
rect -179 120 -145 182
rect 145 120 179 182
rect -33 80 -17 114
rect 17 80 33 114
rect -65 30 -31 46
rect -65 -46 -31 -30
rect 31 30 65 46
rect 31 -46 65 -30
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -179 -182 -145 -120
rect 145 -182 179 -120
rect -179 -216 -83 -182
rect 83 -216 179 -182
<< viali >>
rect -17 80 17 114
rect -65 -30 -31 30
rect 31 -30 65 30
rect -17 -114 17 -80
<< metal1 >>
rect -29 114 29 120
rect -29 80 -17 114
rect 17 80 29 114
rect -29 74 29 80
rect -71 30 -25 42
rect -71 -30 -65 30
rect -31 -30 -25 30
rect -71 -42 -25 -30
rect 25 30 71 42
rect 25 -30 31 30
rect 65 -30 71 30
rect 25 -42 71 -30
rect -29 -80 29 -74
rect -29 -114 -17 -80
rect 17 -114 29 -80
rect -29 -120 29 -114
<< properties >>
string FIXED_BBOX -162 -199 162 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.193 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
