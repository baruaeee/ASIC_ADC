magic
tech sky130A
timestamp 1704418840
<< pwell >>
rect -173 -126 173 126
<< nmos >>
rect -75 -21 75 21
<< ndiff >>
rect -104 15 -75 21
rect -104 -15 -98 15
rect -81 -15 -75 15
rect -104 -21 -75 -15
rect 75 15 104 21
rect 75 -15 81 15
rect 98 -15 104 15
rect 75 -21 104 -15
<< ndiffc >>
rect -98 -15 -81 15
rect 81 -15 98 15
<< psubdiff >>
rect -155 91 -107 108
rect 107 91 155 108
rect -155 60 -138 91
rect 138 60 155 91
rect -155 -91 -138 -60
rect 138 -91 155 -60
rect -155 -108 -107 -91
rect 107 -108 155 -91
<< psubdiffcont >>
rect -107 91 107 108
rect -155 -60 -138 60
rect 138 -60 155 60
rect -107 -108 107 -91
<< poly >>
rect -75 57 75 65
rect -75 40 -67 57
rect 67 40 75 57
rect -75 21 75 40
rect -75 -40 75 -21
rect -75 -57 -67 -40
rect 67 -57 75 -40
rect -75 -65 75 -57
<< polycont >>
rect -67 40 67 57
rect -67 -57 67 -40
<< locali >>
rect -155 91 -107 108
rect 107 91 155 108
rect -155 60 -138 91
rect 138 60 155 91
rect -75 40 -67 57
rect 67 40 75 57
rect -98 15 -81 23
rect -98 -23 -81 -15
rect 81 15 98 23
rect 81 -23 98 -15
rect -75 -57 -67 -40
rect 67 -57 75 -40
rect -155 -91 -138 -60
rect 138 -91 155 -60
rect -155 -108 -107 -91
rect 107 -108 155 -91
<< viali >>
rect -67 40 67 57
rect -98 -15 -81 15
rect 81 -15 98 15
rect -67 -57 67 -40
<< metal1 >>
rect -73 57 73 60
rect -73 40 -67 57
rect 67 40 73 57
rect -73 37 73 40
rect -101 15 -78 21
rect -101 -15 -98 15
rect -81 -15 -78 15
rect -101 -21 -78 -15
rect 78 15 101 21
rect 78 -15 81 15
rect 98 -15 101 15
rect 78 -21 101 -15
rect -73 -40 73 -37
rect -73 -57 -67 -40
rect 67 -57 73 -40
rect -73 -60 73 -57
<< properties >>
string FIXED_BBOX -146 -99 146 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 1.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
