magic
tech sky130A
timestamp 1702941818
<< checkpaint >>
rect -649 1202 787 1226
rect -649 1178 944 1202
rect -649 1154 1147 1178
rect -649 1130 1396 1154
rect -649 1106 1553 1130
rect -649 1082 1802 1106
rect -649 1058 1959 1082
rect -649 1034 2116 1058
rect -649 1010 2273 1034
rect -649 986 2522 1010
rect -649 962 2771 986
rect -649 938 2928 962
rect -649 914 3131 938
rect -649 890 3288 914
rect -649 866 3491 890
rect -649 842 3786 866
rect -649 818 3943 842
rect -649 794 4192 818
rect -649 770 4441 794
rect -649 746 4690 770
rect -649 722 4939 746
rect -649 698 5280 722
rect -649 674 5483 698
rect -649 650 5732 674
rect -649 626 5935 650
rect -649 602 6276 626
rect -649 578 6571 602
rect -649 554 6866 578
rect -649 530 7207 554
rect -649 506 7548 530
rect -649 482 7843 506
rect -649 458 8000 482
rect -649 434 8203 458
rect -649 410 8360 434
rect -649 386 8609 410
rect -649 362 8812 386
rect -649 338 8969 362
rect -649 314 9172 338
rect -649 290 9467 314
rect -649 -354 9624 290
rect -630 -522 9624 -354
rect -630 -1830 730 -522
rect 837 -546 9624 -522
rect 994 -570 9624 -546
rect 1243 -594 9624 -570
rect 1492 -618 9624 -594
rect 1649 -642 9624 -618
rect 1852 -666 9624 -642
rect 2009 -690 9624 -666
rect 2212 -714 9624 -690
rect 2507 -738 9624 -714
rect 2664 -762 9624 -738
rect 2913 -786 9624 -762
rect 3162 -810 9624 -786
rect 3411 -834 9624 -810
rect 3660 -858 9624 -834
rect 4001 -882 9624 -858
rect 4204 -906 9624 -882
rect 4453 -930 9624 -906
rect 4656 -954 9624 -930
rect 4997 -978 9624 -954
rect 5292 -1002 9624 -978
rect 5587 -1026 9624 -1002
rect 5928 -1050 9624 -1026
rect 6269 -1074 9624 -1050
rect 6564 -1098 9624 -1074
rect 6721 -1122 9624 -1098
rect 6924 -1146 9624 -1122
rect 7081 -1170 9624 -1146
rect 7330 -1194 9624 -1170
rect 7533 -1218 9624 -1194
rect 7690 -1242 9624 -1218
rect 7893 -1266 9624 -1242
rect 8188 -1290 9624 -1266
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
use sky130_fd_sc_hd__clkinv_1  x0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 0 0 1 300
box -19 -24 157 296
use sky130_fd_sc_hd__nand2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 157 0 1 276
box -19 -24 157 296
use sky130_fd_sc_hd__nand3_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 314 0 1 252
box -19 -24 203 296
use sky130_fd_sc_hd__nand4_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 517 0 1 228
box -19 -24 249 296
use sky130_fd_sc_hd__nand2_1  x4
timestamp 1696625445
transform 1 0 766 0 1 204
box -19 -24 157 296
use sky130_fd_sc_hd__nand4_1  x5
timestamp 1696625445
transform 1 0 923 0 1 180
box -19 -24 249 296
use sky130_fd_sc_hd__nor2_1  x6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 1172 0 1 156
box -19 -24 157 296
use sky130_fd_sc_hd__nand2_1  x7
timestamp 1696625445
transform 1 0 1329 0 1 132
box -19 -24 157 296
use sky130_fd_sc_hd__nand2_1  x8
timestamp 1696625445
transform 1 0 1486 0 1 108
box -19 -24 157 296
use sky130_fd_sc_hd__nor4_1  x9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 1643 0 1 84
box -19 -24 249 296
use sky130_fd_sc_hd__and2_0  x10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 1892 0 1 60
box -19 -24 249 296
use sky130_fd_sc_hd__nand2_1  x11
timestamp 1696625445
transform 1 0 2141 0 1 36
box -19 -24 157 296
use sky130_fd_sc_hd__nand3_1  x12
timestamp 1696625445
transform 1 0 2298 0 1 12
box -19 -24 203 296
use sky130_fd_sc_hd__nor2_1  x13
timestamp 1696625445
transform 1 0 2501 0 1 -12
box -19 -24 157 296
use sky130_fd_sc_hd__nor3_1  x14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 2658 0 1 -36
box -19 -24 203 296
use sky130_fd_sc_hd__a22oi_1  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 2861 0 1 -60
box -19 -24 295 296
use sky130_fd_sc_hd__nor2_1  x16
timestamp 1696625445
transform 1 0 3156 0 1 -84
box -19 -24 157 296
use sky130_fd_sc_hd__or3_1  x17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3313 0 1 -108
box -19 -24 249 296
use sky130_fd_sc_hd__lpflow_inputiso1p_1  x18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 3562 0 1 -132
box -19 -24 249 296
use sky130_fd_sc_hd__nor4_1  x19
timestamp 1696625445
transform 1 0 3811 0 1 -156
box -19 -24 249 296
use sky130_fd_sc_hd__nand2b_1  x20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 4060 0 1 -180
box -19 -24 249 296
use sky130_fd_sc_hd__nor4b_1  x21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 4309 0 1 -204
box -19 -24 341 296
use sky130_fd_sc_hd__nor3_1  x22
timestamp 1696625445
transform 1 0 4650 0 1 -228
box -19 -24 203 296
use sky130_fd_sc_hd__nor4_1  x23
timestamp 1696625445
transform 1 0 4853 0 1 -252
box -19 -24 249 296
use sky130_fd_sc_hd__o21ai_0  x24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 5102 0 1 -276
box -19 -24 203 296
use sky130_fd_sc_hd__or3b_1  x25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 5305 0 1 -300
box -19 -24 341 296
use sky130_fd_sc_hd__or4_1  x26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 5646 0 1 -324
box -19 -24 295 296
use sky130_fd_sc_hd__a211oi_1  x27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 5941 0 1 -348
box -19 -24 295 296
use sky130_fd_sc_hd__a32oi_1  x28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 6236 0 1 -372
box -19 -24 341 296
use sky130_fd_sc_hd__o2111ai_1  x29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 6577 0 1 -396
box -19 -24 341 296
use sky130_fd_sc_hd__nand3b_1  x30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 6918 0 1 -420
box -19 -24 295 296
use sky130_fd_sc_hd__nand2_1  x31
timestamp 1696625445
transform 1 0 7213 0 1 -444
box -19 -24 157 296
use sky130_fd_sc_hd__nor3_1  x32
timestamp 1696625445
transform 1 0 7370 0 1 -468
box -19 -24 203 296
use sky130_fd_sc_hd__nand2_1  x33
timestamp 1696625445
transform 1 0 7573 0 1 -492
box -19 -24 157 296
use sky130_fd_sc_hd__nand4_1  x34
timestamp 1696625445
transform 1 0 7730 0 1 -516
box -19 -24 249 296
use sky130_fd_sc_hd__o21ai_0  x35
timestamp 1696625445
transform 1 0 7979 0 1 -540
box -19 -24 203 296
use sky130_fd_sc_hd__nor2_1  x36
timestamp 1696625445
transform 1 0 8182 0 1 -564
box -19 -24 157 296
use sky130_fd_sc_hd__o21ai_0  x37
timestamp 1696625445
transform 1 0 8339 0 1 -588
box -19 -24 203 296
use sky130_fd_sc_hd__o31ai_1  x38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1696625445
transform 1 0 8542 0 1 -612
box -19 -24 295 296
use sky130_fd_sc_hd__nand2_1  x39
timestamp 1696625445
transform 1 0 8837 0 1 -636
box -19 -24 157 296
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 Vp
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 Vin
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 b0
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 b1
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 b2
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 b3
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 128 0 0 0 Vn
port 6 nsew
<< end >>
