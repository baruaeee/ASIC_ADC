magic
tech sky130A
timestamp 1703732895
<< pwell >>
rect -1298 -126 1298 126
<< nmos >>
rect -1200 -21 1200 21
<< ndiff >>
rect -1229 15 -1200 21
rect -1229 -15 -1223 15
rect -1206 -15 -1200 15
rect -1229 -21 -1200 -15
rect 1200 15 1229 21
rect 1200 -15 1206 15
rect 1223 -15 1229 15
rect 1200 -21 1229 -15
<< ndiffc >>
rect -1223 -15 -1206 15
rect 1206 -15 1223 15
<< psubdiff >>
rect -1280 91 -1232 108
rect 1232 91 1280 108
rect -1280 60 -1263 91
rect 1263 60 1280 91
rect -1280 -91 -1263 -60
rect 1263 -91 1280 -60
rect -1280 -108 -1232 -91
rect 1232 -108 1280 -91
<< psubdiffcont >>
rect -1232 91 1232 108
rect -1280 -60 -1263 60
rect 1263 -60 1280 60
rect -1232 -108 1232 -91
<< poly >>
rect -1200 57 1200 65
rect -1200 40 -1192 57
rect 1192 40 1200 57
rect -1200 21 1200 40
rect -1200 -40 1200 -21
rect -1200 -57 -1192 -40
rect 1192 -57 1200 -40
rect -1200 -65 1200 -57
<< polycont >>
rect -1192 40 1192 57
rect -1192 -57 1192 -40
<< locali >>
rect -1280 91 -1232 108
rect 1232 91 1280 108
rect -1280 60 -1263 91
rect 1263 60 1280 91
rect -1200 40 -1192 57
rect 1192 40 1200 57
rect -1223 15 -1206 23
rect -1223 -23 -1206 -15
rect 1206 15 1223 23
rect 1206 -23 1223 -15
rect -1200 -57 -1192 -40
rect 1192 -57 1200 -40
rect -1280 -91 -1263 -60
rect 1263 -91 1280 -60
rect -1280 -108 -1232 -91
rect 1232 -108 1280 -91
<< viali >>
rect -1192 40 1192 57
rect -1223 -15 -1206 15
rect 1206 -15 1223 15
rect -1192 -57 1192 -40
<< metal1 >>
rect -1198 57 1198 60
rect -1198 40 -1192 57
rect 1192 40 1198 57
rect -1198 37 1198 40
rect -1226 15 -1203 21
rect -1226 -15 -1223 15
rect -1206 -15 -1203 15
rect -1226 -21 -1203 -15
rect 1203 15 1226 21
rect 1203 -15 1206 15
rect 1223 -15 1226 15
rect 1203 -21 1226 -15
rect -1198 -40 1198 -37
rect -1198 -57 -1192 -40
rect 1192 -57 1198 -40
rect -1198 -60 1198 -57
<< properties >>
string FIXED_BBOX -1271 -99 1271 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 24.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
