************************************************************************
* auCdl Netlist:
* 
* Library Name:  ADC
* Top Cell Name: inv03f
* View Name:     schematic
* Netlisted on:  Nov 18 14:04:15 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: ADC
* Cell Name:    inv03f
* View Name:    schematic
************************************************************************

.SUBCKT inv03f A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MNM1 Y A VSS VSS nfet_01v8 W=765n L=295n M=1
MPM1 Y A VDD VDD pfet_01v8 W=630n L=345n M=1
.ENDS

