magic
tech sky130A
magscale 1 2
timestamp 1703732895
<< error_p >>
rect -29 373 29 379
rect -29 339 -17 373
rect -29 333 29 339
rect -29 -339 29 -333
rect -29 -373 -17 -339
rect -29 -379 29 -373
<< nwell >>
rect -211 -511 211 511
<< pmos >>
rect -15 -292 15 292
<< pdiff >>
rect -73 280 -15 292
rect -73 -280 -61 280
rect -27 -280 -15 280
rect -73 -292 -15 -280
rect 15 280 73 292
rect 15 -280 27 280
rect 61 -280 73 280
rect 15 -292 73 -280
<< pdiffc >>
rect -61 -280 -27 280
rect 27 -280 61 280
<< nsubdiff >>
rect -175 441 -79 475
rect 79 441 175 475
rect -175 379 -141 441
rect 141 379 175 441
rect -175 -441 -141 -379
rect 141 -441 175 -379
rect -175 -475 -79 -441
rect 79 -475 175 -441
<< nsubdiffcont >>
rect -79 441 79 475
rect -175 -379 -141 379
rect 141 -379 175 379
rect -79 -475 79 -441
<< poly >>
rect -33 373 33 389
rect -33 339 -17 373
rect 17 339 33 373
rect -33 323 33 339
rect -15 292 15 323
rect -15 -323 15 -292
rect -33 -339 33 -323
rect -33 -373 -17 -339
rect 17 -373 33 -339
rect -33 -389 33 -373
<< polycont >>
rect -17 339 17 373
rect -17 -373 17 -339
<< locali >>
rect -175 441 -79 475
rect 79 441 175 475
rect -175 379 -141 441
rect 141 379 175 441
rect -33 339 -17 373
rect 17 339 33 373
rect -61 280 -27 296
rect -61 -296 -27 -280
rect 27 280 61 296
rect 27 -296 61 -280
rect -33 -373 -17 -339
rect 17 -373 33 -339
rect -175 -441 -141 -379
rect 141 -441 175 -379
rect -175 -475 -79 -441
rect 79 -475 175 -441
<< viali >>
rect -17 339 17 373
rect -61 -280 -27 280
rect 27 -280 61 280
rect -17 -373 17 -339
<< metal1 >>
rect -29 373 29 379
rect -29 339 -17 373
rect 17 339 29 373
rect -29 333 29 339
rect -67 280 -21 292
rect -67 -280 -61 280
rect -27 -280 -21 280
rect -67 -292 -21 -280
rect 21 280 67 292
rect 21 -280 27 280
rect 61 -280 67 280
rect 21 -292 67 -280
rect -29 -339 29 -333
rect -29 -373 -17 -339
rect 17 -373 29 -339
rect -29 -379 29 -373
<< properties >>
string FIXED_BBOX -158 -458 158 458
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.92 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
