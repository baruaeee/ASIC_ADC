magic
tech sky130A
magscale 1 2
timestamp 1706663412
<< pwell >>
rect 1376 -640 1410 -580
rect 1354 -756 1388 -696
<< psubdiff >>
rect 1119 -842 1221 -808
<< nsubdiff >>
rect 875 396 964 430
<< locali >>
rect 909 396 964 430
rect 1123 -842 1214 -808
rect 1332 -842 1408 -696
<< viali >>
rect 875 396 909 430
<< metal1 >>
rect 834 430 934 468
rect 834 429 875 430
rect 501 396 875 429
rect 909 396 934 430
rect 501 395 934 396
rect 501 229 535 395
rect 834 368 934 395
rect 644 290 708 344
rect 617 229 651 237
rect 501 195 651 229
rect 881 222 915 368
rect 1169 223 1203 233
rect 617 171 651 195
rect 705 187 815 221
rect 881 188 1046 222
rect 1169 189 1410 223
rect 471 87 703 121
rect 781 105 815 187
rect 1169 169 1203 189
rect 1072 105 1142 118
rect 471 -370 505 87
rect 781 71 1323 105
rect 604 -127 1167 -93
rect 604 -181 638 -127
rect 1131 -139 1167 -127
rect 1131 -173 1187 -139
rect 1133 -175 1187 -173
rect 714 -202 868 -184
rect 714 -214 730 -202
rect 724 -254 730 -214
rect 782 -214 868 -202
rect 782 -254 788 -214
rect 468 -470 568 -370
rect 471 -734 505 -470
rect 1059 -600 1065 -596
rect 577 -654 583 -602
rect 635 -654 650 -602
rect 1036 -648 1065 -600
rect 1117 -648 1123 -596
rect 1036 -658 1106 -648
rect 679 -734 879 -707
rect 471 -768 879 -734
rect 1153 -776 1187 -175
rect 1289 -401 1323 71
rect 1230 -435 1323 -401
rect 1376 -344 1410 189
rect 1230 -493 1264 -435
rect 1376 -444 1500 -344
rect 1216 -499 1268 -493
rect 1216 -557 1268 -551
rect 1230 -684 1264 -557
rect 1376 -605 1410 -444
rect 1331 -639 1410 -605
rect 1376 -640 1410 -639
rect 1331 -729 1409 -695
rect 1454 -698 1506 -634
rect 1153 -817 1254 -776
rect 1154 -839 1254 -817
rect 1354 -839 1389 -729
rect 1154 -873 1389 -839
rect 1154 -876 1254 -873
<< via1 >>
rect 730 -254 782 -202
rect 583 -654 635 -602
rect 1065 -648 1117 -596
rect 1216 -551 1268 -499
<< metal2 >>
rect 730 -202 782 -196
rect 724 -254 730 -248
rect 724 -260 782 -254
rect 724 -267 773 -260
rect 592 -301 773 -267
rect 592 -596 626 -301
rect 1210 -508 1216 -499
rect 1074 -542 1216 -508
rect 1074 -590 1108 -542
rect 1210 -551 1216 -542
rect 1268 -551 1274 -499
rect 1065 -596 1117 -590
rect 583 -602 635 -596
rect 1065 -654 1117 -648
rect 583 -660 635 -654
use sky130_fd_pr__pfet_01v8_XGAKDL  XM0
timestamp 1706241174
transform 0 -1 885 1 0 -155
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_4X3CDA  XM1
timestamp 1706241174
transform 1 0 844 0 1 -628
box -376 -252 376 252
use sky130_fd_pr__pfet_01v8_MWB9BZ  XM2
timestamp 1706241174
transform 1 0 677 0 1 206
box -211 -262 211 262
use sky130_fd_pr__pfet_01v8_JM8GTH  XM3
timestamp 1706231216
transform 1 0 1106 0 1 205
box -246 -261 246 261
use sky130_fd_pr__nfet_01v8_L9ESAD  XM4
timestamp 1706241174
transform 0 -1 1370 1 0 -667
box -211 -260 211 260
<< labels >>
flabel metal1 468 -470 568 -370 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 1154 -876 1254 -776 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 834 368 934 468 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 1400 -444 1500 -344 0 FreeSans 256 0 0 0 V11
port 1 nsew
<< end >>
