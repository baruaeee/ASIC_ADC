magic
tech sky130A
magscale 1 2
timestamp 1706473616
<< psubdiff >>
rect 1648 -517 1682 -459
<< viali >>
rect 949 658 983 692
rect 1023 92 1057 126
rect 1648 -493 1682 -459
<< metal1 >>
rect 526 727 626 728
rect 526 693 1092 727
rect 526 628 679 693
rect 937 692 995 693
rect 937 658 949 692
rect 983 658 995 692
rect 937 652 995 658
rect 617 601 679 628
rect 645 495 679 601
rect 645 423 707 495
rect 891 469 925 503
rect 891 435 999 469
rect 1058 436 1092 693
rect 1787 437 1859 497
rect 891 419 925 435
rect 965 373 999 435
rect 736 336 864 362
rect 736 328 776 336
rect 828 328 864 336
rect 965 339 1427 373
rect 776 278 828 284
rect 965 239 999 339
rect 965 205 1156 239
rect 1825 227 1859 437
rect 1825 216 1893 227
rect 1825 205 1974 216
rect 713 135 813 159
rect 1017 135 1059 139
rect 713 126 1063 135
rect 713 125 1023 126
rect 771 93 1023 125
rect 641 -11 707 63
rect 641 -285 675 -11
rect 771 -73 819 93
rect 1017 92 1023 93
rect 1057 92 1063 126
rect 1017 59 1063 92
rect 711 -107 819 -73
rect 1021 -49 1063 59
rect 1122 -2 1156 205
rect 1652 171 1974 205
rect 1652 77 1686 171
rect 1874 116 1974 171
rect 1241 43 1686 77
rect 1652 42 1686 43
rect 1770 36 1776 42
rect 1736 32 1776 36
rect 1734 -2 1776 32
rect 1736 -10 1776 -2
rect 1828 -10 1834 42
rect 1239 -49 1417 -13
rect 1021 -91 1417 -49
rect 881 -202 887 -150
rect 939 -164 945 -150
rect 939 -198 1416 -164
rect 939 -202 963 -198
rect 929 -212 963 -202
rect 1563 -250 1569 -248
rect 1132 -251 1166 -250
rect 1132 -276 1199 -251
rect 1132 -285 1166 -276
rect 641 -318 1179 -285
rect 1534 -300 1569 -250
rect 1621 -300 1627 -248
rect 1534 -310 1568 -300
rect 568 -394 668 -366
rect 730 -394 782 -390
rect 568 -396 784 -394
rect 568 -448 730 -396
rect 782 -448 784 -396
rect 1750 -446 1850 -428
rect 568 -450 784 -448
rect 568 -466 668 -450
rect 730 -454 782 -450
rect 1636 -459 1850 -446
rect 1636 -493 1648 -459
rect 1682 -493 1850 -459
rect 1636 -505 1850 -493
rect 1750 -528 1850 -505
<< via1 >>
rect 776 284 828 336
rect 1776 -10 1828 42
rect 887 -202 939 -150
rect 1569 -300 1621 -248
rect 730 -448 782 -396
<< metal2 >>
rect 770 284 776 336
rect 828 327 834 336
rect 828 293 930 327
rect 828 284 834 293
rect 896 -144 930 293
rect 1776 42 1828 48
rect 1776 -16 1828 -10
rect 1785 -115 1819 -16
rect 887 -150 939 -144
rect 887 -208 939 -202
rect 1578 -149 1819 -115
rect 724 -448 730 -396
rect 782 -405 788 -396
rect 896 -405 930 -208
rect 1578 -242 1612 -149
rect 1569 -248 1621 -242
rect 1569 -306 1621 -300
rect 782 -439 930 -405
rect 782 -448 788 -439
use sky130_fd_pr__pfet_01v8_HPNF99  XM0
timestamp 1706473616
transform 1 0 743 0 1 25
box -219 -269 219 269
use sky130_fd_pr__nfet_01v8_JZU22M  XM1
timestamp 1706400305
transform 1 0 1367 0 1 -280
box -351 -252 351 252
use sky130_fd_pr__pfet_01v8_TM5S5A  XM2
timestamp 1706457568
transform 1 0 800 0 1 459
box -276 -269 276 269
use sky130_fd_pr__pfet_01v8_AM8GZ5  XM3
timestamp 1706454272
transform 1 0 1446 0 1 467
box -526 -261 526 261
use sky130_fd_pr__nfet_01v8_H7HSAV  XM4
timestamp 1706454272
transform 0 1 1446 1 0 15
box -211 -460 157 460
<< labels >>
flabel metal1 1874 116 1974 216 0 FreeSans 256 0 0 0 V14
port 1 nsew
flabel metal1 526 628 626 728 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 1750 -528 1850 -428 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 568 -466 668 -366 0 FreeSans 256 0 0 0 Vin
port 2 nsew
<< end >>
