magic
tech sky130A
magscale 1 2
timestamp 1706231216
<< pwell >>
rect 436 -852 470 -792
<< psubdiff >>
rect 605 -940 703 -906
<< nsubdiff >>
rect 601 -68 704 -34
<< locali >>
rect 269 -67 631 -33
rect 665 -67 704 -34
rect 269 -251 304 -67
rect 611 -68 704 -67
rect 269 -285 383 -251
rect 422 -940 482 -792
rect 603 -940 699 -906
rect 798 -940 858 -792
<< viali >>
rect 631 -67 665 -33
<< metal1 >>
rect 608 -33 708 2
rect 608 -67 631 -33
rect 665 -67 708 -33
rect 608 -98 708 -67
rect 536 -229 570 -228
rect 505 -289 570 -229
rect 645 -242 679 -98
rect 645 -276 786 -242
rect 897 -273 1053 -239
rect 263 -387 479 -353
rect 263 -420 297 -387
rect 200 -463 300 -420
rect 200 -520 340 -463
rect 290 -548 340 -520
rect 306 -782 340 -548
rect 536 -521 570 -289
rect 690 -385 871 -351
rect 690 -521 724 -385
rect 1019 -420 1053 -273
rect 980 -513 1080 -420
rect 536 -555 724 -521
rect 809 -520 1080 -513
rect 809 -547 1053 -520
rect 536 -569 570 -555
rect 437 -603 570 -569
rect 437 -737 471 -603
rect 436 -941 470 -792
rect 524 -796 580 -734
rect 690 -749 724 -555
rect 810 -555 1053 -547
rect 810 -738 844 -555
rect 690 -783 745 -749
rect 588 -941 688 -874
rect 813 -941 847 -793
rect 904 -796 964 -736
rect 436 -975 847 -941
use sky130_fd_pr__nfet_01v8_DD6SHA  XM0
timestamp 1706229878
transform 0 -1 452 1 0 -765
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_7DPLFP  XM1
timestamp 1706229878
transform 1 0 445 0 1 -259
box -245 -261 245 261
use sky130_fd_pr__pfet_01v8_MDPZBH  XM2
timestamp 1706229878
transform 1 0 840 0 1 -259
box -240 -261 240 261
use sky130_fd_pr__nfet_01v8_MYA4RC  XM3
timestamp 1706229878
transform 0 -1 828 1 0 -765
box -211 -256 211 256
<< labels >>
flabel metal1 980 -520 1080 -420 0 FreeSans 256 0 0 0 V06
port 2 nsew
flabel metal1 608 -98 708 2 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 200 -520 300 -420 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 588 -974 688 -874 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
