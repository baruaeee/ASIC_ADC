magic
tech sky130A
magscale 1 2
timestamp 1704135479
<< error_p >>
rect 80662 7523 80720 7529
rect 80662 7489 80674 7523
rect 80662 7483 80720 7489
rect 108165 7311 108223 7317
rect 108165 7277 108177 7311
rect 108165 7271 108223 7277
rect 80832 6526 80866 6544
rect 80832 6490 80902 6526
rect 80849 6456 80920 6490
rect 1221 4705 1256 4722
rect 1222 4704 1256 4705
rect 1222 4668 1292 4704
rect 3978 4668 4031 4669
rect 1239 4634 1310 4668
rect 3960 4634 4031 4668
rect 1239 4289 1309 4634
rect 3961 4633 4031 4634
rect 3978 4599 4049 4633
rect 4329 4599 4364 4616
rect 1239 4253 1292 4289
rect 3978 4236 4048 4599
rect 4330 4598 4364 4599
rect 4330 4562 4400 4598
rect 5586 4562 5639 4563
rect 4160 4531 4218 4537
rect 4160 4497 4172 4531
rect 4347 4528 4418 4562
rect 5568 4528 5639 4562
rect 4160 4491 4218 4497
rect 4160 4319 4218 4325
rect 4160 4285 4172 4319
rect 4160 4279 4218 4285
rect 3978 4200 4031 4236
rect 4347 4183 4417 4528
rect 5569 4527 5639 4528
rect 5586 4493 5657 4527
rect 6907 4493 6942 4510
rect 4347 4147 4400 4183
rect 5586 4130 5656 4493
rect 6908 4492 6942 4493
rect 6908 4456 6978 4492
rect 7294 4456 7347 4457
rect 6925 4422 6996 4456
rect 7276 4422 7347 4456
rect 5586 4094 5639 4130
rect 6925 4077 6995 4422
rect 7277 4421 7347 4422
rect 7294 4387 7365 4421
rect 10015 4387 10050 4404
rect 7107 4354 7165 4360
rect 7107 4320 7119 4354
rect 7107 4314 7165 4320
rect 7107 4160 7165 4166
rect 7107 4126 7119 4160
rect 7107 4120 7165 4126
rect 6925 4041 6978 4077
rect 7294 4024 7364 4387
rect 10016 4386 10050 4387
rect 10016 4350 10086 4386
rect 10033 4316 10104 4350
rect 7294 3988 7347 4024
rect 10033 3971 10103 4316
rect 10033 3935 10086 3971
rect 14677 2780 14711 2834
rect 19789 2816 19823 2834
rect 14507 2519 14565 2525
rect 14507 2485 14519 2519
rect 14507 2479 14565 2485
rect 14696 2383 14711 2780
rect 14730 2746 14765 2780
rect 14730 2383 14764 2746
rect 14730 2349 14745 2383
rect 19753 2330 19823 2816
rect 20105 2656 20139 2710
rect 19935 2413 19993 2419
rect 19935 2379 19947 2413
rect 19935 2373 19993 2379
rect 19753 2294 19806 2330
rect 20124 2277 20139 2656
rect 20158 2622 20193 2656
rect 25153 2622 25188 2656
rect 20158 2277 20192 2622
rect 25154 2603 25188 2622
rect 20158 2243 20173 2277
rect 25173 2224 25188 2603
rect 25207 2569 25242 2603
rect 30292 2569 30327 2603
rect 25207 2224 25241 2569
rect 30293 2550 30327 2569
rect 25207 2190 25222 2224
rect 30312 2171 30327 2550
rect 30346 2516 30381 2550
rect 30346 2171 30380 2516
rect 75123 2799 75158 2833
rect 80516 2816 80550 2834
rect 75124 2780 75158 2799
rect 75143 2383 75158 2780
rect 75177 2746 75212 2780
rect 75177 2383 75211 2746
rect 75177 2349 75192 2383
rect 80480 2330 80550 2816
rect 80662 2413 80720 2419
rect 80662 2379 80674 2413
rect 80662 2373 80720 2379
rect 80480 2294 80533 2330
rect 80849 2277 80919 6456
rect 81031 6388 81089 6394
rect 81031 6354 81043 6388
rect 81031 6348 81089 6354
rect 91569 2728 91604 2762
rect 96962 2756 96997 2763
rect 96962 2745 96996 2756
rect 81201 2639 81235 2657
rect 81201 2603 81271 2639
rect 81218 2569 81289 2603
rect 81031 2360 81089 2366
rect 81031 2326 81043 2360
rect 81031 2320 81089 2326
rect 80849 2241 80902 2277
rect 81218 2224 81288 2569
rect 81218 2188 81271 2224
rect 91570 2709 91604 2728
rect 91589 2330 91604 2709
rect 91623 2675 91658 2709
rect 91623 2330 91657 2675
rect 91623 2296 91638 2330
rect 96926 2277 96996 2745
rect 97113 2688 97171 2694
rect 97113 2654 97125 2688
rect 97113 2648 97171 2654
rect 97288 2621 97322 2675
rect 97113 2360 97171 2366
rect 97113 2326 97125 2360
rect 97113 2320 97171 2326
rect 96926 2241 96979 2277
rect 97307 2224 97322 2621
rect 97341 2587 97376 2621
rect 102626 2587 102661 2621
rect 108019 2604 108053 2622
rect 97341 2224 97375 2587
rect 102627 2568 102661 2587
rect 97341 2190 97356 2224
rect 102646 2171 102661 2568
rect 102680 2534 102715 2568
rect 102680 2171 102714 2534
rect 30346 2137 30361 2171
rect 102680 2137 102695 2171
rect 107983 2118 108053 2604
rect 108165 2201 108223 2207
rect 108165 2167 108177 2201
rect 108165 2161 108223 2167
rect 107983 2082 108036 2118
<< error_s >>
rect 86061 7647 86119 7653
rect 86061 7613 86073 7647
rect 86061 7607 86119 7613
rect 67385 5283 67443 5289
rect 67385 5249 67397 5283
rect 67385 5243 67443 5249
rect 67555 3726 67589 3744
rect 67555 3690 67625 3726
rect 67572 3656 67643 3690
rect 38171 3470 38229 3476
rect 38171 3436 38183 3470
rect 38171 3430 38229 3436
rect 57258 3231 57316 3237
rect 57258 3197 57270 3231
rect 57258 3191 57316 3197
rect 35684 3107 35742 3113
rect 35684 3073 35696 3107
rect 35684 3067 35742 3073
rect 60765 2948 60823 2954
rect 50703 2939 50756 2942
rect 50685 2906 50756 2939
rect 60765 2914 60777 2948
rect 55662 2909 55715 2910
rect 40325 2869 40360 2878
rect 42587 2869 42622 2887
rect 40289 2844 40360 2869
rect 42551 2868 42622 2869
rect 43841 2870 43899 2876
rect 50703 2872 50774 2906
rect 55644 2875 55715 2909
rect 60765 2908 60823 2914
rect 55645 2874 55715 2875
rect 35854 2798 35888 2816
rect 35854 2762 35924 2798
rect 38025 2763 38059 2781
rect 36650 2762 36703 2763
rect 35871 2728 35942 2762
rect 36632 2728 36703 2762
rect 35684 2519 35742 2525
rect 35684 2485 35696 2519
rect 35684 2479 35742 2485
rect 35871 2383 35941 2728
rect 36633 2727 36703 2728
rect 36650 2693 36721 2727
rect 35871 2347 35924 2383
rect 36650 2330 36720 2693
rect 36650 2294 36703 2330
rect 37989 2277 38059 2763
rect 38341 2603 38375 2657
rect 38171 2360 38229 2366
rect 38171 2326 38183 2360
rect 38171 2320 38229 2326
rect 37989 2241 38042 2277
rect 38360 2224 38375 2603
rect 38394 2569 38429 2603
rect 38394 2224 38428 2569
rect 40289 2383 40359 2844
rect 40471 2776 40529 2782
rect 40471 2742 40483 2776
rect 40641 2763 40675 2781
rect 41233 2763 41268 2772
rect 40471 2736 40529 2742
rect 40641 2727 40711 2763
rect 41197 2738 41268 2763
rect 40658 2693 40729 2727
rect 40471 2466 40529 2472
rect 40471 2432 40483 2466
rect 40471 2426 40529 2432
rect 40289 2347 40342 2383
rect 40658 2330 40728 2693
rect 40658 2294 40711 2330
rect 41197 2277 41267 2738
rect 41379 2670 41437 2676
rect 41379 2636 41391 2670
rect 41379 2630 41437 2636
rect 41549 2611 41583 2665
rect 41379 2360 41437 2366
rect 41379 2326 41391 2360
rect 41379 2320 41437 2326
rect 41197 2241 41250 2277
rect 41568 2224 41583 2611
rect 41602 2577 41637 2611
rect 41602 2224 41636 2577
rect 41748 2509 41806 2515
rect 41748 2475 41760 2509
rect 41748 2469 41806 2475
rect 42551 2383 42621 2868
rect 43841 2836 43853 2870
rect 50516 2837 50574 2843
rect 43841 2830 43899 2836
rect 44490 2806 44525 2824
rect 46147 2806 46182 2824
rect 47742 2808 47777 2826
rect 42733 2800 42791 2806
rect 42733 2766 42745 2800
rect 44490 2799 44561 2806
rect 46147 2799 46218 2806
rect 47742 2799 47813 2808
rect 42733 2760 42791 2766
rect 42903 2763 42937 2781
rect 43695 2763 43729 2781
rect 44491 2770 44561 2799
rect 46148 2770 46218 2799
rect 47743 2772 47813 2799
rect 48129 2777 48182 2808
rect 49661 2799 49696 2833
rect 50370 2816 50404 2834
rect 49662 2780 49696 2799
rect 42903 2727 42973 2763
rect 42920 2693 42991 2727
rect 42733 2466 42791 2472
rect 42733 2432 42745 2466
rect 42733 2426 42791 2432
rect 42551 2347 42604 2383
rect 42920 2330 42990 2693
rect 41748 2307 41806 2313
rect 41748 2273 41760 2307
rect 42920 2294 42973 2330
rect 43659 2277 43729 2763
rect 44508 2736 44579 2770
rect 44859 2763 44894 2770
rect 44859 2736 44930 2763
rect 44508 2383 44578 2736
rect 44860 2727 44930 2736
rect 46165 2736 46236 2770
rect 46516 2763 46551 2770
rect 46516 2736 46587 2763
rect 44877 2693 44948 2727
rect 45292 2693 45327 2710
rect 44690 2668 44748 2674
rect 44690 2634 44702 2668
rect 44690 2628 44748 2634
rect 44690 2466 44748 2472
rect 44690 2432 44702 2466
rect 44690 2426 44748 2432
rect 43841 2360 43899 2366
rect 43841 2326 43853 2360
rect 44508 2347 44561 2383
rect 44877 2330 44947 2693
rect 45293 2692 45327 2693
rect 45293 2656 45363 2692
rect 45310 2622 45381 2656
rect 43841 2320 43899 2326
rect 44877 2294 44930 2330
rect 45310 2277 45380 2622
rect 45492 2554 45550 2560
rect 45492 2520 45504 2554
rect 45492 2514 45550 2520
rect 46165 2383 46235 2736
rect 46517 2727 46587 2736
rect 47760 2738 47831 2772
rect 48129 2743 48200 2777
rect 46534 2693 46605 2727
rect 46885 2693 46920 2710
rect 46347 2668 46405 2674
rect 46347 2634 46359 2668
rect 46347 2628 46405 2634
rect 46347 2466 46405 2472
rect 46347 2432 46359 2466
rect 46347 2426 46405 2432
rect 45492 2360 45550 2366
rect 45492 2326 45504 2360
rect 46165 2347 46218 2383
rect 46534 2330 46604 2693
rect 46886 2692 46920 2693
rect 46886 2656 46956 2692
rect 46716 2625 46774 2631
rect 46716 2591 46728 2625
rect 46903 2622 46974 2656
rect 46716 2585 46774 2591
rect 46716 2413 46774 2419
rect 46716 2379 46728 2413
rect 46716 2373 46774 2379
rect 45492 2320 45550 2326
rect 46534 2294 46587 2330
rect 46903 2277 46973 2622
rect 47086 2554 47144 2560
rect 47086 2520 47098 2554
rect 47086 2514 47144 2520
rect 47760 2383 47830 2738
rect 47942 2670 48000 2676
rect 47942 2636 47954 2670
rect 47942 2630 48000 2636
rect 47942 2466 48000 2472
rect 47942 2432 47954 2466
rect 47942 2426 48000 2432
rect 47086 2360 47144 2366
rect 47086 2326 47098 2360
rect 47760 2347 47813 2383
rect 48129 2330 48199 2743
rect 48481 2692 48515 2710
rect 48311 2675 48369 2681
rect 48311 2641 48323 2675
rect 48481 2656 48551 2692
rect 48311 2635 48369 2641
rect 48498 2622 48569 2656
rect 48311 2413 48369 2419
rect 48311 2379 48323 2413
rect 48311 2373 48369 2379
rect 47086 2320 47144 2326
rect 48129 2294 48182 2330
rect 48498 2277 48568 2622
rect 49681 2383 49696 2780
rect 49715 2746 49750 2780
rect 49715 2383 49749 2746
rect 49715 2349 49730 2383
rect 50334 2330 50404 2816
rect 50516 2803 50528 2837
rect 50516 2797 50574 2803
rect 50516 2413 50574 2419
rect 50516 2379 50528 2413
rect 50516 2373 50574 2379
rect 50334 2294 50387 2330
rect 50703 2277 50773 2872
rect 55662 2840 55733 2874
rect 50885 2804 50943 2810
rect 50885 2770 50897 2804
rect 52131 2799 52166 2816
rect 52132 2798 52166 2799
rect 52554 2809 52589 2816
rect 52554 2798 52588 2809
rect 54652 2799 54687 2833
rect 55329 2816 55363 2834
rect 50885 2764 50943 2770
rect 52132 2762 52202 2798
rect 51962 2731 52020 2737
rect 51962 2697 51974 2731
rect 52149 2728 52220 2762
rect 51962 2691 52020 2697
rect 51055 2639 51089 2657
rect 51055 2603 51125 2639
rect 51072 2569 51143 2603
rect 50885 2360 50943 2366
rect 50885 2326 50897 2360
rect 50885 2320 50943 2326
rect 41748 2267 41806 2273
rect 43659 2241 43712 2277
rect 45310 2241 45363 2277
rect 46903 2241 46956 2277
rect 48498 2241 48551 2277
rect 50703 2241 50756 2277
rect 51072 2224 51142 2569
rect 51962 2519 52020 2525
rect 51962 2485 51974 2519
rect 51962 2479 52020 2485
rect 52149 2383 52219 2728
rect 52331 2660 52389 2666
rect 52331 2626 52343 2660
rect 52331 2620 52389 2626
rect 52331 2466 52389 2472
rect 52331 2432 52343 2466
rect 52331 2426 52389 2432
rect 52149 2347 52202 2383
rect 52518 2330 52588 2798
rect 54653 2780 54687 2799
rect 52700 2741 52758 2747
rect 52700 2707 52712 2741
rect 52700 2701 52758 2707
rect 52870 2674 52904 2728
rect 52700 2413 52758 2419
rect 52700 2379 52712 2413
rect 52700 2373 52758 2379
rect 52518 2294 52571 2330
rect 52889 2277 52904 2674
rect 52923 2640 52958 2674
rect 53238 2640 53273 2674
rect 52923 2277 52957 2640
rect 53239 2621 53273 2640
rect 53069 2572 53127 2578
rect 53069 2538 53081 2572
rect 53069 2532 53127 2538
rect 53069 2360 53127 2366
rect 53069 2326 53081 2360
rect 53069 2320 53127 2326
rect 52923 2243 52938 2277
rect 53258 2224 53273 2621
rect 53292 2587 53327 2621
rect 53607 2587 53642 2604
rect 53292 2224 53326 2587
rect 53608 2586 53642 2587
rect 53608 2550 53678 2586
rect 53438 2519 53496 2525
rect 53438 2485 53450 2519
rect 53625 2516 53696 2550
rect 53438 2479 53496 2485
rect 53438 2307 53496 2313
rect 53438 2273 53450 2307
rect 53438 2267 53496 2273
rect 38394 2190 38409 2224
rect 41602 2190 41617 2224
rect 51072 2188 51125 2224
rect 53292 2190 53307 2224
rect 53625 2171 53695 2516
rect 53807 2448 53865 2454
rect 53807 2414 53819 2448
rect 53807 2408 53865 2414
rect 54672 2383 54687 2780
rect 54706 2746 54741 2780
rect 54706 2383 54740 2746
rect 54706 2349 54721 2383
rect 55293 2330 55363 2816
rect 55475 2807 55533 2813
rect 55475 2773 55487 2807
rect 55475 2767 55533 2773
rect 55475 2413 55533 2419
rect 55475 2379 55487 2413
rect 55475 2373 55533 2379
rect 55293 2294 55346 2330
rect 55662 2277 55732 2840
rect 57428 2798 57462 2816
rect 58404 2809 58439 2816
rect 58404 2798 58438 2809
rect 64086 2799 64121 2833
rect 67239 2816 67273 2834
rect 55844 2772 55902 2778
rect 55844 2738 55856 2772
rect 57428 2762 57498 2798
rect 55844 2732 55902 2738
rect 57445 2728 57516 2762
rect 56014 2639 56048 2657
rect 56690 2650 56725 2657
rect 56690 2639 56724 2650
rect 56014 2603 56084 2639
rect 56031 2569 56102 2603
rect 55844 2360 55902 2366
rect 55844 2326 55856 2360
rect 55844 2320 55902 2326
rect 53807 2254 53865 2260
rect 53807 2220 53819 2254
rect 55662 2241 55715 2277
rect 56031 2224 56101 2569
rect 53807 2214 53865 2220
rect 56031 2188 56084 2224
rect 56654 2171 56724 2639
rect 56836 2582 56894 2588
rect 56836 2548 56848 2582
rect 56836 2542 56894 2548
rect 57258 2519 57316 2525
rect 57258 2485 57270 2519
rect 57258 2479 57316 2485
rect 57445 2383 57515 2728
rect 57445 2347 57498 2383
rect 58368 2330 58438 2798
rect 64087 2780 64121 2799
rect 58550 2741 58608 2747
rect 58550 2707 58562 2741
rect 58550 2701 58608 2707
rect 58720 2674 58754 2728
rect 58550 2413 58608 2419
rect 58550 2379 58562 2413
rect 58550 2373 58608 2379
rect 58368 2294 58421 2330
rect 58739 2277 58754 2674
rect 58773 2640 58808 2674
rect 59642 2640 59677 2674
rect 60619 2657 60653 2675
rect 58773 2277 58807 2640
rect 59643 2621 59677 2640
rect 56836 2254 56894 2260
rect 56836 2220 56848 2254
rect 58773 2243 58788 2277
rect 59662 2224 59677 2621
rect 59696 2587 59731 2621
rect 59696 2224 59730 2587
rect 56836 2214 56894 2220
rect 59696 2190 59711 2224
rect 60583 2171 60653 2657
rect 64106 2383 64121 2780
rect 64140 2746 64175 2780
rect 64140 2383 64174 2746
rect 64140 2349 64155 2383
rect 67203 2330 67273 2816
rect 67385 2413 67443 2419
rect 67385 2379 67397 2413
rect 67385 2373 67443 2379
rect 67203 2294 67256 2330
rect 67572 2277 67642 3656
rect 67754 3588 67812 3594
rect 67754 3554 67766 3588
rect 67754 3548 67812 3554
rect 67924 2639 67958 2657
rect 69416 2650 69451 2657
rect 69416 2639 69450 2650
rect 67924 2603 67994 2639
rect 67941 2569 68012 2603
rect 67754 2360 67812 2366
rect 67754 2326 67766 2360
rect 67754 2320 67812 2326
rect 60765 2254 60823 2260
rect 60765 2220 60777 2254
rect 67572 2241 67625 2277
rect 67941 2224 68011 2569
rect 60765 2214 60823 2220
rect 67941 2188 67994 2224
rect 69380 2171 69450 2639
rect 69562 2582 69620 2588
rect 69562 2548 69574 2582
rect 69562 2542 69620 2548
rect 86231 2798 86265 2816
rect 86231 2762 86301 2798
rect 86248 2728 86319 2762
rect 85457 2622 85510 2639
rect 85457 2588 85528 2622
rect 69562 2254 69620 2260
rect 69562 2220 69574 2254
rect 69562 2214 69620 2220
rect 85457 2171 85527 2588
rect 85639 2520 85697 2526
rect 85639 2486 85651 2520
rect 86061 2519 86119 2525
rect 85639 2480 85697 2486
rect 86061 2485 86073 2519
rect 86061 2479 86119 2485
rect 86248 2383 86318 2728
rect 86248 2347 86301 2383
rect 85639 2254 85697 2260
rect 85639 2220 85651 2254
rect 85639 2214 85697 2220
rect 53625 2135 53678 2171
rect 56654 2135 56707 2171
rect 60583 2135 60636 2171
rect 69380 2135 69433 2171
rect 85457 2135 85510 2171
use th01  x1
timestamp 1704135479
transform 1 0 -1447 0 1 3706
box -53 -1200 14272 1069
use th02  x2
timestamp 1704135479
transform 1 0 14378 0 1 1800
box -53 -1200 21124 5785
use th03  x3
timestamp 1704135479
transform 1 0 35555 0 1 1800
box -53 -1200 4195 1808
use th04  x4
timestamp 1704135479
transform 1 0 39803 0 1 1800
box -53 -1200 2185 1114
use th05  x5
timestamp 1704135479
transform 1 0 42041 0 1 1800
box -53 -1200 2040 1208
use th06  x6
timestamp 1704135479
transform 1 0 44134 0 1 1800
box -53 -1200 1598 1069
use th07  x7
timestamp 1704135479
transform 1 0 45785 0 1 1800
box -53 -1200 1542 1069
use th08  x8
timestamp 1704135479
transform 1 0 47380 0 1 1800
box -53 -1200 1644 1069
use th09  x9
timestamp 1704135479
transform 1 0 49077 0 1 1800
box -53 -1200 2703 1175
use th10  x10
timestamp 1704135479
transform 1 0 51833 0 1 1800
box -53 -1200 2214 1079
use th11  x11
timestamp 1704135479
transform 1 0 54100 0 1 1800
box -53 -1200 2976 1145
use th12  x12
timestamp 1704135479
transform 1 0 57129 0 1 1800
box -53 -1200 3876 1569
use th13  x13
timestamp 1704135479
transform 1 0 61058 0 1 1800
box -53 -1200 8744 3621
use th14  x14
timestamp 1704135479
transform 1 0 69855 0 1 1800
box -53 -1200 16024 5861
use th15  x15
timestamp 1704135479
transform 1 0 85932 0 1 1800
box -53 -1200 22473 5985
<< end >>
