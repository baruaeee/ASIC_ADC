magic
tech sky130A
timestamp 1706204487
<< pwell >>
rect -175 -126 175 126
<< nmos >>
rect -77 -21 77 21
<< ndiff >>
rect -106 15 -77 21
rect -106 -15 -100 15
rect -83 -15 -77 15
rect -106 -21 -77 -15
rect 77 15 106 21
rect 77 -15 83 15
rect 100 -15 106 15
rect 77 -21 106 -15
<< ndiffc >>
rect -100 -15 -83 15
rect 83 -15 100 15
<< psubdiff >>
rect -157 60 -140 91
rect -157 -91 -140 -60
<< psubdiffcont >>
rect -157 -60 -140 60
<< poly >>
rect -77 57 77 65
rect -77 40 -69 57
rect 69 40 77 57
rect -77 21 77 40
rect -77 -40 77 -21
rect -77 -57 -69 -40
rect 69 -57 77 -40
rect -77 -65 77 -57
<< polycont >>
rect -69 40 69 57
rect -69 -57 69 -40
<< locali >>
rect -157 60 -140 91
rect -77 40 -69 57
rect 69 40 77 57
rect -100 15 -83 23
rect -100 -23 -83 -15
rect 83 15 100 23
rect 83 -23 100 -15
rect -77 -57 -69 -40
rect 69 -57 77 -40
rect -157 -91 -140 -60
<< viali >>
rect -69 40 69 57
rect -100 -15 -83 15
rect 83 -15 100 15
rect -69 -57 69 -40
<< metal1 >>
rect -75 57 75 60
rect -75 40 -69 57
rect 69 40 75 57
rect -75 37 75 40
rect -103 15 -80 21
rect -103 -15 -100 15
rect -83 -15 -80 15
rect -103 -21 -80 -15
rect 80 15 103 21
rect 80 -15 83 15
rect 100 -15 103 15
rect 80 -21 103 -15
rect -75 -40 75 -37
rect -75 -57 -69 -40
rect 69 -57 75 -40
rect -75 -60 75 -57
<< properties >>
string FIXED_BBOX -148 -99 148 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 1.54 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
