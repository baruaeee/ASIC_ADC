magic
tech sky130A
magscale 1 2
timestamp 1704674176
<< nwell >>
rect -828 -261 828 261
<< pmos >>
rect -632 -42 632 42
<< pdiff >>
rect -690 30 -632 42
rect -690 -30 -678 30
rect -644 -30 -632 30
rect -690 -42 -632 -30
rect 632 30 690 42
rect 632 -30 644 30
rect 678 -30 690 30
rect 632 -42 690 -30
<< pdiffc >>
rect -678 -30 -644 30
rect 644 -30 678 30
<< nsubdiff >>
rect -792 191 -696 225
rect 696 191 792 225
rect -792 129 -758 191
rect 758 129 792 191
rect -792 -191 -758 -129
rect 758 -191 792 -129
rect -792 -225 -696 -191
rect 696 -225 792 -191
<< nsubdiffcont >>
rect -696 191 696 225
rect -792 -129 -758 129
rect 758 -129 792 129
rect -696 -225 696 -191
<< poly >>
rect -632 123 632 139
rect -632 89 -616 123
rect 616 89 632 123
rect -632 42 632 89
rect -632 -89 632 -42
rect -632 -123 -616 -89
rect 616 -123 632 -89
rect -632 -139 632 -123
<< polycont >>
rect -616 89 616 123
rect -616 -123 616 -89
<< locali >>
rect -792 191 -696 225
rect 696 191 792 225
rect -792 129 -758 191
rect 758 129 792 191
rect -632 89 -616 123
rect 616 89 632 123
rect -678 30 -644 46
rect -678 -46 -644 -30
rect 644 30 678 46
rect 644 -46 678 -30
rect -632 -123 -616 -89
rect 616 -123 632 -89
rect -792 -191 -758 -129
rect 758 -191 792 -129
rect -792 -225 -696 -191
rect 696 -225 792 -191
<< viali >>
rect -616 89 616 123
rect -678 -30 -644 30
rect 644 -30 678 30
rect -616 -123 616 -89
<< metal1 >>
rect -628 123 628 129
rect -628 89 -616 123
rect 616 89 628 123
rect -628 83 628 89
rect -684 30 -638 42
rect -684 -30 -678 30
rect -644 -30 -638 30
rect -684 -42 -638 -30
rect 638 30 684 42
rect 638 -30 644 30
rect 678 -30 684 30
rect 638 -42 684 -30
rect -628 -89 628 -83
rect -628 -123 -616 -89
rect 616 -123 628 -89
rect -628 -129 628 -123
<< properties >>
string FIXED_BBOX -775 -208 775 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 6.323 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
