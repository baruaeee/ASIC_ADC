magic
tech sky130A
magscale 1 2
timestamp 1704302491
<< locali >>
rect 3416 1600 3580 1660
rect 3520 1568 3580 1600
rect 3520 1508 3988 1568
rect 3520 1486 3580 1508
rect 3390 1072 3482 1076
rect 3390 1016 3580 1072
rect 3520 268 3580 1016
rect 3928 774 3988 1508
rect 3372 208 3580 268
rect 1410 -328 3402 -268
rect 1410 -452 1470 -328
rect 3520 -352 3580 208
rect 3520 -412 4008 -352
rect 3520 -450 3580 -412
rect 1324 -512 1470 -452
rect 2060 -510 3580 -450
rect 3948 -422 4008 -412
rect 4246 -422 4306 -334
rect 3948 -482 4306 -422
rect 2060 -548 2120 -510
<< viali >>
rect 3520 1428 3580 1486
rect 3402 -328 3460 -268
rect 2060 -606 2120 -548
<< metal1 >>
rect 3149 1858 3659 1862
rect 3149 1804 3824 1858
rect 965 1619 1139 1677
rect 3149 1671 3207 1804
rect 965 562 1023 1619
rect 1249 1413 1307 1615
rect 3304 1612 3362 1670
rect 3624 1658 3824 1804
rect 3508 1486 3592 1492
rect 3508 1428 3520 1486
rect 3580 1483 3592 1486
rect 3624 1483 3682 1658
rect 3580 1455 3682 1483
rect 3580 1428 4105 1455
rect 3508 1425 4105 1428
rect 3508 1422 3592 1425
rect 1076 1355 3395 1413
rect 1076 902 1134 1355
rect 2543 1354 2601 1355
rect 3337 1331 3395 1355
rect 3624 1397 4105 1425
rect 3456 1331 3514 1336
rect 3337 1330 3514 1331
rect 3337 1273 3456 1330
rect 3456 1266 3514 1272
rect 1076 814 1152 902
rect 3265 845 3369 903
rect 3270 820 3369 845
rect 1088 812 1152 814
rect 960 490 1160 562
rect 1309 490 1367 781
rect 960 452 1368 490
rect 958 432 1368 452
rect 958 362 1160 432
rect 1309 430 1367 432
rect 3311 425 3369 820
rect 1475 367 3369 425
rect 958 -43 1016 362
rect 1475 285 1533 367
rect 1074 227 1533 285
rect 1074 6 1132 227
rect 3267 3 3357 91
rect 1172 -43 1280 -32
rect 958 -101 1283 -43
rect 3299 -185 3357 3
rect 3209 -243 3357 -185
rect 3209 -337 3267 -243
rect 915 -395 3267 -337
rect 3396 -268 3466 -256
rect 3396 -328 3402 -268
rect 3460 -270 3466 -268
rect 3624 -270 3682 1397
rect 6213 1379 6301 1469
rect 3753 1330 3811 1336
rect 3811 1311 3856 1324
rect 4189 1311 4234 1338
rect 3811 1272 4234 1311
rect 3753 1266 4234 1272
rect 3460 -328 3682 -270
rect 3811 563 3856 1266
rect 6243 1138 6301 1379
rect 4024 1080 6301 1138
rect 4024 701 4082 1080
rect 4024 607 4115 701
rect 4024 602 4082 607
rect 6229 603 6327 693
rect 3811 518 4188 563
rect 3811 -283 3856 518
rect 6269 280 6327 603
rect 5706 260 6327 280
rect 5706 222 6436 260
rect 5706 -281 5764 222
rect 6236 60 6436 222
rect 3811 -328 4113 -283
rect 3396 -340 3466 -328
rect 6178 -338 6238 -276
rect 915 -656 973 -395
rect 1148 -600 1216 -538
rect 1956 -548 2156 -540
rect 1956 -606 2060 -548
rect 2120 -606 2156 -548
rect 915 -714 1153 -656
rect 1209 -697 1339 -639
rect 1281 -783 1339 -697
rect 1956 -783 2156 -606
rect 1149 -841 2156 -783
rect 1956 -912 2156 -841
<< via1 >>
rect 3456 1272 3514 1330
rect 3753 1272 3811 1330
<< metal2 >>
rect 3450 1272 3456 1330
rect 3514 1272 3753 1330
rect 3811 1272 3817 1330
use sky130_fd_pr__pfet_01v8_MYW2PY  XM0
timestamp 1704301096
transform 1 0 1183 0 1 -683
box -211 -267 211 267
use sky130_fd_pr__nfet_01v8_JRGCPP  XM1
timestamp 1704301096
transform 1 0 2206 0 1 50
box -1246 -252 1246 252
use sky130_fd_pr__nfet_01v8_JRGCPP  XM2
timestamp 1704301096
transform 1 0 2210 0 1 860
box -1246 -252 1246 252
use sky130_fd_pr__pfet_01v8_XJ78MR  XM3
timestamp 1704301096
transform 0 -1 2217 1 0 1643
box -211 -1269 211 1269
use sky130_fd_pr__pfet_01v8_6M437L  XM4
timestamp 1704301096
transform 1 0 5162 0 1 1427
box -1246 -261 1246 261
use sky130_fd_pr__nfet_01v8_A5ES5P  XM5
timestamp 1704301096
transform 0 -1 5148 1 0 -307
box -211 -1210 211 1210
use sky130_fd_pr__pfet_01v8_6M437L  XM7
timestamp 1704301096
transform 1 0 5170 0 1 651
box -1246 -261 1246 261
<< labels >>
flabel metal1 1956 -912 2156 -712 0 FreeSans 256 0 0 0 Vn
port 3 nsew
flabel metal1 3624 1658 3824 1858 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 960 362 1160 562 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 6236 60 6436 260 0 FreeSans 256 0 0 0 Vout
port 1 nsew
<< end >>
