magic
tech sky130A
magscale 1 2
timestamp 1705440694
<< locali >>
rect 558 -344 680 -198
rect 794 -978 964 -852
rect 682 -1102 824 -1046
<< metal1 >>
rect 488 -148 688 52
rect 550 -180 626 -148
rect 550 -228 1090 -180
rect 420 -413 513 -337
rect 550 -346 626 -228
rect 1207 -249 1319 -167
rect 1123 -333 1185 -299
rect 420 -598 466 -413
rect 567 -435 682 -401
rect 730 -402 786 -342
rect 1129 -395 1163 -333
rect 336 -742 536 -598
rect 332 -798 536 -742
rect 648 -613 682 -435
rect 1081 -429 1163 -395
rect 1081 -613 1115 -429
rect 1273 -474 1319 -249
rect 648 -647 1135 -613
rect 332 -1182 380 -798
rect 648 -849 682 -647
rect 1081 -837 1135 -647
rect 1196 -674 1396 -474
rect 451 -883 682 -849
rect 451 -1035 485 -883
rect 936 -938 1080 -890
rect 451 -1105 521 -1035
rect 678 -1112 786 -1038
rect 538 -1182 652 -1146
rect 330 -1230 660 -1182
rect 738 -1268 786 -1112
rect 936 -1192 984 -938
rect 1032 -966 1080 -938
rect 1133 -933 1179 -881
rect 1273 -933 1319 -674
rect 1133 -970 1319 -933
rect 1074 -1058 1136 -1010
rect 900 -1268 1100 -1192
rect 738 -1316 1100 -1268
rect 900 -1392 1100 -1316
use sky130_fd_pr__nfet_01v8_LNCAWD  XM0
timestamp 1704374400
transform 1 0 601 0 1 -1068
box -263 -252 263 252
use sky130_fd_pr__pfet_01v8_M6KFPY  XM1
timestamp 1704374400
transform 0 -1 624 1 0 -371
box -211 -286 211 286
use sky130_fd_pr__pfet_01v8_NZD9V2  XM2
timestamp 1704374400
transform 1 0 1153 0 1 -207
box -243 -261 243 261
use sky130_fd_pr__nfet_01v8_NCP4B2  XM3
timestamp 1704374400
transform 1 0 1107 0 1 -923
box -211 -257 211 257
<< labels >>
flabel metal1 488 -148 688 52 0 FreeSans 256 0 0 0 Vp
port 0 nsew
flabel metal1 336 -798 536 -598 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 1196 -674 1396 -474 0 FreeSans 256 0 0 0 V08
port 1 nsew
flabel metal1 900 -1392 1100 -1192 0 FreeSans 256 0 0 0 Vn
port 3 nsew
<< end >>
