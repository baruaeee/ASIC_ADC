************************************************************************
* auCdl Netlist:
* 
* Library Name:  ADC
* Top Cell Name: inv10f
* View Name:     schematic
* Netlisted on:  Dec  1 05:22:32 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: ADC
* Cell Name:    inv10f
* View Name:    schematic
************************************************************************

.SUBCKT inv10f A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MNM1 Y A VSS VSS nfet_01v8 W=945n L=155n M=1
MPM1 Y A VDD VDD pfet_01v8 W=865n L=245n M=1
.ENDS

