* NGSPICE file created from therm.ext - technology: scmos

* Black-box entry subcircuit for sky130_fd_sc_hs__fill_1 abstract view
.subckt sky130_fd_sc_hs__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__o21ai_1 abstract view
.subckt sky130_fd_sc_hs__o21ai_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__fill_4 abstract view
.subckt sky130_fd_sc_hs__fill_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nand3b_1 abstract view
.subckt sky130_fd_sc_hs__nand3b_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nand3_1 abstract view
.subckt sky130_fd_sc_hs__nand3_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__and2b_1 abstract view
.subckt sky130_fd_sc_hs__and2b_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nor3b_1 abstract view
.subckt sky130_fd_sc_hs__nor3b_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__diode_2 abstract view
.subckt sky130_fd_sc_hs__diode_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nor3_1 abstract view
.subckt sky130_fd_sc_hs__nor3_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__and3_1 abstract view
.subckt sky130_fd_sc_hs__and3_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__o2111ai_1 abstract view
.subckt sky130_fd_sc_hs__o2111ai_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nand2_1 abstract view
.subckt sky130_fd_sc_hs__nand2_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__buf_1 abstract view
.subckt sky130_fd_sc_hs__buf_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkinv_1 abstract view
.subckt sky130_fd_sc_hs__clkinv_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nor2_1 abstract view
.subckt sky130_fd_sc_hs__nor2_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__or3_1 abstract view
.subckt sky130_fd_sc_hs__or3_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hs__o2bb2ai_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__o221ai_1 abstract view
.subckt sky130_fd_sc_hs__o221ai_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__and2_1 abstract view
.subckt sky130_fd_sc_hs__and2_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__or2b_1 abstract view
.subckt sky130_fd_sc_hs__or2b_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__a41oi_1 abstract view
.subckt sky130_fd_sc_hs__a41oi_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hs__a2bb2oi_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nor3_2 abstract view
.subckt sky130_fd_sc_hs__nor3_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfrtp_1 abstract view
.subckt sky130_fd_sc_hs__dfrtp_1 RESET_B VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nand4_1 abstract view
.subckt sky130_fd_sc_hs__nand4_1 VGND VNB VPB VPWR
.ends

.subckt therm VPWR VGND clk rst p[0] p[1] p[2] p[3] p[4] p[5] p[6] p[7] p[8] p[9]
+ p[10] p[11] p[12] p[13] p[14] b[0] b[1] b[2] b[3]
Xsky130_fd_sc_hs__fill_1_0_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__o21ai_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__fill_1_5_0_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__fill_4_6_1_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__o21ai_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__fill_1_5_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__nand3b_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__nand3b_1
Xsky130_fd_sc_hs__fill_1_3_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__fill_4_1_0_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__nand3_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__nand3_1
Xsky130_fd_sc_hs__and2b_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__and2b_1
Xsky130_fd_sc_hs__fill_1_3_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__nand3_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__nand3_1
Xsky130_fd_sc_hs__and2b_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__and2b_1
Xsky130_fd_sc_hs__fill_1_6_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__nand3_1_3 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__nand3_1
Xsky130_fd_sc_hs__nor3b_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__nor3b_1
Xsky130_fd_sc_hs__diode_2_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__and2b_1_3 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__and2b_1
Xsky130_fd_sc_hs__fill_4_4_0_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__nand3_1_4 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__nand3_1
Xsky130_fd_sc_hs__diode_2_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__nand3_1_5 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__nand3_1
Xsky130_fd_sc_hs__diode_2_3 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__nor3_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__fill_1_1_0_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__fill_4_2_1_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__nor3_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__nand3_1_6 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__nand3_1
Xsky130_fd_sc_hs__and3_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__and3_1
Xsky130_fd_sc_hs__diode_2_4 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__nand3_1_7 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__nand3_1
Xsky130_fd_sc_hs__nor3_1_3 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__diode_2_5 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__and3_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__and3_1
Xsky130_fd_sc_hs__diode_2_6 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__fill_1_4_0_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__fill_4_5_1_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__diode_2_7 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__diode_2_8 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__fill_1_2_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__o2111ai_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__o2111ai_1
Xsky130_fd_sc_hs__diode_2_9 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__fill_4_0_0_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__nand2_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__buf_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__buf_1
Xsky130_fd_sc_hs__nand2_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__buf_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__buf_1
Xsky130_fd_sc_hs__fill_1_5_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__nand2_1_3 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__fill_4_3_0_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__clkinv_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__clkinv_1
Xsky130_fd_sc_hs__buf_1_3 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__buf_1
Xsky130_fd_sc_hs__nand2_1_4 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__fill_1_6_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__clkinv_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__clkinv_1
Xsky130_fd_sc_hs__buf_1_4 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__buf_1
Xsky130_fd_sc_hs__nand2_1_5 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__fill_1_0_0_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__or3_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__or3_1
Xsky130_fd_sc_hs__o2bb2ai_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__o2bb2ai_1
Xsky130_fd_sc_hs__nand2_1_6 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__fill_4_1_1_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__nor2_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__fill_4_6_0_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__o221ai_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__o221ai_1
Xsky130_fd_sc_hs__and2_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__o2bb2ai_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__o2bb2ai_1
Xsky130_fd_sc_hs__nor2_1_3 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__and2_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__fill_1_4_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__nor2_1_4 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__or2b_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__or2b_1
Xsky130_fd_sc_hs__diode_2_10 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__fill_1_3_0_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__a41oi_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__a41oi_1
Xsky130_fd_sc_hs__and2_1_3 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__a2bb2oi_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__a2bb2oi_1
Xsky130_fd_sc_hs__fill_4_4_1_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__nor2_1_5 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__diode_2_11 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__and2_1_4 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__and2_1
Xsky130_fd_sc_hs__nor2_1_6 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__diode_2_12 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__nor3_2_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__nor3_2
Xsky130_fd_sc_hs__fill_1_1_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__fill_1_2_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__diode_2_13 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__fill_1_6_0_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__nor2_1_7 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__diode_2_14 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__nor2_1_8 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__diode_2_15 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__dfrtp_1_1 sky130_fd_sc_hs__dfrtp_1_4/RESET_B VGND sky130_fd_sc_hs__or3_1_1/VNB
+ sky130_fd_sc_hs__or3_1_1/VPB VPWR sky130_fd_sc_hs__dfrtp_1
Xsky130_fd_sc_hs__fill_1_4_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__diode_2_16 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__fill_4_2_0_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__dfrtp_1_2 sky130_fd_sc_hs__dfrtp_1_4/RESET_B VGND sky130_fd_sc_hs__or3_1_1/VNB
+ sky130_fd_sc_hs__nor3_2_1/VPB VPWR sky130_fd_sc_hs__dfrtp_1
Xsky130_fd_sc_hs__nand4_1_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__nand4_1
Xsky130_fd_sc_hs__diode_2_17 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__dfrtp_1_3 sky130_fd_sc_hs__dfrtp_1_4/RESET_B VGND sky130_fd_sc_hs__or3_1_1/VNB
+ sky130_fd_sc_hs__buf_1_4/VPB VPWR sky130_fd_sc_hs__dfrtp_1
Xsky130_fd_sc_hs__nand4_1_2 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__nand4_1
Xsky130_fd_sc_hs__dfrtp_1_4 sky130_fd_sc_hs__dfrtp_1_4/RESET_B VGND sky130_fd_sc_hs__or3_1_1/VNB
+ sky130_fd_sc_hs__buf_1_4/VPB VPWR sky130_fd_sc_hs__dfrtp_1
Xsky130_fd_sc_hs__fill_4_0_1_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_2/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__nand4_1_3 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__nand4_1
Xsky130_fd_sc_hs__fill_4_5_0_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__fill_1_2_0_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__or3_1_1/VPB
+ VPWR sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__fill_4_3_1_0 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__nor3_2_1/VPB
+ VPWR sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__fill_1_7_1 VGND sky130_fd_sc_hs__or3_1_1/VNB sky130_fd_sc_hs__buf_1_4/VPB
+ VPWR sky130_fd_sc_hs__fill_1
.ends

